module ibex_load_store_unit (addr_incr_req_o,
    busy_o,
    clk_i,
    data_err_i,
    data_gnt_i,
    data_pmp_err_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    load_err_o,
    lsu_rdata_valid_o,
    lsu_req_done_o,
    lsu_req_i,
    lsu_resp_valid_o,
    lsu_sign_ext_i,
    lsu_we_i,
    perf_load_o,
    perf_store_o,
    rst_ni,
    store_err_o,
    adder_result_ex_i,
    addr_last_o,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    lsu_rdata_o,
    lsu_type_i,
    lsu_wdata_i);
 output addr_incr_req_o;
 output busy_o;
 input clk_i;
 input data_err_i;
 input data_gnt_i;
 input data_pmp_err_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 output load_err_o;
 output lsu_rdata_valid_o;
 output lsu_req_done_o;
 input lsu_req_i;
 output lsu_resp_valid_o;
 input lsu_sign_ext_i;
 input lsu_we_i;
 output perf_load_o;
 output perf_store_o;
 input rst_ni;
 output store_err_o;
 input [31:0] adder_result_ex_i;
 output [31:0] addr_last_o;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 output [31:0] lsu_rdata_o;
 input [1:0] lsu_type_i;
 input [31:0] lsu_wdata_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire clknet_0_clk_i;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire data_sign_ext_q;
 wire \data_type_q[0] ;
 wire \data_type_q[1] ;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire data_we_q;
 wire handle_misaligned_q;
 wire net208;
 wire \ls_fsm_cs[0] ;
 wire \ls_fsm_cs[1] ;
 wire \ls_fsm_cs[2] ;
 wire \ls_fsm_ns[0] ;
 wire \ls_fsm_ns[1] ;
 wire \ls_fsm_ns[2] ;
 wire lsu_err_q;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire pmp_err_q;
 wire \rdata_offset_q[0] ;
 wire \rdata_offset_q[1] ;
 wire \rdata_q[10] ;
 wire \rdata_q[11] ;
 wire \rdata_q[12] ;
 wire \rdata_q[13] ;
 wire \rdata_q[14] ;
 wire \rdata_q[15] ;
 wire \rdata_q[16] ;
 wire \rdata_q[17] ;
 wire \rdata_q[18] ;
 wire \rdata_q[19] ;
 wire \rdata_q[20] ;
 wire \rdata_q[21] ;
 wire \rdata_q[22] ;
 wire \rdata_q[23] ;
 wire \rdata_q[24] ;
 wire \rdata_q[25] ;
 wire \rdata_q[26] ;
 wire \rdata_q[27] ;
 wire \rdata_q[28] ;
 wire \rdata_q[29] ;
 wire \rdata_q[30] ;
 wire \rdata_q[31] ;
 wire \rdata_q[8] ;
 wire \rdata_q[9] ;
 wire net246;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net247;
 wire net248;
 wire clknet_3_0__leaf_clk_i;
 wire clknet_3_1__leaf_clk_i;
 wire clknet_3_2__leaf_clk_i;
 wire clknet_3_3__leaf_clk_i;
 wire clknet_3_4__leaf_clk_i;
 wire clknet_3_5__leaf_clk_i;
 wire clknet_3_6__leaf_clk_i;
 wire clknet_3_7__leaf_clk_i;

 sky130_fd_sc_hd__clkbuf_4 _0449_ (.A(\ls_fsm_cs[2] ),
    .X(_0065_));
 sky130_fd_sc_hd__buf_6 _0450_ (.A(\ls_fsm_cs[1] ),
    .X(_0066_));
 sky130_fd_sc_hd__or3_1 _0451_ (.A(_0065_),
    .B(_0066_),
    .C(\ls_fsm_cs[0] ),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_2 _0452_ (.A(_0067_),
    .X(net139));
 sky130_fd_sc_hd__clkinvlp_4 _0453_ (.A(handle_misaligned_q),
    .Y(_0432_));
 sky130_fd_sc_hd__buf_2 _0454_ (.A(_0066_),
    .X(_0068_));
 sky130_fd_sc_hd__buf_2 _0455_ (.A(pmp_err_q),
    .X(_0069_));
 sky130_fd_sc_hd__o21ai_1 _0456_ (.A1(_0069_),
    .A2(net34),
    .B1(\ls_fsm_cs[0] ),
    .Y(_0070_));
 sky130_fd_sc_hd__buf_4 _0457_ (.A(\ls_fsm_cs[0] ),
    .X(_0071_));
 sky130_fd_sc_hd__nand2_1 _0458_ (.A(_0071_),
    .B(_0069_),
    .Y(_0072_));
 sky130_fd_sc_hd__nor2b_1 _0459_ (.A(net34),
    .B_N(_0068_),
    .Y(_0073_));
 sky130_fd_sc_hd__a2bb2oi_1 _0460_ (.A1_N(_0068_),
    .A2_N(_0070_),
    .B1(_0072_),
    .B2(_0073_),
    .Y(_0074_));
 sky130_fd_sc_hd__buf_2 _0461_ (.A(_0444_),
    .X(_0075_));
 sky130_fd_sc_hd__buf_2 _0462_ (.A(lsu_type_i[0]),
    .X(_0076_));
 sky130_fd_sc_hd__nor2b_1 _0463_ (.A(_0075_),
    .B_N(_0076_),
    .Y(_0077_));
 sky130_fd_sc_hd__nor2b_1 _0464_ (.A(_0076_),
    .B_N(_0438_),
    .Y(_0078_));
 sky130_fd_sc_hd__nor4b_2 _0465_ (.A(\ls_fsm_cs[2] ),
    .B(_0066_),
    .C(\ls_fsm_cs[0] ),
    .D_N(net69),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_1 _0466_ (.A(net34),
    .Y(_0080_));
 sky130_fd_sc_hd__o311ai_1 _0467_ (.A1(net71),
    .A2(_0077_),
    .A3(_0078_),
    .B1(_0079_),
    .C1(_0080_),
    .Y(_0081_));
 sky130_fd_sc_hd__and2_0 _0468_ (.A(_0076_),
    .B(_0075_),
    .X(_0082_));
 sky130_fd_sc_hd__nor2_1 _0469_ (.A(_0076_),
    .B(_0438_),
    .Y(_0083_));
 sky130_fd_sc_hd__clkbuf_4 _0470_ (.A(net71),
    .X(_0084_));
 sky130_fd_sc_hd__inv_1 _0471_ (.A(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__o2111ai_1 _0472_ (.A1(_0082_),
    .A2(_0083_),
    .B1(net34),
    .C1(_0085_),
    .D1(_0079_),
    .Y(_0086_));
 sky130_fd_sc_hd__o211ai_1 _0473_ (.A1(_0065_),
    .A2(_0074_),
    .B1(_0081_),
    .C1(_0086_),
    .Y(\ls_fsm_ns[1] ));
 sky130_fd_sc_hd__nor2b_1 _0474_ (.A(_0069_),
    .B_N(_0071_),
    .Y(_0087_));
 sky130_fd_sc_hd__nor3b_1 _0475_ (.A(_0068_),
    .B(_0071_),
    .C_N(net69),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_1 _0476_ (.A(_0065_),
    .Y(_0089_));
 sky130_fd_sc_hd__o211ai_2 _0477_ (.A1(_0087_),
    .A2(_0088_),
    .B1(_0089_),
    .C1(_0080_),
    .Y(_0090_));
 sky130_fd_sc_hd__nor4b_1 _0478_ (.A(_0065_),
    .B(_0071_),
    .C(net34),
    .D_N(_0068_),
    .Y(_0091_));
 sky130_fd_sc_hd__o21ai_0 _0479_ (.A1(_0069_),
    .A2(net68),
    .B1(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _0480_ (.A(_0090_),
    .B(_0092_),
    .Y(\ls_fsm_ns[0] ));
 sky130_fd_sc_hd__inv_1 _0481_ (.A(_0069_),
    .Y(_0093_));
 sky130_fd_sc_hd__and2b_1 _0482_ (.A_N(\ls_fsm_cs[2] ),
    .B(_0066_),
    .X(_0094_));
 sky130_fd_sc_hd__and2b_1 _0483_ (.A_N(_0066_),
    .B(\ls_fsm_cs[2] ),
    .X(_0095_));
 sky130_fd_sc_hd__a31oi_2 _0484_ (.A1(_0093_),
    .A2(net34),
    .A3(_0094_),
    .B1(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__nor3_1 _0485_ (.A(_0071_),
    .B(net68),
    .C(_0096_),
    .Y(\ls_fsm_ns[2] ));
 sky130_fd_sc_hd__inv_1 _0486_ (.A(net1),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_1 _0487_ (.A(_0438_),
    .Y(_0097_));
 sky130_fd_sc_hd__buf_2 _0488_ (.A(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_4 _0489_ (.A(_0098_),
    .X(_0433_));
 sky130_fd_sc_hd__inv_1 _0490_ (.A(net12),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2b_1 _0491_ (.A_N(net33),
    .B(net68),
    .Y(_0099_));
 sky130_fd_sc_hd__a211o_1 _0492_ (.A1(_0066_),
    .A2(lsu_err_q),
    .B1(_0070_),
    .C1(\ls_fsm_cs[2] ),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _0493_ (.A(net34),
    .B(_0079_),
    .Y(_0101_));
 sky130_fd_sc_hd__o311ai_4 _0494_ (.A1(\ls_fsm_cs[0] ),
    .A2(_0096_),
    .A3(_0099_),
    .B1(_0100_),
    .C1(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__buf_6 _0495_ (.A(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0496_ (.A0(net107),
    .A1(net1),
    .S(_0103_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _0497_ (.A0(net108),
    .A1(net2),
    .S(_0103_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0498_ (.A0(net109),
    .A1(net3),
    .S(_0103_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0499_ (.A0(net110),
    .A1(net4),
    .S(_0103_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0500_ (.A0(net111),
    .A1(net5),
    .S(_0103_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0501_ (.A0(net112),
    .A1(net6),
    .S(_0103_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _0502_ (.A0(net113),
    .A1(net7),
    .S(_0103_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0503_ (.A0(net114),
    .A1(net8),
    .S(_0103_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0504_ (.A0(net115),
    .A1(net9),
    .S(_0103_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0505_ (.A0(net116),
    .A1(net10),
    .S(_0103_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_6 _0506_ (.A(_0102_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0507_ (.A0(net117),
    .A1(net11),
    .S(_0104_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0508_ (.A0(net118),
    .A1(net12),
    .S(_0104_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0509_ (.A0(net119),
    .A1(net13),
    .S(_0104_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0510_ (.A0(net120),
    .A1(net14),
    .S(_0104_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0511_ (.A0(net121),
    .A1(net15),
    .S(_0104_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0512_ (.A0(net122),
    .A1(net16),
    .S(_0104_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0513_ (.A0(net123),
    .A1(net17),
    .S(_0104_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0514_ (.A0(net124),
    .A1(net18),
    .S(_0104_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0515_ (.A0(net125),
    .A1(net19),
    .S(_0104_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0516_ (.A0(net126),
    .A1(net20),
    .S(_0104_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_6 _0517_ (.A(_0102_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0518_ (.A0(net127),
    .A1(net21),
    .S(_0105_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0519_ (.A0(net128),
    .A1(net22),
    .S(_0105_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0520_ (.A0(net129),
    .A1(net23),
    .S(_0105_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0521_ (.A0(net130),
    .A1(net24),
    .S(_0105_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0522_ (.A0(net131),
    .A1(net25),
    .S(_0105_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0523_ (.A0(net132),
    .A1(net26),
    .S(_0105_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0524_ (.A0(net133),
    .A1(net27),
    .S(_0105_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0525_ (.A0(net134),
    .A1(net28),
    .S(_0105_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0526_ (.A0(net135),
    .A1(net29),
    .S(_0105_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0527_ (.A0(net136),
    .A1(net30),
    .S(_0105_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0528_ (.A0(net137),
    .A1(net31),
    .S(_0102_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0529_ (.A0(net138),
    .A1(net32),
    .S(_0102_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2b_1 _0530_ (.A(_0066_),
    .B_N(net69),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ai_1 _0531_ (.A1(\ls_fsm_cs[0] ),
    .A2(_0106_),
    .B1(net34),
    .Y(_0107_));
 sky130_fd_sc_hd__a21oi_4 _0532_ (.A1(_0072_),
    .A2(_0107_),
    .B1(_0065_),
    .Y(_0108_));
 sky130_fd_sc_hd__mux2_1 _0533_ (.A0(data_sign_ext_q),
    .A1(net70),
    .S(_0108_),
    .X(_0032_));
 sky130_fd_sc_hd__buf_4 _0534_ (.A(\data_type_q[0] ),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0535_ (.A0(_0109_),
    .A1(_0076_),
    .S(_0108_),
    .X(_0033_));
 sky130_fd_sc_hd__buf_8 _0536_ (.A(\data_type_q[1] ),
    .X(_0110_));
 sky130_fd_sc_hd__buf_4 _0537_ (.A(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0538_ (.A0(_0111_),
    .A1(_0084_),
    .S(_0108_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0539_ (.A0(data_we_q),
    .A1(net104),
    .S(_0108_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_1 _0540_ (.A(_0069_),
    .B(net68),
    .Y(_0112_));
 sky130_fd_sc_hd__nor3_1 _0541_ (.A(_0068_),
    .B(_0071_),
    .C(net69),
    .Y(_0113_));
 sky130_fd_sc_hd__a211oi_1 _0542_ (.A1(_0112_),
    .A2(_0091_),
    .B1(_0113_),
    .C1(_0065_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_1 _0543_ (.A(_0071_),
    .Y(_0115_));
 sky130_fd_sc_hd__o31a_1 _0544_ (.A1(_0065_),
    .A2(_0068_),
    .A3(_0115_),
    .B1(_0092_),
    .X(_0116_));
 sky130_fd_sc_hd__or2b_1 _0545_ (.A(\ls_fsm_cs[2] ),
    .B_N(_0066_),
    .X(_0117_));
 sky130_fd_sc_hd__o211ai_1 _0546_ (.A1(_0082_),
    .A2(_0083_),
    .B1(_0117_),
    .C1(_0085_),
    .Y(_0118_));
 sky130_fd_sc_hd__a21oi_1 _0547_ (.A1(_0090_),
    .A2(_0114_),
    .B1(handle_misaligned_q),
    .Y(_0119_));
 sky130_fd_sc_hd__a41oi_1 _0548_ (.A1(_0090_),
    .A2(_0114_),
    .A3(_0116_),
    .A4(_0118_),
    .B1(_0119_),
    .Y(_0036_));
 sky130_fd_sc_hd__o21ai_0 _0549_ (.A1(_0069_),
    .A2(net33),
    .B1(_0094_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand2_1 _0550_ (.A(net33),
    .B(_0095_),
    .Y(_0121_));
 sky130_fd_sc_hd__a21oi_1 _0551_ (.A1(_0120_),
    .A2(_0121_),
    .B1(_0071_),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2b_1 _0552_ (.A_N(_0066_),
    .B(net68),
    .Y(_0123_));
 sky130_fd_sc_hd__a21oi_1 _0553_ (.A1(_0065_),
    .A2(_0123_),
    .B1(_0071_),
    .Y(_0124_));
 sky130_fd_sc_hd__nand2_1 _0554_ (.A(_0068_),
    .B(_0112_),
    .Y(_0125_));
 sky130_fd_sc_hd__o311ai_1 _0555_ (.A1(_0065_),
    .A2(_0068_),
    .A3(net69),
    .B1(_0124_),
    .C1(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__mux2_1 _0556_ (.A0(_0122_),
    .A1(lsu_err_q),
    .S(_0126_),
    .X(_0037_));
 sky130_fd_sc_hd__o21ai_0 _0557_ (.A1(_0068_),
    .A2(net69),
    .B1(net35),
    .Y(_0127_));
 sky130_fd_sc_hd__nand2_1 _0558_ (.A(_0089_),
    .B(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__o21ai_0 _0559_ (.A1(net35),
    .A2(_0123_),
    .B1(_0128_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2b_1 _0560_ (.A_N(net68),
    .B(_0068_),
    .Y(_0130_));
 sky130_fd_sc_hd__a21oi_1 _0561_ (.A1(_0124_),
    .A2(_0130_),
    .B1(_0069_),
    .Y(_0131_));
 sky130_fd_sc_hd__a21oi_1 _0562_ (.A1(_0115_),
    .A2(_0129_),
    .B1(_0131_),
    .Y(_0038_));
 sky130_fd_sc_hd__buf_2 _0563_ (.A(\rdata_offset_q[0] ),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_4 _0564_ (.A(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_4 _0565_ (.A(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_8 _0566_ (.A(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0567_ (.A0(_0135_),
    .A1(net1),
    .S(_0108_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_2 _0568_ (.A(\rdata_offset_q[1] ),
    .X(_0136_));
 sky130_fd_sc_hd__buf_4 _0569_ (.A(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__buf_4 _0570_ (.A(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__buf_8 _0571_ (.A(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0572_ (.A0(_0139_),
    .A1(net12),
    .S(_0108_),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_1 _0573_ (.A(_0089_),
    .B(_0123_),
    .Y(_0140_));
 sky130_fd_sc_hd__nor2_1 _0574_ (.A(_0112_),
    .B(_0117_),
    .Y(_0141_));
 sky130_fd_sc_hd__nor2_1 _0575_ (.A(\ls_fsm_cs[0] ),
    .B(data_we_q),
    .Y(_0142_));
 sky130_fd_sc_hd__o21ai_4 _0576_ (.A1(_0140_),
    .A2(_0141_),
    .B1(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__buf_6 _0577_ (.A(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0578_ (.A0(net66),
    .A1(\rdata_q[8] ),
    .S(_0144_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0579_ (.A0(net45),
    .A1(\rdata_q[18] ),
    .S(_0144_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0580_ (.A0(net46),
    .A1(\rdata_q[19] ),
    .S(_0144_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0581_ (.A0(net48),
    .A1(\rdata_q[20] ),
    .S(_0144_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0582_ (.A0(net49),
    .A1(\rdata_q[21] ),
    .S(_0144_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0583_ (.A0(net50),
    .A1(\rdata_q[22] ),
    .S(_0144_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(net51),
    .A1(\rdata_q[23] ),
    .S(_0144_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(net52),
    .A1(\rdata_q[24] ),
    .S(_0144_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0586_ (.A0(net53),
    .A1(\rdata_q[25] ),
    .S(_0144_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0587_ (.A0(net54),
    .A1(\rdata_q[26] ),
    .S(_0144_),
    .X(_0050_));
 sky130_fd_sc_hd__buf_6 _0588_ (.A(_0143_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(net55),
    .A1(\rdata_q[27] ),
    .S(_0145_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0590_ (.A0(net67),
    .A1(\rdata_q[9] ),
    .S(_0145_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(net56),
    .A1(\rdata_q[28] ),
    .S(_0145_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0592_ (.A0(net57),
    .A1(\rdata_q[29] ),
    .S(_0145_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0593_ (.A0(net59),
    .A1(\rdata_q[30] ),
    .S(_0145_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(net60),
    .A1(\rdata_q[31] ),
    .S(_0145_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0595_ (.A0(net37),
    .A1(\rdata_q[10] ),
    .S(_0145_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(net38),
    .A1(\rdata_q[11] ),
    .S(_0145_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0597_ (.A0(net39),
    .A1(\rdata_q[12] ),
    .S(_0145_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(net40),
    .A1(\rdata_q[13] ),
    .S(_0145_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0599_ (.A0(net41),
    .A1(\rdata_q[14] ),
    .S(_0143_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0600_ (.A0(net42),
    .A1(\rdata_q[15] ),
    .S(_0143_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0601_ (.A0(net43),
    .A1(\rdata_q[16] ),
    .S(_0143_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(net44),
    .A1(\rdata_q[17] ),
    .S(_0143_),
    .X(_0064_));
 sky130_fd_sc_hd__a21oi_1 _0603_ (.A1(_0071_),
    .A2(_0432_),
    .B1(_0117_),
    .Y(_0146_));
 sky130_fd_sc_hd__a21o_1 _0604_ (.A1(_0115_),
    .A2(_0095_),
    .B1(_0146_),
    .X(net106));
 sky130_fd_sc_hd__inv_1 _0605_ (.A(_0434_),
    .Y(_0147_));
 sky130_fd_sc_hd__mux2i_1 _0606_ (.A0(_0435_),
    .A1(_0147_),
    .S(_0076_),
    .Y(_0148_));
 sky130_fd_sc_hd__nand2_1 _0607_ (.A(_0084_),
    .B(_0438_),
    .Y(_0149_));
 sky130_fd_sc_hd__o21ai_1 _0608_ (.A1(_0084_),
    .A2(_0148_),
    .B1(_0149_),
    .Y(net170));
 sky130_fd_sc_hd__clkbuf_2 _0609_ (.A(_0440_),
    .X(_0150_));
 sky130_fd_sc_hd__nor2_1 _0610_ (.A(_0150_),
    .B(_0075_),
    .Y(_0151_));
 sky130_fd_sc_hd__nor2_1 _0611_ (.A(_0076_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__a21oi_1 _0612_ (.A1(_0098_),
    .A2(_0432_),
    .B1(_0084_),
    .Y(_0153_));
 sky130_fd_sc_hd__clkbuf_2 _0613_ (.A(_0442_),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_4 _0614_ (.A(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__o32a_1 _0615_ (.A1(_0084_),
    .A2(_0432_),
    .A3(_0152_),
    .B1(_0153_),
    .B2(_0155_),
    .X(net171));
 sky130_fd_sc_hd__nor2b_1 _0616_ (.A(_0446_),
    .B_N(handle_misaligned_q),
    .Y(_0156_));
 sky130_fd_sc_hd__a211oi_1 _0617_ (.A1(_0432_),
    .A2(_0075_),
    .B1(_0156_),
    .C1(_0076_),
    .Y(_0157_));
 sky130_fd_sc_hd__a31oi_2 _0618_ (.A1(_0076_),
    .A2(_0432_),
    .A3(_0439_),
    .B1(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__clkbuf_4 _0619_ (.A(_0150_),
    .X(_0159_));
 sky130_fd_sc_hd__nand2_1 _0620_ (.A(_0084_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__o21ai_4 _0621_ (.A1(_0084_),
    .A2(_0158_),
    .B1(_0160_),
    .Y(net172));
 sky130_fd_sc_hd__a211oi_1 _0622_ (.A1(_0076_),
    .A2(_0151_),
    .B1(handle_misaligned_q),
    .C1(_0084_),
    .Y(_0161_));
 sky130_fd_sc_hd__a21o_1 _0623_ (.A1(_0084_),
    .A2(_0446_),
    .B1(_0161_),
    .X(net173));
 sky130_fd_sc_hd__nor2_1 _0624_ (.A(_0065_),
    .B(_0113_),
    .Y(net174));
 sky130_fd_sc_hd__buf_2 _0625_ (.A(_0075_),
    .X(_0162_));
 sky130_fd_sc_hd__a222oi_1 _0626_ (.A1(_0159_),
    .A2(net79),
    .B1(_0162_),
    .B2(net102),
    .C1(net88),
    .C2(_0155_),
    .Y(_0163_));
 sky130_fd_sc_hd__clkbuf_4 _0627_ (.A(_0098_),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_1 _0628_ (.A(_0164_),
    .B(net72),
    .Y(_0165_));
 sky130_fd_sc_hd__a21oi_2 _0629_ (.A1(_0433_),
    .A2(_0163_),
    .B1(_0165_),
    .Y(net175));
 sky130_fd_sc_hd__buf_2 _0630_ (.A(_0150_),
    .X(_0166_));
 sky130_fd_sc_hd__a222oi_1 _0631_ (.A1(_0166_),
    .A2(net90),
    .B1(_0162_),
    .B2(net81),
    .C1(net94),
    .C2(_0155_),
    .Y(_0167_));
 sky130_fd_sc_hd__nor2_1 _0632_ (.A(_0164_),
    .B(net73),
    .Y(_0168_));
 sky130_fd_sc_hd__a21oi_1 _0633_ (.A1(_0433_),
    .A2(_0167_),
    .B1(_0168_),
    .Y(net176));
 sky130_fd_sc_hd__a222oi_1 _0634_ (.A1(_0166_),
    .A2(net91),
    .B1(_0162_),
    .B2(net82),
    .C1(net97),
    .C2(_0155_),
    .Y(_0169_));
 sky130_fd_sc_hd__nor2_1 _0635_ (.A(_0164_),
    .B(net74),
    .Y(_0170_));
 sky130_fd_sc_hd__a21oi_1 _0636_ (.A1(_0433_),
    .A2(_0169_),
    .B1(_0170_),
    .Y(net177));
 sky130_fd_sc_hd__a222oi_1 _0637_ (.A1(_0166_),
    .A2(net92),
    .B1(_0162_),
    .B2(net84),
    .C1(net98),
    .C2(_0155_),
    .Y(_0171_));
 sky130_fd_sc_hd__nor2_1 _0638_ (.A(_0164_),
    .B(net75),
    .Y(_0172_));
 sky130_fd_sc_hd__a21oi_1 _0639_ (.A1(_0433_),
    .A2(_0171_),
    .B1(_0172_),
    .Y(net178));
 sky130_fd_sc_hd__a222oi_1 _0640_ (.A1(_0166_),
    .A2(net93),
    .B1(_0162_),
    .B2(net85),
    .C1(net99),
    .C2(_0155_),
    .Y(_0173_));
 sky130_fd_sc_hd__nor2_1 _0641_ (.A(_0164_),
    .B(net76),
    .Y(_0174_));
 sky130_fd_sc_hd__a21oi_1 _0642_ (.A1(_0433_),
    .A2(_0173_),
    .B1(_0174_),
    .Y(net179));
 sky130_fd_sc_hd__a222oi_1 _0643_ (.A1(_0166_),
    .A2(net95),
    .B1(_0162_),
    .B2(net86),
    .C1(net100),
    .C2(_0155_),
    .Y(_0175_));
 sky130_fd_sc_hd__nor2_1 _0644_ (.A(_0164_),
    .B(net77),
    .Y(_0176_));
 sky130_fd_sc_hd__a21oi_2 _0645_ (.A1(_0433_),
    .A2(_0175_),
    .B1(_0176_),
    .Y(net180));
 sky130_fd_sc_hd__a222oi_1 _0646_ (.A1(_0166_),
    .A2(net96),
    .B1(_0162_),
    .B2(net87),
    .C1(net101),
    .C2(_0155_),
    .Y(_0177_));
 sky130_fd_sc_hd__nor2_1 _0647_ (.A(_0164_),
    .B(net78),
    .Y(_0178_));
 sky130_fd_sc_hd__a21oi_1 _0648_ (.A1(_0433_),
    .A2(_0177_),
    .B1(_0178_),
    .Y(net181));
 sky130_fd_sc_hd__buf_2 _0649_ (.A(_0154_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_4 _0650_ (.A(_0075_),
    .X(_0180_));
 sky130_fd_sc_hd__a222oi_1 _0651_ (.A1(_0179_),
    .A2(net102),
    .B1(net88),
    .B2(_0180_),
    .C1(net72),
    .C2(_0159_),
    .Y(_0181_));
 sky130_fd_sc_hd__clkbuf_4 _0652_ (.A(_0097_),
    .X(_0182_));
 sky130_fd_sc_hd__nor2_1 _0653_ (.A(_0182_),
    .B(net79),
    .Y(_0183_));
 sky130_fd_sc_hd__a21oi_1 _0654_ (.A1(_0433_),
    .A2(_0181_),
    .B1(_0183_),
    .Y(net182));
 sky130_fd_sc_hd__a222oi_1 _0655_ (.A1(_0179_),
    .A2(net103),
    .B1(net89),
    .B2(_0180_),
    .C1(net83),
    .C2(_0159_),
    .Y(_0184_));
 sky130_fd_sc_hd__nor2_1 _0656_ (.A(_0182_),
    .B(net80),
    .Y(_0185_));
 sky130_fd_sc_hd__a21oi_2 _0657_ (.A1(_0433_),
    .A2(_0184_),
    .B1(_0185_),
    .Y(net183));
 sky130_fd_sc_hd__clkbuf_4 _0658_ (.A(_0098_),
    .X(_0186_));
 sky130_fd_sc_hd__a222oi_1 _0659_ (.A1(_0179_),
    .A2(net73),
    .B1(net90),
    .B2(_0180_),
    .C1(net94),
    .C2(_0159_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _0660_ (.A(_0182_),
    .B(net81),
    .Y(_0188_));
 sky130_fd_sc_hd__a21oi_1 _0661_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0188_),
    .Y(net184));
 sky130_fd_sc_hd__a222oi_1 _0662_ (.A1(_0179_),
    .A2(net74),
    .B1(net91),
    .B2(_0180_),
    .C1(net97),
    .C2(_0159_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _0663_ (.A(_0182_),
    .B(net82),
    .Y(_0190_));
 sky130_fd_sc_hd__a21oi_1 _0664_ (.A1(_0186_),
    .A2(_0189_),
    .B1(_0190_),
    .Y(net185));
 sky130_fd_sc_hd__a222oi_1 _0665_ (.A1(_0166_),
    .A2(net80),
    .B1(_0162_),
    .B2(net103),
    .C1(net89),
    .C2(_0155_),
    .Y(_0191_));
 sky130_fd_sc_hd__nor2_1 _0666_ (.A(_0182_),
    .B(net83),
    .Y(_0192_));
 sky130_fd_sc_hd__a21oi_2 _0667_ (.A1(_0186_),
    .A2(_0191_),
    .B1(_0192_),
    .Y(net186));
 sky130_fd_sc_hd__clkbuf_4 _0668_ (.A(_0075_),
    .X(_0193_));
 sky130_fd_sc_hd__a222oi_1 _0669_ (.A1(_0179_),
    .A2(net75),
    .B1(net92),
    .B2(_0193_),
    .C1(net98),
    .C2(_0159_),
    .Y(_0194_));
 sky130_fd_sc_hd__nor2_1 _0670_ (.A(_0182_),
    .B(net84),
    .Y(_0195_));
 sky130_fd_sc_hd__a21oi_1 _0671_ (.A1(_0186_),
    .A2(_0194_),
    .B1(_0195_),
    .Y(net187));
 sky130_fd_sc_hd__a222oi_1 _0672_ (.A1(_0154_),
    .A2(net76),
    .B1(net93),
    .B2(_0193_),
    .C1(net99),
    .C2(_0159_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _0673_ (.A(_0182_),
    .B(net85),
    .Y(_0197_));
 sky130_fd_sc_hd__a21oi_1 _0674_ (.A1(_0186_),
    .A2(_0196_),
    .B1(_0197_),
    .Y(net188));
 sky130_fd_sc_hd__a222oi_1 _0675_ (.A1(_0154_),
    .A2(net77),
    .B1(net95),
    .B2(_0193_),
    .C1(net100),
    .C2(_0159_),
    .Y(_0198_));
 sky130_fd_sc_hd__nor2_1 _0676_ (.A(_0182_),
    .B(net86),
    .Y(_0199_));
 sky130_fd_sc_hd__a21oi_2 _0677_ (.A1(_0186_),
    .A2(_0198_),
    .B1(_0199_),
    .Y(net189));
 sky130_fd_sc_hd__a222oi_1 _0678_ (.A1(_0154_),
    .A2(net78),
    .B1(net96),
    .B2(_0193_),
    .C1(net101),
    .C2(_0159_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _0679_ (.A(_0182_),
    .B(net87),
    .Y(_0201_));
 sky130_fd_sc_hd__a21oi_1 _0680_ (.A1(_0186_),
    .A2(_0200_),
    .B1(_0201_),
    .Y(net190));
 sky130_fd_sc_hd__a222oi_1 _0681_ (.A1(_0166_),
    .A2(net102),
    .B1(net72),
    .B2(_0193_),
    .C1(net79),
    .C2(_0155_),
    .Y(_0202_));
 sky130_fd_sc_hd__nor2_1 _0682_ (.A(_0182_),
    .B(net88),
    .Y(_0203_));
 sky130_fd_sc_hd__a21oi_1 _0683_ (.A1(_0186_),
    .A2(_0202_),
    .B1(_0203_),
    .Y(net191));
 sky130_fd_sc_hd__buf_2 _0684_ (.A(_0154_),
    .X(_0204_));
 sky130_fd_sc_hd__a222oi_1 _0685_ (.A1(_0166_),
    .A2(net103),
    .B1(net83),
    .B2(_0193_),
    .C1(net80),
    .C2(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__clkbuf_4 _0686_ (.A(_0097_),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _0687_ (.A(_0206_),
    .B(net89),
    .Y(_0207_));
 sky130_fd_sc_hd__a21oi_2 _0688_ (.A1(_0186_),
    .A2(_0205_),
    .B1(_0207_),
    .Y(net192));
 sky130_fd_sc_hd__a222oi_1 _0689_ (.A1(_0166_),
    .A2(net73),
    .B1(net94),
    .B2(_0193_),
    .C1(net81),
    .C2(_0204_),
    .Y(_0208_));
 sky130_fd_sc_hd__nor2_1 _0690_ (.A(_0206_),
    .B(net90),
    .Y(_0209_));
 sky130_fd_sc_hd__a21oi_1 _0691_ (.A1(_0186_),
    .A2(_0208_),
    .B1(_0209_),
    .Y(net193));
 sky130_fd_sc_hd__clkbuf_4 _0692_ (.A(_0098_),
    .X(_0210_));
 sky130_fd_sc_hd__buf_2 _0693_ (.A(_0150_),
    .X(_0211_));
 sky130_fd_sc_hd__a222oi_1 _0694_ (.A1(_0211_),
    .A2(net74),
    .B1(net97),
    .B2(_0193_),
    .C1(net82),
    .C2(_0204_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _0695_ (.A(_0206_),
    .B(net91),
    .Y(_0213_));
 sky130_fd_sc_hd__a21oi_1 _0696_ (.A1(_0210_),
    .A2(_0212_),
    .B1(_0213_),
    .Y(net194));
 sky130_fd_sc_hd__a222oi_1 _0697_ (.A1(_0211_),
    .A2(net75),
    .B1(net98),
    .B2(_0193_),
    .C1(net84),
    .C2(_0204_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _0698_ (.A(_0206_),
    .B(net92),
    .Y(_0215_));
 sky130_fd_sc_hd__a21oi_1 _0699_ (.A1(_0210_),
    .A2(_0214_),
    .B1(_0215_),
    .Y(net195));
 sky130_fd_sc_hd__a222oi_1 _0700_ (.A1(_0211_),
    .A2(net76),
    .B1(net99),
    .B2(_0193_),
    .C1(net85),
    .C2(_0204_),
    .Y(_0216_));
 sky130_fd_sc_hd__nor2_1 _0701_ (.A(_0206_),
    .B(net93),
    .Y(_0217_));
 sky130_fd_sc_hd__a21oi_1 _0702_ (.A1(_0210_),
    .A2(_0216_),
    .B1(_0217_),
    .Y(net196));
 sky130_fd_sc_hd__a222oi_1 _0703_ (.A1(_0211_),
    .A2(net81),
    .B1(_0162_),
    .B2(net73),
    .C1(net90),
    .C2(_0204_),
    .Y(_0218_));
 sky130_fd_sc_hd__nor2_1 _0704_ (.A(_0206_),
    .B(net94),
    .Y(_0219_));
 sky130_fd_sc_hd__a21oi_1 _0705_ (.A1(_0210_),
    .A2(_0218_),
    .B1(_0219_),
    .Y(net197));
 sky130_fd_sc_hd__a222oi_1 _0706_ (.A1(_0211_),
    .A2(net77),
    .B1(net100),
    .B2(_0075_),
    .C1(net86),
    .C2(_0204_),
    .Y(_0220_));
 sky130_fd_sc_hd__nor2_1 _0707_ (.A(_0206_),
    .B(net95),
    .Y(_0221_));
 sky130_fd_sc_hd__a21oi_2 _0708_ (.A1(_0210_),
    .A2(_0220_),
    .B1(_0221_),
    .Y(net198));
 sky130_fd_sc_hd__a222oi_1 _0709_ (.A1(_0211_),
    .A2(net78),
    .B1(net101),
    .B2(_0075_),
    .C1(net87),
    .C2(_0204_),
    .Y(_0222_));
 sky130_fd_sc_hd__nor2_1 _0710_ (.A(_0206_),
    .B(net96),
    .Y(_0223_));
 sky130_fd_sc_hd__a21oi_4 _0711_ (.A1(_0210_),
    .A2(_0222_),
    .B1(_0223_),
    .Y(net199));
 sky130_fd_sc_hd__a222oi_1 _0712_ (.A1(_0211_),
    .A2(net82),
    .B1(_0162_),
    .B2(net74),
    .C1(net91),
    .C2(_0204_),
    .Y(_0224_));
 sky130_fd_sc_hd__nor2_1 _0713_ (.A(_0206_),
    .B(net97),
    .Y(_0225_));
 sky130_fd_sc_hd__a21oi_1 _0714_ (.A1(_0210_),
    .A2(_0224_),
    .B1(_0225_),
    .Y(net200));
 sky130_fd_sc_hd__a222oi_1 _0715_ (.A1(_0211_),
    .A2(net84),
    .B1(_0180_),
    .B2(net75),
    .C1(net92),
    .C2(_0204_),
    .Y(_0226_));
 sky130_fd_sc_hd__nor2_1 _0716_ (.A(_0206_),
    .B(net98),
    .Y(_0227_));
 sky130_fd_sc_hd__a21oi_1 _0717_ (.A1(_0210_),
    .A2(_0226_),
    .B1(_0227_),
    .Y(net201));
 sky130_fd_sc_hd__a222oi_1 _0718_ (.A1(_0211_),
    .A2(net85),
    .B1(_0180_),
    .B2(net76),
    .C1(net93),
    .C2(_0179_),
    .Y(_0228_));
 sky130_fd_sc_hd__nor2_1 _0719_ (.A(_0098_),
    .B(net99),
    .Y(_0229_));
 sky130_fd_sc_hd__a21oi_1 _0720_ (.A1(_0210_),
    .A2(_0228_),
    .B1(_0229_),
    .Y(net202));
 sky130_fd_sc_hd__a222oi_1 _0721_ (.A1(_0211_),
    .A2(net86),
    .B1(_0180_),
    .B2(net77),
    .C1(net95),
    .C2(_0179_),
    .Y(_0230_));
 sky130_fd_sc_hd__nor2_1 _0722_ (.A(_0098_),
    .B(net100),
    .Y(_0231_));
 sky130_fd_sc_hd__a21oi_2 _0723_ (.A1(_0210_),
    .A2(_0230_),
    .B1(_0231_),
    .Y(net203));
 sky130_fd_sc_hd__a222oi_1 _0724_ (.A1(_0150_),
    .A2(net87),
    .B1(_0180_),
    .B2(net78),
    .C1(net96),
    .C2(_0179_),
    .Y(_0232_));
 sky130_fd_sc_hd__nor2_1 _0725_ (.A(_0098_),
    .B(net101),
    .Y(_0233_));
 sky130_fd_sc_hd__a21oi_1 _0726_ (.A1(_0164_),
    .A2(_0232_),
    .B1(_0233_),
    .Y(net204));
 sky130_fd_sc_hd__a222oi_1 _0727_ (.A1(_0150_),
    .A2(net88),
    .B1(_0180_),
    .B2(net79),
    .C1(net72),
    .C2(_0179_),
    .Y(_0234_));
 sky130_fd_sc_hd__nor2_1 _0728_ (.A(_0098_),
    .B(net102),
    .Y(_0235_));
 sky130_fd_sc_hd__a21oi_1 _0729_ (.A1(_0164_),
    .A2(_0234_),
    .B1(_0235_),
    .Y(net205));
 sky130_fd_sc_hd__a222oi_1 _0730_ (.A1(_0150_),
    .A2(net89),
    .B1(_0180_),
    .B2(net80),
    .C1(net83),
    .C2(_0179_),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _0731_ (.A(_0098_),
    .B(net103),
    .Y(_0237_));
 sky130_fd_sc_hd__a21oi_4 _0732_ (.A1(_0164_),
    .A2(_0236_),
    .B1(_0237_),
    .Y(net206));
 sky130_fd_sc_hd__nor2_1 _0733_ (.A(net139),
    .B(_0112_),
    .Y(net243));
 sky130_fd_sc_hd__o21a_1 _0734_ (.A1(net33),
    .A2(lsu_err_q),
    .B1(net68),
    .X(_0238_));
 sky130_fd_sc_hd__nor2_1 _0735_ (.A(_0069_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nor3_1 _0736_ (.A(data_we_q),
    .B(net139),
    .C(_0239_),
    .Y(net208));
 sky130_fd_sc_hd__nand2b_1 _0737_ (.A_N(_0135_),
    .B(net36),
    .Y(_0240_));
 sky130_fd_sc_hd__mux2i_1 _0738_ (.A0(\rdata_q[24] ),
    .A1(net52),
    .S(_0110_),
    .Y(_0241_));
 sky130_fd_sc_hd__buf_4 _0739_ (.A(_0137_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_8 _0740_ (.A(_0242_),
    .B(_0135_),
    .Y(_0243_));
 sky130_fd_sc_hd__nor2_4 _0741_ (.A(_0109_),
    .B(\data_type_q[1] ),
    .Y(_0244_));
 sky130_fd_sc_hd__buf_4 _0742_ (.A(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_4 _0743_ (.A(_0133_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2b_1 _0744_ (.A_N(_0246_),
    .B(net43),
    .Y(_0247_));
 sky130_fd_sc_hd__buf_4 _0745_ (.A(_0134_),
    .X(_0248_));
 sky130_fd_sc_hd__a21oi_1 _0746_ (.A1(_0248_),
    .A2(net66),
    .B1(_0138_),
    .Y(_0249_));
 sky130_fd_sc_hd__a21oi_1 _0747_ (.A1(_0242_),
    .A2(_0247_),
    .B1(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__nor2b_1 _0748_ (.A(_0136_),
    .B_N(_0132_),
    .Y(_0251_));
 sky130_fd_sc_hd__buf_4 _0749_ (.A(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2b_1 _0750_ (.A(_0132_),
    .B_N(_0136_),
    .Y(_0253_));
 sky130_fd_sc_hd__buf_4 _0751_ (.A(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__or2_0 _0752_ (.A(\data_type_q[0] ),
    .B(\data_type_q[1] ),
    .X(_0255_));
 sky130_fd_sc_hd__clkbuf_4 _0753_ (.A(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__a221o_1 _0754_ (.A1(\rdata_q[8] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[16] ),
    .C1(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__o21ai_0 _0755_ (.A1(_0245_),
    .A2(_0250_),
    .B1(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__o221ai_2 _0756_ (.A1(_0139_),
    .A2(_0240_),
    .B1(_0241_),
    .B2(_0243_),
    .C1(_0258_),
    .Y(net209));
 sky130_fd_sc_hd__clkbuf_4 _0757_ (.A(_0136_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _0758_ (.A(_0246_),
    .B(net45),
    .Y(_0260_));
 sky130_fd_sc_hd__clkbuf_4 _0759_ (.A(_0136_),
    .X(_0261_));
 sky130_fd_sc_hd__nand3b_1 _0760_ (.A_N(_0134_),
    .B(net54),
    .C(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__o21ai_0 _0761_ (.A1(_0259_),
    .A2(_0260_),
    .B1(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__clkbuf_4 _0762_ (.A(_0133_),
    .X(_0264_));
 sky130_fd_sc_hd__buf_4 _0763_ (.A(\data_type_q[0] ),
    .X(_0265_));
 sky130_fd_sc_hd__nand2b_1 _0764_ (.A_N(_0265_),
    .B(\rdata_q[18] ),
    .Y(_0266_));
 sky130_fd_sc_hd__a21oi_1 _0765_ (.A1(_0264_),
    .A2(_0266_),
    .B1(_0138_),
    .Y(_0267_));
 sky130_fd_sc_hd__and2_0 _0766_ (.A(\rdata_offset_q[1] ),
    .B(_0132_),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_4 _0767_ (.A(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_4 _0768_ (.A(_0133_),
    .B(_0265_),
    .Y(_0270_));
 sky130_fd_sc_hd__a22o_1 _0769_ (.A1(net58),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[26] ),
    .X(_0271_));
 sky130_fd_sc_hd__a211oi_1 _0770_ (.A1(_0109_),
    .A2(_0263_),
    .B1(_0267_),
    .C1(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__or2_0 _0771_ (.A(\rdata_offset_q[1] ),
    .B(\rdata_offset_q[0] ),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_4 _0772_ (.A(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_1 _0773_ (.A(net37),
    .B(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_1 _0774_ (.A(data_sign_ext_q),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2b_1 _0775_ (.A_N(\rdata_offset_q[0] ),
    .B(net51),
    .Y(_0277_));
 sky130_fd_sc_hd__a21boi_1 _0776_ (.A1(net42),
    .A2(data_sign_ext_q),
    .B1_N(_0132_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand4_1 _0777_ (.A(_0136_),
    .B(_0132_),
    .C(net60),
    .D(data_sign_ext_q),
    .Y(_0279_));
 sky130_fd_sc_hd__o221ai_4 _0778_ (.A1(_0276_),
    .A2(_0277_),
    .B1(_0278_),
    .B2(_0136_),
    .C1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21o_1 _0779_ (.A1(net65),
    .A2(data_sign_ext_q),
    .B1(_0274_),
    .X(_0281_));
 sky130_fd_sc_hd__nand3_4 _0780_ (.A(_0111_),
    .B(_0280_),
    .C(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__o31ai_2 _0781_ (.A1(_0111_),
    .A2(_0272_),
    .A3(_0275_),
    .B1(_0282_),
    .Y(net210));
 sky130_fd_sc_hd__nand2_1 _0782_ (.A(_0246_),
    .B(net46),
    .Y(_0283_));
 sky130_fd_sc_hd__nand3b_1 _0783_ (.A_N(_0133_),
    .B(net55),
    .C(_0261_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_0 _0784_ (.A1(_0259_),
    .A2(_0283_),
    .B1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand2b_1 _0785_ (.A_N(_0265_),
    .B(\rdata_q[19] ),
    .Y(_0286_));
 sky130_fd_sc_hd__a21oi_1 _0786_ (.A1(_0264_),
    .A2(_0286_),
    .B1(_0259_),
    .Y(_0287_));
 sky130_fd_sc_hd__a22o_1 _0787_ (.A1(net61),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[27] ),
    .X(_0288_));
 sky130_fd_sc_hd__a211oi_1 _0788_ (.A1(_0109_),
    .A2(_0285_),
    .B1(_0287_),
    .C1(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__nor2_1 _0789_ (.A(net38),
    .B(_0274_),
    .Y(_0290_));
 sky130_fd_sc_hd__o31ai_2 _0790_ (.A1(_0111_),
    .A2(_0289_),
    .A3(_0290_),
    .B1(_0282_),
    .Y(net211));
 sky130_fd_sc_hd__nand2_1 _0791_ (.A(_0246_),
    .B(net48),
    .Y(_0291_));
 sky130_fd_sc_hd__nand3b_1 _0792_ (.A_N(_0133_),
    .B(net56),
    .C(_0261_),
    .Y(_0292_));
 sky130_fd_sc_hd__o21ai_0 _0793_ (.A1(_0259_),
    .A2(_0291_),
    .B1(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2b_1 _0794_ (.A_N(_0265_),
    .B(\rdata_q[20] ),
    .Y(_0294_));
 sky130_fd_sc_hd__a21oi_1 _0795_ (.A1(_0264_),
    .A2(_0294_),
    .B1(_0259_),
    .Y(_0295_));
 sky130_fd_sc_hd__a22o_1 _0796_ (.A1(net62),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[28] ),
    .X(_0296_));
 sky130_fd_sc_hd__a211oi_1 _0797_ (.A1(_0109_),
    .A2(_0293_),
    .B1(_0295_),
    .C1(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _0798_ (.A(net39),
    .B(_0274_),
    .Y(_0298_));
 sky130_fd_sc_hd__o31ai_2 _0799_ (.A1(_0111_),
    .A2(_0297_),
    .A3(_0298_),
    .B1(_0282_),
    .Y(net212));
 sky130_fd_sc_hd__nand2_1 _0800_ (.A(_0246_),
    .B(net49),
    .Y(_0299_));
 sky130_fd_sc_hd__nand3b_1 _0801_ (.A_N(_0133_),
    .B(net57),
    .C(_0261_),
    .Y(_0300_));
 sky130_fd_sc_hd__o21ai_0 _0802_ (.A1(_0261_),
    .A2(_0299_),
    .B1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand2b_1 _0803_ (.A_N(_0265_),
    .B(\rdata_q[21] ),
    .Y(_0302_));
 sky130_fd_sc_hd__a21oi_1 _0804_ (.A1(_0264_),
    .A2(_0302_),
    .B1(_0259_),
    .Y(_0303_));
 sky130_fd_sc_hd__a22o_1 _0805_ (.A1(net63),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[29] ),
    .X(_0304_));
 sky130_fd_sc_hd__a211oi_1 _0806_ (.A1(_0109_),
    .A2(_0301_),
    .B1(_0303_),
    .C1(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_1 _0807_ (.A(net40),
    .B(_0274_),
    .Y(_0306_));
 sky130_fd_sc_hd__o31ai_1 _0808_ (.A1(_0111_),
    .A2(_0305_),
    .A3(_0306_),
    .B1(_0282_),
    .Y(net213));
 sky130_fd_sc_hd__nand2_1 _0809_ (.A(_0246_),
    .B(net50),
    .Y(_0307_));
 sky130_fd_sc_hd__nand3b_1 _0810_ (.A_N(_0133_),
    .B(net59),
    .C(_0261_),
    .Y(_0308_));
 sky130_fd_sc_hd__o21ai_0 _0811_ (.A1(_0261_),
    .A2(_0307_),
    .B1(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__nand2b_1 _0812_ (.A_N(_0265_),
    .B(\rdata_q[22] ),
    .Y(_0310_));
 sky130_fd_sc_hd__a21oi_1 _0813_ (.A1(_0264_),
    .A2(_0310_),
    .B1(_0259_),
    .Y(_0311_));
 sky130_fd_sc_hd__a22o_1 _0814_ (.A1(net64),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[30] ),
    .X(_0312_));
 sky130_fd_sc_hd__a211oi_1 _0815_ (.A1(_0109_),
    .A2(_0309_),
    .B1(_0311_),
    .C1(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__nor2_1 _0816_ (.A(net41),
    .B(_0274_),
    .Y(_0314_));
 sky130_fd_sc_hd__o31ai_1 _0817_ (.A1(_0111_),
    .A2(_0313_),
    .A3(_0314_),
    .B1(_0282_),
    .Y(net214));
 sky130_fd_sc_hd__nor2b_1 _0818_ (.A(_0132_),
    .B_N(net60),
    .Y(_0315_));
 sky130_fd_sc_hd__a22o_1 _0819_ (.A1(net51),
    .A2(_0252_),
    .B1(_0315_),
    .B2(_0137_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2b_1 _0820_ (.A_N(_0265_),
    .B(\rdata_q[23] ),
    .Y(_0317_));
 sky130_fd_sc_hd__a21oi_1 _0821_ (.A1(_0264_),
    .A2(_0317_),
    .B1(_0259_),
    .Y(_0318_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(net65),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[31] ),
    .X(_0319_));
 sky130_fd_sc_hd__a211oi_1 _0823_ (.A1(_0109_),
    .A2(_0316_),
    .B1(_0318_),
    .C1(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__nor3_1 _0824_ (.A(_0136_),
    .B(_0132_),
    .C(net42),
    .Y(_0321_));
 sky130_fd_sc_hd__o31ai_2 _0825_ (.A1(_0111_),
    .A2(_0320_),
    .A3(_0321_),
    .B1(_0282_),
    .Y(net215));
 sky130_fd_sc_hd__clkbuf_8 _0826_ (.A(_0136_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2i_1 _0827_ (.A0(net60),
    .A1(net65),
    .S(_0132_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor3b_1 _0828_ (.A(_0136_),
    .B(net51),
    .C_N(_0132_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_1 _0829_ (.A1(_0322_),
    .A2(_0323_),
    .B1(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2_1 _0830_ (.A(_0265_),
    .B(data_sign_ext_q),
    .Y(_0326_));
 sky130_fd_sc_hd__nor3_1 _0831_ (.A(\data_type_q[1] ),
    .B(_0321_),
    .C(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__a32oi_4 _0832_ (.A1(_0110_),
    .A2(_0280_),
    .A3(_0281_),
    .B1(_0325_),
    .B2(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__buf_4 _0833_ (.A(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_4 _0834_ (.A(_0244_),
    .X(_0330_));
 sky130_fd_sc_hd__buf_4 _0835_ (.A(_0134_),
    .X(_0331_));
 sky130_fd_sc_hd__mux4_1 _0836_ (.A0(net43),
    .A1(net36),
    .A2(\rdata_q[24] ),
    .A3(net66),
    .S0(_0137_),
    .S1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _0837_ (.A(_0330_),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand2_1 _0838_ (.A(_0329_),
    .B(_0333_),
    .Y(net216));
 sky130_fd_sc_hd__mux4_1 _0839_ (.A0(net44),
    .A1(net47),
    .A2(\rdata_q[25] ),
    .A3(net67),
    .S0(_0137_),
    .S1(_0331_),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _0840_ (.A(_0330_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _0841_ (.A(_0329_),
    .B(_0335_),
    .Y(net217));
 sky130_fd_sc_hd__mux4_1 _0842_ (.A0(net45),
    .A1(net58),
    .A2(\rdata_q[26] ),
    .A3(net37),
    .S0(_0137_),
    .S1(_0331_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_1 _0843_ (.A(_0330_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _0844_ (.A(_0329_),
    .B(_0337_),
    .Y(net218));
 sky130_fd_sc_hd__mux4_1 _0845_ (.A0(net46),
    .A1(net61),
    .A2(\rdata_q[27] ),
    .A3(net38),
    .S0(_0137_),
    .S1(_0331_),
    .X(_0338_));
 sky130_fd_sc_hd__nand2_1 _0846_ (.A(_0330_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _0847_ (.A(_0329_),
    .B(_0339_),
    .Y(net219));
 sky130_fd_sc_hd__nand2b_1 _0848_ (.A_N(_0135_),
    .B(net47),
    .Y(_0340_));
 sky130_fd_sc_hd__mux2i_2 _0849_ (.A0(\rdata_q[25] ),
    .A1(net53),
    .S(_0110_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand2b_1 _0850_ (.A_N(_0134_),
    .B(net44),
    .Y(_0342_));
 sky130_fd_sc_hd__a21oi_1 _0851_ (.A1(_0248_),
    .A2(net67),
    .B1(_0138_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21oi_1 _0852_ (.A1(_0242_),
    .A2(_0342_),
    .B1(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__a221o_1 _0853_ (.A1(\rdata_q[9] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[17] ),
    .C1(_0256_),
    .X(_0345_));
 sky130_fd_sc_hd__o21ai_2 _0854_ (.A1(_0245_),
    .A2(_0344_),
    .B1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__o221ai_4 _0855_ (.A1(_0139_),
    .A2(_0340_),
    .B1(_0341_),
    .B2(_0243_),
    .C1(_0346_),
    .Y(net220));
 sky130_fd_sc_hd__mux4_1 _0856_ (.A0(net48),
    .A1(net62),
    .A2(\rdata_q[28] ),
    .A3(net39),
    .S0(_0137_),
    .S1(_0331_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_1 _0857_ (.A(_0330_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _0858_ (.A(_0329_),
    .B(_0348_),
    .Y(net221));
 sky130_fd_sc_hd__mux4_1 _0859_ (.A0(net49),
    .A1(net63),
    .A2(\rdata_q[29] ),
    .A3(net40),
    .S0(_0137_),
    .S1(_0331_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _0860_ (.A(_0330_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _0861_ (.A(_0329_),
    .B(_0350_),
    .Y(net222));
 sky130_fd_sc_hd__mux4_1 _0862_ (.A0(net50),
    .A1(net64),
    .A2(\rdata_q[30] ),
    .A3(net41),
    .S0(_0322_),
    .S1(_0331_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _0863_ (.A(_0330_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _0864_ (.A(_0329_),
    .B(_0352_),
    .Y(net223));
 sky130_fd_sc_hd__mux4_1 _0865_ (.A0(net51),
    .A1(net65),
    .A2(\rdata_q[31] ),
    .A3(net42),
    .S0(_0322_),
    .S1(_0331_),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_1 _0866_ (.A(_0330_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _0867_ (.A(_0329_),
    .B(_0354_),
    .Y(net224));
 sky130_fd_sc_hd__mux4_1 _0868_ (.A0(net52),
    .A1(net66),
    .A2(net36),
    .A3(net43),
    .S0(_0322_),
    .S1(_0331_),
    .X(_0355_));
 sky130_fd_sc_hd__nand2_1 _0869_ (.A(_0330_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _0870_ (.A(_0329_),
    .B(_0356_),
    .Y(net225));
 sky130_fd_sc_hd__mux4_1 _0871_ (.A0(net53),
    .A1(net67),
    .A2(net47),
    .A3(net44),
    .S0(_0322_),
    .S1(_0248_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_1 _0872_ (.A(_0330_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _0873_ (.A(_0329_),
    .B(_0358_),
    .Y(net226));
 sky130_fd_sc_hd__mux4_1 _0874_ (.A0(net54),
    .A1(net37),
    .A2(net58),
    .A3(net45),
    .S0(_0322_),
    .S1(_0248_),
    .X(_0359_));
 sky130_fd_sc_hd__nand2_1 _0875_ (.A(_0245_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _0876_ (.A(_0328_),
    .B(_0360_),
    .Y(net227));
 sky130_fd_sc_hd__mux4_1 _0877_ (.A0(net55),
    .A1(net38),
    .A2(net61),
    .A3(net46),
    .S0(_0322_),
    .S1(_0248_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _0878_ (.A(_0245_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2_1 _0879_ (.A(_0328_),
    .B(_0362_),
    .Y(net228));
 sky130_fd_sc_hd__mux4_1 _0880_ (.A0(net56),
    .A1(net39),
    .A2(net62),
    .A3(net48),
    .S0(_0322_),
    .S1(_0248_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _0881_ (.A(_0245_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2_1 _0882_ (.A(_0328_),
    .B(_0364_),
    .Y(net229));
 sky130_fd_sc_hd__mux4_1 _0883_ (.A0(net57),
    .A1(net40),
    .A2(net63),
    .A3(net49),
    .S0(_0322_),
    .S1(_0248_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _0884_ (.A(_0245_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _0885_ (.A(_0328_),
    .B(_0366_),
    .Y(net230));
 sky130_fd_sc_hd__nand2b_1 _0886_ (.A_N(_0135_),
    .B(net58),
    .Y(_0367_));
 sky130_fd_sc_hd__mux2i_2 _0887_ (.A0(\rdata_q[26] ),
    .A1(net54),
    .S(_0110_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2b_1 _0888_ (.A_N(_0134_),
    .B(net45),
    .Y(_0369_));
 sky130_fd_sc_hd__a21oi_1 _0889_ (.A1(_0248_),
    .A2(net37),
    .B1(_0138_),
    .Y(_0370_));
 sky130_fd_sc_hd__a21oi_1 _0890_ (.A1(_0242_),
    .A2(_0369_),
    .B1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__a221o_1 _0891_ (.A1(\rdata_q[10] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[18] ),
    .C1(_0256_),
    .X(_0372_));
 sky130_fd_sc_hd__o21ai_1 _0892_ (.A1(_0245_),
    .A2(_0371_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__o221ai_4 _0893_ (.A1(_0139_),
    .A2(_0367_),
    .B1(_0368_),
    .B2(_0243_),
    .C1(_0373_),
    .Y(net231));
 sky130_fd_sc_hd__mux4_1 _0894_ (.A0(net59),
    .A1(net41),
    .A2(net64),
    .A3(net50),
    .S0(_0322_),
    .S1(_0248_),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _0895_ (.A(_0245_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _0896_ (.A(_0328_),
    .B(_0375_),
    .Y(net232));
 sky130_fd_sc_hd__mux2i_1 _0897_ (.A0(net42),
    .A1(net51),
    .S(_0135_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _0898_ (.A(_0139_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2b_1 _0899_ (.A_N(_0242_),
    .B(_0323_),
    .Y(_0378_));
 sky130_fd_sc_hd__nand3_1 _0900_ (.A(_0245_),
    .B(_0377_),
    .C(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _0901_ (.A(_0328_),
    .B(_0379_),
    .Y(net233));
 sky130_fd_sc_hd__nand2b_1 _0902_ (.A_N(_0135_),
    .B(net61),
    .Y(_0380_));
 sky130_fd_sc_hd__mux2i_2 _0903_ (.A0(\rdata_q[27] ),
    .A1(net55),
    .S(_0110_),
    .Y(_0381_));
 sky130_fd_sc_hd__nand2b_1 _0904_ (.A_N(_0134_),
    .B(net46),
    .Y(_0382_));
 sky130_fd_sc_hd__a21oi_1 _0905_ (.A1(_0248_),
    .A2(net38),
    .B1(_0138_),
    .Y(_0383_));
 sky130_fd_sc_hd__a21oi_1 _0906_ (.A1(_0242_),
    .A2(_0382_),
    .B1(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__a221o_1 _0907_ (.A1(\rdata_q[11] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[19] ),
    .C1(_0256_),
    .X(_0385_));
 sky130_fd_sc_hd__o21ai_1 _0908_ (.A1(_0245_),
    .A2(_0384_),
    .B1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__o221ai_4 _0909_ (.A1(_0139_),
    .A2(_0380_),
    .B1(_0381_),
    .B2(_0243_),
    .C1(_0386_),
    .Y(net234));
 sky130_fd_sc_hd__nand2b_1 _0910_ (.A_N(_0135_),
    .B(net62),
    .Y(_0387_));
 sky130_fd_sc_hd__mux2i_1 _0911_ (.A0(\rdata_q[28] ),
    .A1(net56),
    .S(_0110_),
    .Y(_0388_));
 sky130_fd_sc_hd__nand2b_1 _0912_ (.A_N(_0134_),
    .B(net48),
    .Y(_0389_));
 sky130_fd_sc_hd__a21oi_1 _0913_ (.A1(_0264_),
    .A2(net39),
    .B1(_0138_),
    .Y(_0390_));
 sky130_fd_sc_hd__a21oi_1 _0914_ (.A1(_0242_),
    .A2(_0389_),
    .B1(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a221o_1 _0915_ (.A1(\rdata_q[12] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[20] ),
    .C1(_0256_),
    .X(_0392_));
 sky130_fd_sc_hd__o21ai_0 _0916_ (.A1(_0244_),
    .A2(_0391_),
    .B1(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__o221ai_2 _0917_ (.A1(_0139_),
    .A2(_0387_),
    .B1(_0388_),
    .B2(_0243_),
    .C1(_0393_),
    .Y(net235));
 sky130_fd_sc_hd__nand2b_1 _0918_ (.A_N(_0135_),
    .B(net63),
    .Y(_0394_));
 sky130_fd_sc_hd__mux2i_1 _0919_ (.A0(\rdata_q[29] ),
    .A1(net57),
    .S(_0110_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2b_1 _0920_ (.A_N(_0134_),
    .B(net49),
    .Y(_0396_));
 sky130_fd_sc_hd__a21oi_1 _0921_ (.A1(_0264_),
    .A2(net40),
    .B1(_0138_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21oi_1 _0922_ (.A1(_0242_),
    .A2(_0396_),
    .B1(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__a221o_1 _0923_ (.A1(\rdata_q[13] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[21] ),
    .C1(_0256_),
    .X(_0399_));
 sky130_fd_sc_hd__o21ai_0 _0924_ (.A1(_0244_),
    .A2(_0398_),
    .B1(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__o221ai_2 _0925_ (.A1(_0139_),
    .A2(_0394_),
    .B1(_0395_),
    .B2(_0243_),
    .C1(_0400_),
    .Y(net236));
 sky130_fd_sc_hd__nand2b_1 _0926_ (.A_N(_0135_),
    .B(net64),
    .Y(_0401_));
 sky130_fd_sc_hd__mux2i_1 _0927_ (.A0(\rdata_q[30] ),
    .A1(net59),
    .S(_0110_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2b_1 _0928_ (.A_N(_0134_),
    .B(net50),
    .Y(_0403_));
 sky130_fd_sc_hd__a21oi_1 _0929_ (.A1(_0264_),
    .A2(net41),
    .B1(_0138_),
    .Y(_0404_));
 sky130_fd_sc_hd__a21oi_1 _0930_ (.A1(_0242_),
    .A2(_0403_),
    .B1(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__a221o_1 _0931_ (.A1(\rdata_q[14] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[22] ),
    .C1(_0256_),
    .X(_0406_));
 sky130_fd_sc_hd__o21ai_0 _0932_ (.A1(_0244_),
    .A2(_0405_),
    .B1(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__o221ai_2 _0933_ (.A1(_0139_),
    .A2(_0401_),
    .B1(_0402_),
    .B2(_0243_),
    .C1(_0407_),
    .Y(net237));
 sky130_fd_sc_hd__nand2b_1 _0934_ (.A_N(_0331_),
    .B(net65),
    .Y(_0408_));
 sky130_fd_sc_hd__mux2i_2 _0935_ (.A0(\rdata_q[31] ),
    .A1(net60),
    .S(_0110_),
    .Y(_0409_));
 sky130_fd_sc_hd__a21oi_1 _0936_ (.A1(_0264_),
    .A2(net42),
    .B1(_0138_),
    .Y(_0410_));
 sky130_fd_sc_hd__a21oi_1 _0937_ (.A1(_0242_),
    .A2(_0277_),
    .B1(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__a221o_1 _0938_ (.A1(\rdata_q[15] ),
    .A2(_0252_),
    .B1(_0254_),
    .B2(\rdata_q[23] ),
    .C1(_0256_),
    .X(_0412_));
 sky130_fd_sc_hd__o21ai_1 _0939_ (.A1(_0244_),
    .A2(_0411_),
    .B1(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__o221ai_4 _0940_ (.A1(_0139_),
    .A2(_0408_),
    .B1(_0409_),
    .B2(_0243_),
    .C1(_0413_),
    .Y(net238));
 sky130_fd_sc_hd__nand2_1 _0941_ (.A(_0246_),
    .B(net43),
    .Y(_0414_));
 sky130_fd_sc_hd__nand3b_1 _0942_ (.A_N(_0133_),
    .B(net52),
    .C(_0261_),
    .Y(_0415_));
 sky130_fd_sc_hd__o21ai_0 _0943_ (.A1(_0261_),
    .A2(_0414_),
    .B1(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__nand2b_1 _0944_ (.A_N(_0265_),
    .B(\rdata_q[16] ),
    .Y(_0417_));
 sky130_fd_sc_hd__a21oi_1 _0945_ (.A1(_0246_),
    .A2(_0417_),
    .B1(_0259_),
    .Y(_0418_));
 sky130_fd_sc_hd__a22o_1 _0946_ (.A1(net36),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[24] ),
    .X(_0419_));
 sky130_fd_sc_hd__a211oi_1 _0947_ (.A1(_0109_),
    .A2(_0416_),
    .B1(_0418_),
    .C1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__nor2_1 _0948_ (.A(net66),
    .B(_0274_),
    .Y(_0421_));
 sky130_fd_sc_hd__o31ai_1 _0949_ (.A1(_0111_),
    .A2(_0420_),
    .A3(_0421_),
    .B1(_0282_),
    .Y(net239));
 sky130_fd_sc_hd__nand2_1 _0950_ (.A(_0246_),
    .B(net44),
    .Y(_0422_));
 sky130_fd_sc_hd__nand3b_1 _0951_ (.A_N(_0133_),
    .B(net53),
    .C(_0137_),
    .Y(_0423_));
 sky130_fd_sc_hd__o21ai_0 _0952_ (.A1(_0261_),
    .A2(_0422_),
    .B1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2b_1 _0953_ (.A_N(_0265_),
    .B(\rdata_q[17] ),
    .Y(_0425_));
 sky130_fd_sc_hd__a21oi_1 _0954_ (.A1(_0246_),
    .A2(_0425_),
    .B1(_0259_),
    .Y(_0426_));
 sky130_fd_sc_hd__a22o_1 _0955_ (.A1(net47),
    .A2(_0269_),
    .B1(_0270_),
    .B2(\rdata_q[25] ),
    .X(_0427_));
 sky130_fd_sc_hd__a211oi_1 _0956_ (.A1(_0109_),
    .A2(_0424_),
    .B1(_0426_),
    .C1(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__nor2_1 _0957_ (.A(net67),
    .B(_0274_),
    .Y(_0429_));
 sky130_fd_sc_hd__o31ai_2 _0958_ (.A1(_0111_),
    .A2(_0428_),
    .A3(_0429_),
    .B1(_0282_),
    .Y(net240));
 sky130_fd_sc_hd__or3_1 _0959_ (.A(_0069_),
    .B(lsu_err_q),
    .C(_0099_),
    .X(_0430_));
 sky130_fd_sc_hd__nor3_1 _0960_ (.A(data_we_q),
    .B(net139),
    .C(_0430_),
    .Y(net241));
 sky130_fd_sc_hd__nor2_1 _0961_ (.A(net69),
    .B(net139),
    .Y(_0431_));
 sky130_fd_sc_hd__nor4_1 _0962_ (.A(\ls_fsm_ns[1] ),
    .B(\ls_fsm_ns[0] ),
    .C(\ls_fsm_ns[2] ),
    .D(_0431_),
    .Y(net242));
 sky130_fd_sc_hd__nor2b_1 _0963_ (.A(net104),
    .B_N(_0079_),
    .Y(net244));
 sky130_fd_sc_hd__and2_1 _0964_ (.A(net104),
    .B(_0079_),
    .X(net245));
 sky130_fd_sc_hd__nor3b_2 _0965_ (.A(_0239_),
    .B(net139),
    .C_N(data_we_q),
    .Y(net246));
 sky130_fd_sc_hd__ha_1 _0966_ (.A(_0432_),
    .B(_0433_),
    .COUT(_0434_),
    .SUM(_0435_));
 sky130_fd_sc_hd__ha_1 _0967_ (.A(_0436_),
    .B(_0437_),
    .COUT(_0438_),
    .SUM(_0439_));
 sky130_fd_sc_hd__ha_1 _0968_ (.A(_0436_),
    .B(net12),
    .COUT(_0440_),
    .SUM(_0441_));
 sky130_fd_sc_hd__ha_1 _0969_ (.A(net1),
    .B(_0437_),
    .COUT(_0442_),
    .SUM(_0443_));
 sky130_fd_sc_hd__ha_1 _0970_ (.A(net1),
    .B(net12),
    .COUT(_0444_),
    .SUM(_0445_));
 sky130_fd_sc_hd__ha_1 _0971_ (.A(net1),
    .B(net12),
    .COUT(_0446_),
    .SUM(_0447_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__buf_4 _0973_ (.A(net247),
    .X(data_addr_o[0]));
 sky130_fd_sc_hd__buf_4 _0974_ (.A(net248),
    .X(data_addr_o[1]));
 sky130_fd_sc_hd__clkbuf_1 _0975_ (.A(net23),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _0976_ (.A(net26),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(net27),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 _0978_ (.A(net28),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _0979_ (.A(net29),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(net30),
    .X(net167));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0981_ (.A(net31),
    .X(net168));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0982_ (.A(net32),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(net2),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _0984_ (.A(net3),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(net4),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _0986_ (.A(net5),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 _0987_ (.A(net6),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _0988_ (.A(net7),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(net8),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _0990_ (.A(net9),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _0991_ (.A(net10),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(net11),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _0993_ (.A(net13),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(net14),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _0995_ (.A(net15),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0996_ (.A(net16),
    .X(net153));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0997_ (.A(net17),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(net18),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(net19),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(net20),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(net21),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _1002_ (.A(net22),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(net24),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 _1004_ (.A(net25),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _1005_ (.A(net104),
    .X(net207));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[0]$_DFFE_PN0P_  (.D(_0000_),
    .Q(net107),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[10]$_DFFE_PN0P_  (.D(_0001_),
    .Q(net108),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[11]$_DFFE_PN0P_  (.D(_0002_),
    .Q(net109),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[12]$_DFFE_PN0P_  (.D(_0003_),
    .Q(net110),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[13]$_DFFE_PN0P_  (.D(_0004_),
    .Q(net111),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[14]$_DFFE_PN0P_  (.D(_0005_),
    .Q(net112),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[15]$_DFFE_PN0P_  (.D(_0006_),
    .Q(net113),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[16]$_DFFE_PN0P_  (.D(_0007_),
    .Q(net114),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[17]$_DFFE_PN0P_  (.D(_0008_),
    .Q(net115),
    .RESET_B(net105),
    .CLK(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[18]$_DFFE_PN0P_  (.D(_0009_),
    .Q(net116),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[19]$_DFFE_PN0P_  (.D(_0010_),
    .Q(net117),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[1]$_DFFE_PN0P_  (.D(_0011_),
    .Q(net118),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[20]$_DFFE_PN0P_  (.D(_0012_),
    .Q(net119),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[21]$_DFFE_PN0P_  (.D(_0013_),
    .Q(net120),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[22]$_DFFE_PN0P_  (.D(_0014_),
    .Q(net121),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[23]$_DFFE_PN0P_  (.D(_0015_),
    .Q(net122),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \addr_last_q[24]$_DFFE_PN0P_  (.D(_0016_),
    .Q(net123),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[25]$_DFFE_PN0P_  (.D(_0017_),
    .Q(net124),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[26]$_DFFE_PN0P_  (.D(_0018_),
    .Q(net125),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[27]$_DFFE_PN0P_  (.D(_0019_),
    .Q(net126),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[28]$_DFFE_PN0P_  (.D(_0020_),
    .Q(net127),
    .RESET_B(net105),
    .CLK(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[29]$_DFFE_PN0P_  (.D(_0021_),
    .Q(net128),
    .RESET_B(net105),
    .CLK(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[2]$_DFFE_PN0P_  (.D(_0022_),
    .Q(net129),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[30]$_DFFE_PN0P_  (.D(_0023_),
    .Q(net130),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \addr_last_q[31]$_DFFE_PN0P_  (.D(_0024_),
    .Q(net131),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[3]$_DFFE_PN0P_  (.D(_0025_),
    .Q(net132),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[4]$_DFFE_PN0P_  (.D(_0026_),
    .Q(net133),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[5]$_DFFE_PN0P_  (.D(_0027_),
    .Q(net134),
    .RESET_B(net105),
    .CLK(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[6]$_DFFE_PN0P_  (.D(_0028_),
    .Q(net135),
    .RESET_B(net105),
    .CLK(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[7]$_DFFE_PN0P_  (.D(_0029_),
    .Q(net136),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[8]$_DFFE_PN0P_  (.D(_0030_),
    .Q(net137),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \addr_last_q[9]$_DFFE_PN0P_  (.D(_0031_),
    .Q(net138),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \data_sign_ext_q$_DFFE_PN0P_  (.D(_0032_),
    .Q(data_sign_ext_q),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \data_type_q[0]$_DFFE_PN0P_  (.D(_0033_),
    .Q(\data_type_q[0] ),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \data_type_q[1]$_DFFE_PN0P_  (.D(_0034_),
    .Q(\data_type_q[1] ),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \data_we_q$_DFFE_PN0P_  (.D(_0035_),
    .Q(data_we_q),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \handle_misaligned_q$_DFFE_PN0P_  (.D(_0036_),
    .Q(handle_misaligned_q),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \ls_fsm_cs[0]$_DFF_PN0_  (.D(\ls_fsm_ns[0] ),
    .Q(\ls_fsm_cs[0] ),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \ls_fsm_cs[1]$_DFF_PN0_  (.D(\ls_fsm_ns[1] ),
    .Q(\ls_fsm_cs[1] ),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \ls_fsm_cs[2]$_DFF_PN0_  (.D(\ls_fsm_ns[2] ),
    .Q(\ls_fsm_cs[2] ),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \lsu_err_q$_DFFE_PN0P_  (.D(_0037_),
    .Q(lsu_err_q),
    .RESET_B(net105),
    .CLK(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \pmp_err_q$_DFFE_PN0P_  (.D(_0038_),
    .Q(pmp_err_q),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_offset_q[0]$_DFFE_PN0P_  (.D(_0039_),
    .Q(\rdata_offset_q[0] ),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_offset_q[1]$_DFFE_PN0P_  (.D(_0040_),
    .Q(\rdata_offset_q[1] ),
    .RESET_B(net105),
    .CLK(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[0]$_DFFE_PN0P_  (.D(_0041_),
    .Q(\rdata_q[8] ),
    .RESET_B(net105),
    .CLK(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[10]$_DFFE_PN0P_  (.D(_0042_),
    .Q(\rdata_q[18] ),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[11]$_DFFE_PN0P_  (.D(_0043_),
    .Q(\rdata_q[19] ),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[12]$_DFFE_PN0P_  (.D(_0044_),
    .Q(\rdata_q[20] ),
    .RESET_B(net105),
    .CLK(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[13]$_DFFE_PN0P_  (.D(_0045_),
    .Q(\rdata_q[21] ),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[14]$_DFFE_PN0P_  (.D(_0046_),
    .Q(\rdata_q[22] ),
    .RESET_B(net105),
    .CLK(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[15]$_DFFE_PN0P_  (.D(_0047_),
    .Q(\rdata_q[23] ),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[16]$_DFFE_PN0P_  (.D(_0048_),
    .Q(\rdata_q[24] ),
    .RESET_B(net105),
    .CLK(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[17]$_DFFE_PN0P_  (.D(_0049_),
    .Q(\rdata_q[25] ),
    .RESET_B(net105),
    .CLK(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[18]$_DFFE_PN0P_  (.D(_0050_),
    .Q(\rdata_q[26] ),
    .RESET_B(net105),
    .CLK(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[19]$_DFFE_PN0P_  (.D(_0051_),
    .Q(\rdata_q[27] ),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[1]$_DFFE_PN0P_  (.D(_0052_),
    .Q(\rdata_q[9] ),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[20]$_DFFE_PN0P_  (.D(_0053_),
    .Q(\rdata_q[28] ),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[21]$_DFFE_PN0P_  (.D(_0054_),
    .Q(\rdata_q[29] ),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[22]$_DFFE_PN0P_  (.D(_0055_),
    .Q(\rdata_q[30] ),
    .RESET_B(net105),
    .CLK(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[23]$_DFFE_PN0P_  (.D(_0056_),
    .Q(\rdata_q[31] ),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[2]$_DFFE_PN0P_  (.D(_0057_),
    .Q(\rdata_q[10] ),
    .RESET_B(net105),
    .CLK(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[3]$_DFFE_PN0P_  (.D(_0058_),
    .Q(\rdata_q[11] ),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[4]$_DFFE_PN0P_  (.D(_0059_),
    .Q(\rdata_q[12] ),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[5]$_DFFE_PN0P_  (.D(_0060_),
    .Q(\rdata_q[13] ),
    .RESET_B(net105),
    .CLK(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[6]$_DFFE_PN0P_  (.D(_0061_),
    .Q(\rdata_q[14] ),
    .RESET_B(net105),
    .CLK(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[7]$_DFFE_PN0P_  (.D(_0062_),
    .Q(\rdata_q[15] ),
    .RESET_B(net105),
    .CLK(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[8]$_DFFE_PN0P_  (.D(_0063_),
    .Q(\rdata_q[16] ),
    .RESET_B(net105),
    .CLK(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rdata_q[9]$_DFFE_PN0P_  (.D(_0064_),
    .Q(\rdata_q[17] ),
    .RESET_B(net105),
    .CLK(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_279 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(adder_result_ex_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(adder_result_ex_i[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(adder_result_ex_i[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(adder_result_ex_i[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(adder_result_ex_i[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(adder_result_ex_i[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(adder_result_ex_i[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(adder_result_ex_i[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(adder_result_ex_i[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(adder_result_ex_i[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(adder_result_ex_i[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(adder_result_ex_i[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(adder_result_ex_i[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(adder_result_ex_i[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(adder_result_ex_i[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(adder_result_ex_i[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(adder_result_ex_i[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(adder_result_ex_i[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(adder_result_ex_i[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(adder_result_ex_i[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(adder_result_ex_i[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(adder_result_ex_i[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(adder_result_ex_i[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(adder_result_ex_i[30]),
    .X(net24));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input25 (.A(adder_result_ex_i[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(adder_result_ex_i[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(adder_result_ex_i[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(adder_result_ex_i[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(adder_result_ex_i[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(adder_result_ex_i[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(adder_result_ex_i[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(adder_result_ex_i[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(data_err_i),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(data_gnt_i),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(data_pmp_err_i),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(data_rdata_i[0]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(data_rdata_i[10]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(data_rdata_i[11]),
    .X(net38));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input39 (.A(data_rdata_i[12]),
    .X(net39));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input40 (.A(data_rdata_i[13]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(data_rdata_i[14]),
    .X(net41));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input42 (.A(data_rdata_i[15]),
    .X(net42));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input43 (.A(data_rdata_i[16]),
    .X(net43));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input44 (.A(data_rdata_i[17]),
    .X(net44));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input45 (.A(data_rdata_i[18]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(data_rdata_i[19]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(data_rdata_i[1]),
    .X(net47));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input48 (.A(data_rdata_i[20]),
    .X(net48));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input49 (.A(data_rdata_i[21]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(data_rdata_i[22]),
    .X(net50));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input51 (.A(data_rdata_i[23]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(data_rdata_i[24]),
    .X(net52));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input53 (.A(data_rdata_i[25]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(data_rdata_i[26]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(data_rdata_i[27]),
    .X(net55));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input56 (.A(data_rdata_i[28]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(data_rdata_i[29]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(data_rdata_i[2]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(data_rdata_i[30]),
    .X(net59));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input60 (.A(data_rdata_i[31]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(data_rdata_i[3]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(data_rdata_i[4]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(data_rdata_i[5]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(data_rdata_i[6]),
    .X(net64));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input65 (.A(data_rdata_i[7]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(data_rdata_i[8]),
    .X(net66));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input67 (.A(data_rdata_i[9]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(data_rvalid_i),
    .X(net68));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input69 (.A(lsu_req_i),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(lsu_sign_ext_i),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(lsu_type_i[1]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(lsu_wdata_i[0]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(lsu_wdata_i[10]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(lsu_wdata_i[11]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(lsu_wdata_i[12]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(lsu_wdata_i[13]),
    .X(net76));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input77 (.A(lsu_wdata_i[14]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(lsu_wdata_i[15]),
    .X(net78));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input79 (.A(lsu_wdata_i[16]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(lsu_wdata_i[17]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(lsu_wdata_i[18]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(lsu_wdata_i[19]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(lsu_wdata_i[1]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(lsu_wdata_i[20]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(lsu_wdata_i[21]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(lsu_wdata_i[22]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(lsu_wdata_i[23]),
    .X(net87));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input88 (.A(lsu_wdata_i[24]),
    .X(net88));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input89 (.A(lsu_wdata_i[25]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(lsu_wdata_i[26]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(lsu_wdata_i[27]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(lsu_wdata_i[28]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(lsu_wdata_i[29]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(lsu_wdata_i[2]),
    .X(net94));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input95 (.A(lsu_wdata_i[30]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 input96 (.A(lsu_wdata_i[31]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(lsu_wdata_i[3]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(lsu_wdata_i[4]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(lsu_wdata_i[5]),
    .X(net99));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input100 (.A(lsu_wdata_i[6]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(lsu_wdata_i[7]),
    .X(net101));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input102 (.A(lsu_wdata_i[8]),
    .X(net102));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input103 (.A(lsu_wdata_i[9]),
    .X(net103));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input104 (.A(lsu_we_i),
    .X(net104));
 sky130_fd_sc_hd__buf_16 input105 (.A(rst_ni),
    .X(net105));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(addr_incr_req_o));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(addr_last_o[0]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(addr_last_o[10]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(addr_last_o[11]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(addr_last_o[12]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(addr_last_o[13]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(addr_last_o[14]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(addr_last_o[15]));
 sky130_fd_sc_hd__buf_1 output114 (.A(net114),
    .X(addr_last_o[16]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(addr_last_o[17]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(addr_last_o[18]));
 sky130_fd_sc_hd__buf_1 output117 (.A(net117),
    .X(addr_last_o[19]));
 sky130_fd_sc_hd__buf_1 output118 (.A(net118),
    .X(addr_last_o[1]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(addr_last_o[20]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(addr_last_o[21]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(addr_last_o[22]));
 sky130_fd_sc_hd__buf_1 output122 (.A(net122),
    .X(addr_last_o[23]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(addr_last_o[24]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(addr_last_o[25]));
 sky130_fd_sc_hd__buf_1 output125 (.A(net125),
    .X(addr_last_o[26]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(addr_last_o[27]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(addr_last_o[28]));
 sky130_fd_sc_hd__buf_1 output128 (.A(net128),
    .X(addr_last_o[29]));
 sky130_fd_sc_hd__buf_1 output129 (.A(net129),
    .X(addr_last_o[2]));
 sky130_fd_sc_hd__buf_1 output130 (.A(net130),
    .X(addr_last_o[30]));
 sky130_fd_sc_hd__buf_1 output131 (.A(net131),
    .X(addr_last_o[31]));
 sky130_fd_sc_hd__buf_1 output132 (.A(net132),
    .X(addr_last_o[3]));
 sky130_fd_sc_hd__buf_1 output133 (.A(net133),
    .X(addr_last_o[4]));
 sky130_fd_sc_hd__buf_1 output134 (.A(net134),
    .X(addr_last_o[5]));
 sky130_fd_sc_hd__buf_1 output135 (.A(net135),
    .X(addr_last_o[6]));
 sky130_fd_sc_hd__buf_1 output136 (.A(net136),
    .X(addr_last_o[7]));
 sky130_fd_sc_hd__buf_1 output137 (.A(net137),
    .X(addr_last_o[8]));
 sky130_fd_sc_hd__buf_1 output138 (.A(net138),
    .X(addr_last_o[9]));
 sky130_fd_sc_hd__buf_1 output139 (.A(net139),
    .X(busy_o));
 sky130_fd_sc_hd__buf_1 output140 (.A(net140),
    .X(data_addr_o[10]));
 sky130_fd_sc_hd__buf_1 output141 (.A(net141),
    .X(data_addr_o[11]));
 sky130_fd_sc_hd__buf_1 output142 (.A(net142),
    .X(data_addr_o[12]));
 sky130_fd_sc_hd__buf_1 output143 (.A(net143),
    .X(data_addr_o[13]));
 sky130_fd_sc_hd__buf_1 output144 (.A(net144),
    .X(data_addr_o[14]));
 sky130_fd_sc_hd__buf_1 output145 (.A(net145),
    .X(data_addr_o[15]));
 sky130_fd_sc_hd__buf_1 output146 (.A(net146),
    .X(data_addr_o[16]));
 sky130_fd_sc_hd__buf_1 output147 (.A(net147),
    .X(data_addr_o[17]));
 sky130_fd_sc_hd__buf_1 output148 (.A(net148),
    .X(data_addr_o[18]));
 sky130_fd_sc_hd__buf_1 output149 (.A(net149),
    .X(data_addr_o[19]));
 sky130_fd_sc_hd__buf_1 output150 (.A(net150),
    .X(data_addr_o[20]));
 sky130_fd_sc_hd__buf_1 output151 (.A(net151),
    .X(data_addr_o[21]));
 sky130_fd_sc_hd__buf_1 output152 (.A(net152),
    .X(data_addr_o[22]));
 sky130_fd_sc_hd__buf_1 output153 (.A(net153),
    .X(data_addr_o[23]));
 sky130_fd_sc_hd__buf_1 output154 (.A(net154),
    .X(data_addr_o[24]));
 sky130_fd_sc_hd__buf_1 output155 (.A(net155),
    .X(data_addr_o[25]));
 sky130_fd_sc_hd__buf_1 output156 (.A(net156),
    .X(data_addr_o[26]));
 sky130_fd_sc_hd__buf_1 output157 (.A(net157),
    .X(data_addr_o[27]));
 sky130_fd_sc_hd__buf_1 output158 (.A(net158),
    .X(data_addr_o[28]));
 sky130_fd_sc_hd__buf_1 output159 (.A(net159),
    .X(data_addr_o[29]));
 sky130_fd_sc_hd__buf_1 output160 (.A(net160),
    .X(data_addr_o[2]));
 sky130_fd_sc_hd__buf_1 output161 (.A(net161),
    .X(data_addr_o[30]));
 sky130_fd_sc_hd__buf_1 output162 (.A(net162),
    .X(data_addr_o[31]));
 sky130_fd_sc_hd__buf_1 output163 (.A(net163),
    .X(data_addr_o[3]));
 sky130_fd_sc_hd__buf_1 output164 (.A(net164),
    .X(data_addr_o[4]));
 sky130_fd_sc_hd__buf_1 output165 (.A(net165),
    .X(data_addr_o[5]));
 sky130_fd_sc_hd__buf_1 output166 (.A(net166),
    .X(data_addr_o[6]));
 sky130_fd_sc_hd__buf_1 output167 (.A(net167),
    .X(data_addr_o[7]));
 sky130_fd_sc_hd__buf_1 output168 (.A(net168),
    .X(data_addr_o[8]));
 sky130_fd_sc_hd__buf_1 output169 (.A(net169),
    .X(data_addr_o[9]));
 sky130_fd_sc_hd__buf_1 output170 (.A(net170),
    .X(data_be_o[0]));
 sky130_fd_sc_hd__buf_1 output171 (.A(net171),
    .X(data_be_o[1]));
 sky130_fd_sc_hd__buf_1 output172 (.A(net172),
    .X(data_be_o[2]));
 sky130_fd_sc_hd__buf_1 output173 (.A(net173),
    .X(data_be_o[3]));
 sky130_fd_sc_hd__buf_1 output174 (.A(net174),
    .X(data_req_o));
 sky130_fd_sc_hd__buf_1 output175 (.A(net175),
    .X(data_wdata_o[0]));
 sky130_fd_sc_hd__buf_1 output176 (.A(net176),
    .X(data_wdata_o[10]));
 sky130_fd_sc_hd__buf_1 output177 (.A(net177),
    .X(data_wdata_o[11]));
 sky130_fd_sc_hd__buf_1 output178 (.A(net178),
    .X(data_wdata_o[12]));
 sky130_fd_sc_hd__buf_1 output179 (.A(net179),
    .X(data_wdata_o[13]));
 sky130_fd_sc_hd__buf_1 output180 (.A(net180),
    .X(data_wdata_o[14]));
 sky130_fd_sc_hd__buf_1 output181 (.A(net181),
    .X(data_wdata_o[15]));
 sky130_fd_sc_hd__buf_1 output182 (.A(net182),
    .X(data_wdata_o[16]));
 sky130_fd_sc_hd__buf_1 output183 (.A(net183),
    .X(data_wdata_o[17]));
 sky130_fd_sc_hd__buf_1 output184 (.A(net184),
    .X(data_wdata_o[18]));
 sky130_fd_sc_hd__buf_1 output185 (.A(net185),
    .X(data_wdata_o[19]));
 sky130_fd_sc_hd__buf_1 output186 (.A(net186),
    .X(data_wdata_o[1]));
 sky130_fd_sc_hd__buf_1 output187 (.A(net187),
    .X(data_wdata_o[20]));
 sky130_fd_sc_hd__buf_1 output188 (.A(net188),
    .X(data_wdata_o[21]));
 sky130_fd_sc_hd__buf_1 output189 (.A(net189),
    .X(data_wdata_o[22]));
 sky130_fd_sc_hd__buf_1 output190 (.A(net190),
    .X(data_wdata_o[23]));
 sky130_fd_sc_hd__buf_1 output191 (.A(net191),
    .X(data_wdata_o[24]));
 sky130_fd_sc_hd__buf_1 output192 (.A(net192),
    .X(data_wdata_o[25]));
 sky130_fd_sc_hd__buf_1 output193 (.A(net193),
    .X(data_wdata_o[26]));
 sky130_fd_sc_hd__buf_1 output194 (.A(net194),
    .X(data_wdata_o[27]));
 sky130_fd_sc_hd__buf_1 output195 (.A(net195),
    .X(data_wdata_o[28]));
 sky130_fd_sc_hd__buf_1 output196 (.A(net196),
    .X(data_wdata_o[29]));
 sky130_fd_sc_hd__buf_1 output197 (.A(net197),
    .X(data_wdata_o[2]));
 sky130_fd_sc_hd__buf_1 output198 (.A(net198),
    .X(data_wdata_o[30]));
 sky130_fd_sc_hd__buf_1 output199 (.A(net199),
    .X(data_wdata_o[31]));
 sky130_fd_sc_hd__buf_1 output200 (.A(net200),
    .X(data_wdata_o[3]));
 sky130_fd_sc_hd__buf_1 output201 (.A(net201),
    .X(data_wdata_o[4]));
 sky130_fd_sc_hd__buf_1 output202 (.A(net202),
    .X(data_wdata_o[5]));
 sky130_fd_sc_hd__buf_1 output203 (.A(net203),
    .X(data_wdata_o[6]));
 sky130_fd_sc_hd__buf_1 output204 (.A(net204),
    .X(data_wdata_o[7]));
 sky130_fd_sc_hd__buf_1 output205 (.A(net205),
    .X(data_wdata_o[8]));
 sky130_fd_sc_hd__buf_1 output206 (.A(net206),
    .X(data_wdata_o[9]));
 sky130_fd_sc_hd__buf_1 output207 (.A(net207),
    .X(data_we_o));
 sky130_fd_sc_hd__buf_1 output208 (.A(net208),
    .X(load_err_o));
 sky130_fd_sc_hd__buf_1 output209 (.A(net209),
    .X(lsu_rdata_o[0]));
 sky130_fd_sc_hd__buf_1 output210 (.A(net210),
    .X(lsu_rdata_o[10]));
 sky130_fd_sc_hd__buf_1 output211 (.A(net211),
    .X(lsu_rdata_o[11]));
 sky130_fd_sc_hd__buf_1 output212 (.A(net212),
    .X(lsu_rdata_o[12]));
 sky130_fd_sc_hd__buf_1 output213 (.A(net213),
    .X(lsu_rdata_o[13]));
 sky130_fd_sc_hd__buf_1 output214 (.A(net214),
    .X(lsu_rdata_o[14]));
 sky130_fd_sc_hd__buf_1 output215 (.A(net215),
    .X(lsu_rdata_o[15]));
 sky130_fd_sc_hd__buf_1 output216 (.A(net216),
    .X(lsu_rdata_o[16]));
 sky130_fd_sc_hd__buf_1 output217 (.A(net217),
    .X(lsu_rdata_o[17]));
 sky130_fd_sc_hd__buf_1 output218 (.A(net218),
    .X(lsu_rdata_o[18]));
 sky130_fd_sc_hd__buf_1 output219 (.A(net219),
    .X(lsu_rdata_o[19]));
 sky130_fd_sc_hd__buf_1 output220 (.A(net220),
    .X(lsu_rdata_o[1]));
 sky130_fd_sc_hd__buf_1 output221 (.A(net221),
    .X(lsu_rdata_o[20]));
 sky130_fd_sc_hd__buf_1 output222 (.A(net222),
    .X(lsu_rdata_o[21]));
 sky130_fd_sc_hd__buf_1 output223 (.A(net223),
    .X(lsu_rdata_o[22]));
 sky130_fd_sc_hd__buf_1 output224 (.A(net224),
    .X(lsu_rdata_o[23]));
 sky130_fd_sc_hd__buf_1 output225 (.A(net225),
    .X(lsu_rdata_o[24]));
 sky130_fd_sc_hd__buf_1 output226 (.A(net226),
    .X(lsu_rdata_o[25]));
 sky130_fd_sc_hd__buf_1 output227 (.A(net227),
    .X(lsu_rdata_o[26]));
 sky130_fd_sc_hd__buf_1 output228 (.A(net228),
    .X(lsu_rdata_o[27]));
 sky130_fd_sc_hd__buf_1 output229 (.A(net229),
    .X(lsu_rdata_o[28]));
 sky130_fd_sc_hd__buf_1 output230 (.A(net230),
    .X(lsu_rdata_o[29]));
 sky130_fd_sc_hd__buf_1 output231 (.A(net231),
    .X(lsu_rdata_o[2]));
 sky130_fd_sc_hd__buf_1 output232 (.A(net232),
    .X(lsu_rdata_o[30]));
 sky130_fd_sc_hd__buf_1 output233 (.A(net233),
    .X(lsu_rdata_o[31]));
 sky130_fd_sc_hd__buf_1 output234 (.A(net234),
    .X(lsu_rdata_o[3]));
 sky130_fd_sc_hd__buf_1 output235 (.A(net235),
    .X(lsu_rdata_o[4]));
 sky130_fd_sc_hd__buf_1 output236 (.A(net236),
    .X(lsu_rdata_o[5]));
 sky130_fd_sc_hd__buf_1 output237 (.A(net237),
    .X(lsu_rdata_o[6]));
 sky130_fd_sc_hd__buf_1 output238 (.A(net238),
    .X(lsu_rdata_o[7]));
 sky130_fd_sc_hd__buf_1 output239 (.A(net239),
    .X(lsu_rdata_o[8]));
 sky130_fd_sc_hd__buf_1 output240 (.A(net240),
    .X(lsu_rdata_o[9]));
 sky130_fd_sc_hd__buf_1 output241 (.A(net241),
    .X(lsu_rdata_valid_o));
 sky130_fd_sc_hd__buf_1 output242 (.A(net242),
    .X(lsu_req_done_o));
 sky130_fd_sc_hd__buf_1 output243 (.A(net243),
    .X(lsu_resp_valid_o));
 sky130_fd_sc_hd__buf_1 output244 (.A(net244),
    .X(perf_load_o));
 sky130_fd_sc_hd__buf_1 output245 (.A(net245),
    .X(perf_store_o));
 sky130_fd_sc_hd__buf_1 output246 (.A(net246),
    .X(store_err_o));
 sky130_fd_sc_hd__conb_1 _0973__247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 _0974__248 (.LO(net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload3 (.A(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__clkinvlp_4 clkload5 (.A(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload6 (.A(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(lsu_type_i[0]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_5 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_323 ();
endmodule
