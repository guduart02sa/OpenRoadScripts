module ibex_register_file_ff (clk_i,
    dummy_instr_id_i,
    rst_ni,
    test_en_i,
    we_a_i,
    raddr_a_i,
    raddr_b_i,
    rdata_a_o,
    rdata_b_o,
    waddr_a_i,
    wdata_a_i);
 input clk_i;
 input dummy_instr_id_i;
 input rst_ni;
 input test_en_i;
 input we_a_i;
 input [4:0] raddr_a_i;
 input [4:0] raddr_b_i;
 output [31:0] rdata_a_o;
 output [31:0] rdata_b_o;
 input [4:0] waddr_a_i;
 input [31:0] wdata_a_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire \rf_reg[1000] ;
 wire \rf_reg[1001] ;
 wire \rf_reg[1002] ;
 wire \rf_reg[1003] ;
 wire \rf_reg[1004] ;
 wire \rf_reg[1005] ;
 wire \rf_reg[1006] ;
 wire \rf_reg[1007] ;
 wire \rf_reg[1008] ;
 wire \rf_reg[1009] ;
 wire \rf_reg[100] ;
 wire \rf_reg[1010] ;
 wire \rf_reg[1011] ;
 wire \rf_reg[1012] ;
 wire \rf_reg[1013] ;
 wire \rf_reg[1014] ;
 wire \rf_reg[1015] ;
 wire \rf_reg[1016] ;
 wire \rf_reg[1017] ;
 wire \rf_reg[1018] ;
 wire \rf_reg[1019] ;
 wire \rf_reg[101] ;
 wire \rf_reg[1020] ;
 wire \rf_reg[1021] ;
 wire \rf_reg[1022] ;
 wire \rf_reg[1023] ;
 wire \rf_reg[102] ;
 wire \rf_reg[103] ;
 wire \rf_reg[104] ;
 wire \rf_reg[105] ;
 wire \rf_reg[106] ;
 wire \rf_reg[107] ;
 wire \rf_reg[108] ;
 wire \rf_reg[109] ;
 wire \rf_reg[110] ;
 wire \rf_reg[111] ;
 wire \rf_reg[112] ;
 wire \rf_reg[113] ;
 wire \rf_reg[114] ;
 wire \rf_reg[115] ;
 wire \rf_reg[116] ;
 wire \rf_reg[117] ;
 wire \rf_reg[118] ;
 wire \rf_reg[119] ;
 wire \rf_reg[120] ;
 wire \rf_reg[121] ;
 wire \rf_reg[122] ;
 wire \rf_reg[123] ;
 wire \rf_reg[124] ;
 wire \rf_reg[125] ;
 wire \rf_reg[126] ;
 wire \rf_reg[127] ;
 wire \rf_reg[128] ;
 wire \rf_reg[129] ;
 wire \rf_reg[130] ;
 wire \rf_reg[131] ;
 wire \rf_reg[132] ;
 wire \rf_reg[133] ;
 wire \rf_reg[134] ;
 wire \rf_reg[135] ;
 wire \rf_reg[136] ;
 wire \rf_reg[137] ;
 wire \rf_reg[138] ;
 wire \rf_reg[139] ;
 wire \rf_reg[140] ;
 wire \rf_reg[141] ;
 wire \rf_reg[142] ;
 wire \rf_reg[143] ;
 wire \rf_reg[144] ;
 wire \rf_reg[145] ;
 wire \rf_reg[146] ;
 wire \rf_reg[147] ;
 wire \rf_reg[148] ;
 wire \rf_reg[149] ;
 wire \rf_reg[150] ;
 wire \rf_reg[151] ;
 wire \rf_reg[152] ;
 wire \rf_reg[153] ;
 wire \rf_reg[154] ;
 wire \rf_reg[155] ;
 wire \rf_reg[156] ;
 wire \rf_reg[157] ;
 wire \rf_reg[158] ;
 wire \rf_reg[159] ;
 wire \rf_reg[160] ;
 wire \rf_reg[161] ;
 wire \rf_reg[162] ;
 wire \rf_reg[163] ;
 wire \rf_reg[164] ;
 wire \rf_reg[165] ;
 wire \rf_reg[166] ;
 wire \rf_reg[167] ;
 wire \rf_reg[168] ;
 wire \rf_reg[169] ;
 wire \rf_reg[170] ;
 wire \rf_reg[171] ;
 wire \rf_reg[172] ;
 wire \rf_reg[173] ;
 wire \rf_reg[174] ;
 wire \rf_reg[175] ;
 wire \rf_reg[176] ;
 wire \rf_reg[177] ;
 wire \rf_reg[178] ;
 wire \rf_reg[179] ;
 wire \rf_reg[180] ;
 wire \rf_reg[181] ;
 wire \rf_reg[182] ;
 wire \rf_reg[183] ;
 wire \rf_reg[184] ;
 wire \rf_reg[185] ;
 wire \rf_reg[186] ;
 wire \rf_reg[187] ;
 wire \rf_reg[188] ;
 wire \rf_reg[189] ;
 wire \rf_reg[190] ;
 wire \rf_reg[191] ;
 wire \rf_reg[192] ;
 wire \rf_reg[193] ;
 wire \rf_reg[194] ;
 wire \rf_reg[195] ;
 wire \rf_reg[196] ;
 wire \rf_reg[197] ;
 wire \rf_reg[198] ;
 wire \rf_reg[199] ;
 wire \rf_reg[200] ;
 wire \rf_reg[201] ;
 wire \rf_reg[202] ;
 wire \rf_reg[203] ;
 wire \rf_reg[204] ;
 wire \rf_reg[205] ;
 wire \rf_reg[206] ;
 wire \rf_reg[207] ;
 wire \rf_reg[208] ;
 wire \rf_reg[209] ;
 wire \rf_reg[210] ;
 wire \rf_reg[211] ;
 wire \rf_reg[212] ;
 wire \rf_reg[213] ;
 wire \rf_reg[214] ;
 wire \rf_reg[215] ;
 wire \rf_reg[216] ;
 wire \rf_reg[217] ;
 wire \rf_reg[218] ;
 wire \rf_reg[219] ;
 wire \rf_reg[220] ;
 wire \rf_reg[221] ;
 wire \rf_reg[222] ;
 wire \rf_reg[223] ;
 wire \rf_reg[224] ;
 wire \rf_reg[225] ;
 wire \rf_reg[226] ;
 wire \rf_reg[227] ;
 wire \rf_reg[228] ;
 wire \rf_reg[229] ;
 wire \rf_reg[230] ;
 wire \rf_reg[231] ;
 wire \rf_reg[232] ;
 wire \rf_reg[233] ;
 wire \rf_reg[234] ;
 wire \rf_reg[235] ;
 wire \rf_reg[236] ;
 wire \rf_reg[237] ;
 wire \rf_reg[238] ;
 wire \rf_reg[239] ;
 wire \rf_reg[240] ;
 wire \rf_reg[241] ;
 wire \rf_reg[242] ;
 wire \rf_reg[243] ;
 wire \rf_reg[244] ;
 wire \rf_reg[245] ;
 wire \rf_reg[246] ;
 wire \rf_reg[247] ;
 wire \rf_reg[248] ;
 wire \rf_reg[249] ;
 wire \rf_reg[250] ;
 wire \rf_reg[251] ;
 wire \rf_reg[252] ;
 wire \rf_reg[253] ;
 wire \rf_reg[254] ;
 wire \rf_reg[255] ;
 wire \rf_reg[256] ;
 wire \rf_reg[257] ;
 wire \rf_reg[258] ;
 wire \rf_reg[259] ;
 wire \rf_reg[260] ;
 wire \rf_reg[261] ;
 wire \rf_reg[262] ;
 wire \rf_reg[263] ;
 wire \rf_reg[264] ;
 wire \rf_reg[265] ;
 wire \rf_reg[266] ;
 wire \rf_reg[267] ;
 wire \rf_reg[268] ;
 wire \rf_reg[269] ;
 wire \rf_reg[270] ;
 wire \rf_reg[271] ;
 wire \rf_reg[272] ;
 wire \rf_reg[273] ;
 wire \rf_reg[274] ;
 wire \rf_reg[275] ;
 wire \rf_reg[276] ;
 wire \rf_reg[277] ;
 wire \rf_reg[278] ;
 wire \rf_reg[279] ;
 wire \rf_reg[280] ;
 wire \rf_reg[281] ;
 wire \rf_reg[282] ;
 wire \rf_reg[283] ;
 wire \rf_reg[284] ;
 wire \rf_reg[285] ;
 wire \rf_reg[286] ;
 wire \rf_reg[287] ;
 wire \rf_reg[288] ;
 wire \rf_reg[289] ;
 wire \rf_reg[290] ;
 wire \rf_reg[291] ;
 wire \rf_reg[292] ;
 wire \rf_reg[293] ;
 wire \rf_reg[294] ;
 wire \rf_reg[295] ;
 wire \rf_reg[296] ;
 wire \rf_reg[297] ;
 wire \rf_reg[298] ;
 wire \rf_reg[299] ;
 wire \rf_reg[300] ;
 wire \rf_reg[301] ;
 wire \rf_reg[302] ;
 wire \rf_reg[303] ;
 wire \rf_reg[304] ;
 wire \rf_reg[305] ;
 wire \rf_reg[306] ;
 wire \rf_reg[307] ;
 wire \rf_reg[308] ;
 wire \rf_reg[309] ;
 wire \rf_reg[310] ;
 wire \rf_reg[311] ;
 wire \rf_reg[312] ;
 wire \rf_reg[313] ;
 wire \rf_reg[314] ;
 wire \rf_reg[315] ;
 wire \rf_reg[316] ;
 wire \rf_reg[317] ;
 wire \rf_reg[318] ;
 wire \rf_reg[319] ;
 wire \rf_reg[320] ;
 wire \rf_reg[321] ;
 wire \rf_reg[322] ;
 wire \rf_reg[323] ;
 wire \rf_reg[324] ;
 wire \rf_reg[325] ;
 wire \rf_reg[326] ;
 wire \rf_reg[327] ;
 wire \rf_reg[328] ;
 wire \rf_reg[329] ;
 wire \rf_reg[32] ;
 wire \rf_reg[330] ;
 wire \rf_reg[331] ;
 wire \rf_reg[332] ;
 wire \rf_reg[333] ;
 wire \rf_reg[334] ;
 wire \rf_reg[335] ;
 wire \rf_reg[336] ;
 wire \rf_reg[337] ;
 wire \rf_reg[338] ;
 wire \rf_reg[339] ;
 wire \rf_reg[33] ;
 wire \rf_reg[340] ;
 wire \rf_reg[341] ;
 wire \rf_reg[342] ;
 wire \rf_reg[343] ;
 wire \rf_reg[344] ;
 wire \rf_reg[345] ;
 wire \rf_reg[346] ;
 wire \rf_reg[347] ;
 wire \rf_reg[348] ;
 wire \rf_reg[349] ;
 wire \rf_reg[34] ;
 wire \rf_reg[350] ;
 wire \rf_reg[351] ;
 wire \rf_reg[352] ;
 wire \rf_reg[353] ;
 wire \rf_reg[354] ;
 wire \rf_reg[355] ;
 wire \rf_reg[356] ;
 wire \rf_reg[357] ;
 wire \rf_reg[358] ;
 wire \rf_reg[359] ;
 wire \rf_reg[35] ;
 wire \rf_reg[360] ;
 wire \rf_reg[361] ;
 wire \rf_reg[362] ;
 wire \rf_reg[363] ;
 wire \rf_reg[364] ;
 wire \rf_reg[365] ;
 wire \rf_reg[366] ;
 wire \rf_reg[367] ;
 wire \rf_reg[368] ;
 wire \rf_reg[369] ;
 wire \rf_reg[36] ;
 wire \rf_reg[370] ;
 wire \rf_reg[371] ;
 wire \rf_reg[372] ;
 wire \rf_reg[373] ;
 wire \rf_reg[374] ;
 wire \rf_reg[375] ;
 wire \rf_reg[376] ;
 wire \rf_reg[377] ;
 wire \rf_reg[378] ;
 wire \rf_reg[379] ;
 wire \rf_reg[37] ;
 wire \rf_reg[380] ;
 wire \rf_reg[381] ;
 wire \rf_reg[382] ;
 wire \rf_reg[383] ;
 wire \rf_reg[384] ;
 wire \rf_reg[385] ;
 wire \rf_reg[386] ;
 wire \rf_reg[387] ;
 wire \rf_reg[388] ;
 wire \rf_reg[389] ;
 wire \rf_reg[38] ;
 wire \rf_reg[390] ;
 wire \rf_reg[391] ;
 wire \rf_reg[392] ;
 wire \rf_reg[393] ;
 wire \rf_reg[394] ;
 wire \rf_reg[395] ;
 wire \rf_reg[396] ;
 wire \rf_reg[397] ;
 wire \rf_reg[398] ;
 wire \rf_reg[399] ;
 wire \rf_reg[39] ;
 wire \rf_reg[400] ;
 wire \rf_reg[401] ;
 wire \rf_reg[402] ;
 wire \rf_reg[403] ;
 wire \rf_reg[404] ;
 wire \rf_reg[405] ;
 wire \rf_reg[406] ;
 wire \rf_reg[407] ;
 wire \rf_reg[408] ;
 wire \rf_reg[409] ;
 wire \rf_reg[40] ;
 wire \rf_reg[410] ;
 wire \rf_reg[411] ;
 wire \rf_reg[412] ;
 wire \rf_reg[413] ;
 wire \rf_reg[414] ;
 wire \rf_reg[415] ;
 wire \rf_reg[416] ;
 wire \rf_reg[417] ;
 wire \rf_reg[418] ;
 wire \rf_reg[419] ;
 wire \rf_reg[41] ;
 wire \rf_reg[420] ;
 wire \rf_reg[421] ;
 wire \rf_reg[422] ;
 wire \rf_reg[423] ;
 wire \rf_reg[424] ;
 wire \rf_reg[425] ;
 wire \rf_reg[426] ;
 wire \rf_reg[427] ;
 wire \rf_reg[428] ;
 wire \rf_reg[429] ;
 wire \rf_reg[42] ;
 wire \rf_reg[430] ;
 wire \rf_reg[431] ;
 wire \rf_reg[432] ;
 wire \rf_reg[433] ;
 wire \rf_reg[434] ;
 wire \rf_reg[435] ;
 wire \rf_reg[436] ;
 wire \rf_reg[437] ;
 wire \rf_reg[438] ;
 wire \rf_reg[439] ;
 wire \rf_reg[43] ;
 wire \rf_reg[440] ;
 wire \rf_reg[441] ;
 wire \rf_reg[442] ;
 wire \rf_reg[443] ;
 wire \rf_reg[444] ;
 wire \rf_reg[445] ;
 wire \rf_reg[446] ;
 wire \rf_reg[447] ;
 wire \rf_reg[448] ;
 wire \rf_reg[449] ;
 wire \rf_reg[44] ;
 wire \rf_reg[450] ;
 wire \rf_reg[451] ;
 wire \rf_reg[452] ;
 wire \rf_reg[453] ;
 wire \rf_reg[454] ;
 wire \rf_reg[455] ;
 wire \rf_reg[456] ;
 wire \rf_reg[457] ;
 wire \rf_reg[458] ;
 wire \rf_reg[459] ;
 wire \rf_reg[45] ;
 wire \rf_reg[460] ;
 wire \rf_reg[461] ;
 wire \rf_reg[462] ;
 wire \rf_reg[463] ;
 wire \rf_reg[464] ;
 wire \rf_reg[465] ;
 wire \rf_reg[466] ;
 wire \rf_reg[467] ;
 wire \rf_reg[468] ;
 wire \rf_reg[469] ;
 wire \rf_reg[46] ;
 wire \rf_reg[470] ;
 wire \rf_reg[471] ;
 wire \rf_reg[472] ;
 wire \rf_reg[473] ;
 wire \rf_reg[474] ;
 wire \rf_reg[475] ;
 wire \rf_reg[476] ;
 wire \rf_reg[477] ;
 wire \rf_reg[478] ;
 wire \rf_reg[479] ;
 wire \rf_reg[47] ;
 wire \rf_reg[480] ;
 wire \rf_reg[481] ;
 wire \rf_reg[482] ;
 wire \rf_reg[483] ;
 wire \rf_reg[484] ;
 wire \rf_reg[485] ;
 wire \rf_reg[486] ;
 wire \rf_reg[487] ;
 wire \rf_reg[488] ;
 wire \rf_reg[489] ;
 wire \rf_reg[48] ;
 wire \rf_reg[490] ;
 wire \rf_reg[491] ;
 wire \rf_reg[492] ;
 wire \rf_reg[493] ;
 wire \rf_reg[494] ;
 wire \rf_reg[495] ;
 wire \rf_reg[496] ;
 wire \rf_reg[497] ;
 wire \rf_reg[498] ;
 wire \rf_reg[499] ;
 wire \rf_reg[49] ;
 wire \rf_reg[500] ;
 wire \rf_reg[501] ;
 wire \rf_reg[502] ;
 wire \rf_reg[503] ;
 wire \rf_reg[504] ;
 wire \rf_reg[505] ;
 wire \rf_reg[506] ;
 wire \rf_reg[507] ;
 wire \rf_reg[508] ;
 wire \rf_reg[509] ;
 wire \rf_reg[50] ;
 wire \rf_reg[510] ;
 wire \rf_reg[511] ;
 wire \rf_reg[512] ;
 wire \rf_reg[513] ;
 wire \rf_reg[514] ;
 wire \rf_reg[515] ;
 wire \rf_reg[516] ;
 wire \rf_reg[517] ;
 wire \rf_reg[518] ;
 wire \rf_reg[519] ;
 wire \rf_reg[51] ;
 wire \rf_reg[520] ;
 wire \rf_reg[521] ;
 wire \rf_reg[522] ;
 wire \rf_reg[523] ;
 wire \rf_reg[524] ;
 wire \rf_reg[525] ;
 wire \rf_reg[526] ;
 wire \rf_reg[527] ;
 wire \rf_reg[528] ;
 wire \rf_reg[529] ;
 wire \rf_reg[52] ;
 wire \rf_reg[530] ;
 wire \rf_reg[531] ;
 wire \rf_reg[532] ;
 wire \rf_reg[533] ;
 wire \rf_reg[534] ;
 wire \rf_reg[535] ;
 wire \rf_reg[536] ;
 wire \rf_reg[537] ;
 wire \rf_reg[538] ;
 wire \rf_reg[539] ;
 wire \rf_reg[53] ;
 wire \rf_reg[540] ;
 wire \rf_reg[541] ;
 wire \rf_reg[542] ;
 wire \rf_reg[543] ;
 wire \rf_reg[544] ;
 wire \rf_reg[545] ;
 wire \rf_reg[546] ;
 wire \rf_reg[547] ;
 wire \rf_reg[548] ;
 wire \rf_reg[549] ;
 wire \rf_reg[54] ;
 wire \rf_reg[550] ;
 wire \rf_reg[551] ;
 wire \rf_reg[552] ;
 wire \rf_reg[553] ;
 wire \rf_reg[554] ;
 wire \rf_reg[555] ;
 wire \rf_reg[556] ;
 wire \rf_reg[557] ;
 wire \rf_reg[558] ;
 wire \rf_reg[559] ;
 wire \rf_reg[55] ;
 wire \rf_reg[560] ;
 wire \rf_reg[561] ;
 wire \rf_reg[562] ;
 wire \rf_reg[563] ;
 wire \rf_reg[564] ;
 wire \rf_reg[565] ;
 wire \rf_reg[566] ;
 wire \rf_reg[567] ;
 wire \rf_reg[568] ;
 wire \rf_reg[569] ;
 wire \rf_reg[56] ;
 wire \rf_reg[570] ;
 wire \rf_reg[571] ;
 wire \rf_reg[572] ;
 wire \rf_reg[573] ;
 wire \rf_reg[574] ;
 wire \rf_reg[575] ;
 wire \rf_reg[576] ;
 wire \rf_reg[577] ;
 wire \rf_reg[578] ;
 wire \rf_reg[579] ;
 wire \rf_reg[57] ;
 wire \rf_reg[580] ;
 wire \rf_reg[581] ;
 wire \rf_reg[582] ;
 wire \rf_reg[583] ;
 wire \rf_reg[584] ;
 wire \rf_reg[585] ;
 wire \rf_reg[586] ;
 wire \rf_reg[587] ;
 wire \rf_reg[588] ;
 wire \rf_reg[589] ;
 wire \rf_reg[58] ;
 wire \rf_reg[590] ;
 wire \rf_reg[591] ;
 wire \rf_reg[592] ;
 wire \rf_reg[593] ;
 wire \rf_reg[594] ;
 wire \rf_reg[595] ;
 wire \rf_reg[596] ;
 wire \rf_reg[597] ;
 wire \rf_reg[598] ;
 wire \rf_reg[599] ;
 wire \rf_reg[59] ;
 wire \rf_reg[600] ;
 wire \rf_reg[601] ;
 wire \rf_reg[602] ;
 wire \rf_reg[603] ;
 wire \rf_reg[604] ;
 wire \rf_reg[605] ;
 wire \rf_reg[606] ;
 wire \rf_reg[607] ;
 wire \rf_reg[608] ;
 wire \rf_reg[609] ;
 wire \rf_reg[60] ;
 wire \rf_reg[610] ;
 wire \rf_reg[611] ;
 wire \rf_reg[612] ;
 wire \rf_reg[613] ;
 wire \rf_reg[614] ;
 wire \rf_reg[615] ;
 wire \rf_reg[616] ;
 wire \rf_reg[617] ;
 wire \rf_reg[618] ;
 wire \rf_reg[619] ;
 wire \rf_reg[61] ;
 wire \rf_reg[620] ;
 wire \rf_reg[621] ;
 wire \rf_reg[622] ;
 wire \rf_reg[623] ;
 wire \rf_reg[624] ;
 wire \rf_reg[625] ;
 wire \rf_reg[626] ;
 wire \rf_reg[627] ;
 wire \rf_reg[628] ;
 wire \rf_reg[629] ;
 wire \rf_reg[62] ;
 wire \rf_reg[630] ;
 wire \rf_reg[631] ;
 wire \rf_reg[632] ;
 wire \rf_reg[633] ;
 wire \rf_reg[634] ;
 wire \rf_reg[635] ;
 wire \rf_reg[636] ;
 wire \rf_reg[637] ;
 wire \rf_reg[638] ;
 wire \rf_reg[639] ;
 wire \rf_reg[63] ;
 wire \rf_reg[640] ;
 wire \rf_reg[641] ;
 wire \rf_reg[642] ;
 wire \rf_reg[643] ;
 wire \rf_reg[644] ;
 wire \rf_reg[645] ;
 wire \rf_reg[646] ;
 wire \rf_reg[647] ;
 wire \rf_reg[648] ;
 wire \rf_reg[649] ;
 wire \rf_reg[64] ;
 wire \rf_reg[650] ;
 wire \rf_reg[651] ;
 wire \rf_reg[652] ;
 wire \rf_reg[653] ;
 wire \rf_reg[654] ;
 wire \rf_reg[655] ;
 wire \rf_reg[656] ;
 wire \rf_reg[657] ;
 wire \rf_reg[658] ;
 wire \rf_reg[659] ;
 wire \rf_reg[65] ;
 wire \rf_reg[660] ;
 wire \rf_reg[661] ;
 wire \rf_reg[662] ;
 wire \rf_reg[663] ;
 wire \rf_reg[664] ;
 wire \rf_reg[665] ;
 wire \rf_reg[666] ;
 wire \rf_reg[667] ;
 wire \rf_reg[668] ;
 wire \rf_reg[669] ;
 wire \rf_reg[66] ;
 wire \rf_reg[670] ;
 wire \rf_reg[671] ;
 wire \rf_reg[672] ;
 wire \rf_reg[673] ;
 wire \rf_reg[674] ;
 wire \rf_reg[675] ;
 wire \rf_reg[676] ;
 wire \rf_reg[677] ;
 wire \rf_reg[678] ;
 wire \rf_reg[679] ;
 wire \rf_reg[67] ;
 wire \rf_reg[680] ;
 wire \rf_reg[681] ;
 wire \rf_reg[682] ;
 wire \rf_reg[683] ;
 wire \rf_reg[684] ;
 wire \rf_reg[685] ;
 wire \rf_reg[686] ;
 wire \rf_reg[687] ;
 wire \rf_reg[688] ;
 wire \rf_reg[689] ;
 wire \rf_reg[68] ;
 wire \rf_reg[690] ;
 wire \rf_reg[691] ;
 wire \rf_reg[692] ;
 wire \rf_reg[693] ;
 wire \rf_reg[694] ;
 wire \rf_reg[695] ;
 wire \rf_reg[696] ;
 wire \rf_reg[697] ;
 wire \rf_reg[698] ;
 wire \rf_reg[699] ;
 wire \rf_reg[69] ;
 wire \rf_reg[700] ;
 wire \rf_reg[701] ;
 wire \rf_reg[702] ;
 wire \rf_reg[703] ;
 wire \rf_reg[704] ;
 wire \rf_reg[705] ;
 wire \rf_reg[706] ;
 wire \rf_reg[707] ;
 wire \rf_reg[708] ;
 wire \rf_reg[709] ;
 wire \rf_reg[70] ;
 wire \rf_reg[710] ;
 wire \rf_reg[711] ;
 wire \rf_reg[712] ;
 wire \rf_reg[713] ;
 wire \rf_reg[714] ;
 wire \rf_reg[715] ;
 wire \rf_reg[716] ;
 wire \rf_reg[717] ;
 wire \rf_reg[718] ;
 wire \rf_reg[719] ;
 wire \rf_reg[71] ;
 wire \rf_reg[720] ;
 wire \rf_reg[721] ;
 wire \rf_reg[722] ;
 wire \rf_reg[723] ;
 wire \rf_reg[724] ;
 wire \rf_reg[725] ;
 wire \rf_reg[726] ;
 wire \rf_reg[727] ;
 wire \rf_reg[728] ;
 wire \rf_reg[729] ;
 wire \rf_reg[72] ;
 wire \rf_reg[730] ;
 wire \rf_reg[731] ;
 wire \rf_reg[732] ;
 wire \rf_reg[733] ;
 wire \rf_reg[734] ;
 wire \rf_reg[735] ;
 wire \rf_reg[736] ;
 wire \rf_reg[737] ;
 wire \rf_reg[738] ;
 wire \rf_reg[739] ;
 wire \rf_reg[73] ;
 wire \rf_reg[740] ;
 wire \rf_reg[741] ;
 wire \rf_reg[742] ;
 wire \rf_reg[743] ;
 wire \rf_reg[744] ;
 wire \rf_reg[745] ;
 wire \rf_reg[746] ;
 wire \rf_reg[747] ;
 wire \rf_reg[748] ;
 wire \rf_reg[749] ;
 wire \rf_reg[74] ;
 wire \rf_reg[750] ;
 wire \rf_reg[751] ;
 wire \rf_reg[752] ;
 wire \rf_reg[753] ;
 wire \rf_reg[754] ;
 wire \rf_reg[755] ;
 wire \rf_reg[756] ;
 wire \rf_reg[757] ;
 wire \rf_reg[758] ;
 wire \rf_reg[759] ;
 wire \rf_reg[75] ;
 wire \rf_reg[760] ;
 wire \rf_reg[761] ;
 wire \rf_reg[762] ;
 wire \rf_reg[763] ;
 wire \rf_reg[764] ;
 wire \rf_reg[765] ;
 wire \rf_reg[766] ;
 wire \rf_reg[767] ;
 wire \rf_reg[768] ;
 wire \rf_reg[769] ;
 wire \rf_reg[76] ;
 wire \rf_reg[770] ;
 wire \rf_reg[771] ;
 wire \rf_reg[772] ;
 wire \rf_reg[773] ;
 wire \rf_reg[774] ;
 wire \rf_reg[775] ;
 wire \rf_reg[776] ;
 wire \rf_reg[777] ;
 wire \rf_reg[778] ;
 wire \rf_reg[779] ;
 wire \rf_reg[77] ;
 wire \rf_reg[780] ;
 wire \rf_reg[781] ;
 wire \rf_reg[782] ;
 wire \rf_reg[783] ;
 wire \rf_reg[784] ;
 wire \rf_reg[785] ;
 wire \rf_reg[786] ;
 wire \rf_reg[787] ;
 wire \rf_reg[788] ;
 wire \rf_reg[789] ;
 wire \rf_reg[78] ;
 wire \rf_reg[790] ;
 wire \rf_reg[791] ;
 wire \rf_reg[792] ;
 wire \rf_reg[793] ;
 wire \rf_reg[794] ;
 wire \rf_reg[795] ;
 wire \rf_reg[796] ;
 wire \rf_reg[797] ;
 wire \rf_reg[798] ;
 wire \rf_reg[799] ;
 wire \rf_reg[79] ;
 wire \rf_reg[800] ;
 wire \rf_reg[801] ;
 wire \rf_reg[802] ;
 wire \rf_reg[803] ;
 wire \rf_reg[804] ;
 wire \rf_reg[805] ;
 wire \rf_reg[806] ;
 wire \rf_reg[807] ;
 wire \rf_reg[808] ;
 wire \rf_reg[809] ;
 wire \rf_reg[80] ;
 wire \rf_reg[810] ;
 wire \rf_reg[811] ;
 wire \rf_reg[812] ;
 wire \rf_reg[813] ;
 wire \rf_reg[814] ;
 wire \rf_reg[815] ;
 wire \rf_reg[816] ;
 wire \rf_reg[817] ;
 wire \rf_reg[818] ;
 wire \rf_reg[819] ;
 wire \rf_reg[81] ;
 wire \rf_reg[820] ;
 wire \rf_reg[821] ;
 wire \rf_reg[822] ;
 wire \rf_reg[823] ;
 wire \rf_reg[824] ;
 wire \rf_reg[825] ;
 wire \rf_reg[826] ;
 wire \rf_reg[827] ;
 wire \rf_reg[828] ;
 wire \rf_reg[829] ;
 wire \rf_reg[82] ;
 wire \rf_reg[830] ;
 wire \rf_reg[831] ;
 wire \rf_reg[832] ;
 wire \rf_reg[833] ;
 wire \rf_reg[834] ;
 wire \rf_reg[835] ;
 wire \rf_reg[836] ;
 wire \rf_reg[837] ;
 wire \rf_reg[838] ;
 wire \rf_reg[839] ;
 wire \rf_reg[83] ;
 wire \rf_reg[840] ;
 wire \rf_reg[841] ;
 wire \rf_reg[842] ;
 wire \rf_reg[843] ;
 wire \rf_reg[844] ;
 wire \rf_reg[845] ;
 wire \rf_reg[846] ;
 wire \rf_reg[847] ;
 wire \rf_reg[848] ;
 wire \rf_reg[849] ;
 wire \rf_reg[84] ;
 wire \rf_reg[850] ;
 wire \rf_reg[851] ;
 wire \rf_reg[852] ;
 wire \rf_reg[853] ;
 wire \rf_reg[854] ;
 wire \rf_reg[855] ;
 wire \rf_reg[856] ;
 wire \rf_reg[857] ;
 wire \rf_reg[858] ;
 wire \rf_reg[859] ;
 wire \rf_reg[85] ;
 wire \rf_reg[860] ;
 wire \rf_reg[861] ;
 wire \rf_reg[862] ;
 wire \rf_reg[863] ;
 wire \rf_reg[864] ;
 wire \rf_reg[865] ;
 wire \rf_reg[866] ;
 wire \rf_reg[867] ;
 wire \rf_reg[868] ;
 wire \rf_reg[869] ;
 wire \rf_reg[86] ;
 wire \rf_reg[870] ;
 wire \rf_reg[871] ;
 wire \rf_reg[872] ;
 wire \rf_reg[873] ;
 wire \rf_reg[874] ;
 wire \rf_reg[875] ;
 wire \rf_reg[876] ;
 wire \rf_reg[877] ;
 wire \rf_reg[878] ;
 wire \rf_reg[879] ;
 wire \rf_reg[87] ;
 wire \rf_reg[880] ;
 wire \rf_reg[881] ;
 wire \rf_reg[882] ;
 wire \rf_reg[883] ;
 wire \rf_reg[884] ;
 wire \rf_reg[885] ;
 wire \rf_reg[886] ;
 wire \rf_reg[887] ;
 wire \rf_reg[888] ;
 wire \rf_reg[889] ;
 wire \rf_reg[88] ;
 wire \rf_reg[890] ;
 wire \rf_reg[891] ;
 wire \rf_reg[892] ;
 wire \rf_reg[893] ;
 wire \rf_reg[894] ;
 wire \rf_reg[895] ;
 wire \rf_reg[896] ;
 wire \rf_reg[897] ;
 wire \rf_reg[898] ;
 wire \rf_reg[899] ;
 wire \rf_reg[89] ;
 wire \rf_reg[900] ;
 wire \rf_reg[901] ;
 wire \rf_reg[902] ;
 wire \rf_reg[903] ;
 wire \rf_reg[904] ;
 wire \rf_reg[905] ;
 wire \rf_reg[906] ;
 wire \rf_reg[907] ;
 wire \rf_reg[908] ;
 wire \rf_reg[909] ;
 wire \rf_reg[90] ;
 wire \rf_reg[910] ;
 wire \rf_reg[911] ;
 wire \rf_reg[912] ;
 wire \rf_reg[913] ;
 wire \rf_reg[914] ;
 wire \rf_reg[915] ;
 wire \rf_reg[916] ;
 wire \rf_reg[917] ;
 wire \rf_reg[918] ;
 wire \rf_reg[919] ;
 wire \rf_reg[91] ;
 wire \rf_reg[920] ;
 wire \rf_reg[921] ;
 wire \rf_reg[922] ;
 wire \rf_reg[923] ;
 wire \rf_reg[924] ;
 wire \rf_reg[925] ;
 wire \rf_reg[926] ;
 wire \rf_reg[927] ;
 wire \rf_reg[928] ;
 wire \rf_reg[929] ;
 wire \rf_reg[92] ;
 wire \rf_reg[930] ;
 wire \rf_reg[931] ;
 wire \rf_reg[932] ;
 wire \rf_reg[933] ;
 wire \rf_reg[934] ;
 wire \rf_reg[935] ;
 wire \rf_reg[936] ;
 wire \rf_reg[937] ;
 wire \rf_reg[938] ;
 wire \rf_reg[939] ;
 wire \rf_reg[93] ;
 wire \rf_reg[940] ;
 wire \rf_reg[941] ;
 wire \rf_reg[942] ;
 wire \rf_reg[943] ;
 wire \rf_reg[944] ;
 wire \rf_reg[945] ;
 wire \rf_reg[946] ;
 wire \rf_reg[947] ;
 wire \rf_reg[948] ;
 wire \rf_reg[949] ;
 wire \rf_reg[94] ;
 wire \rf_reg[950] ;
 wire \rf_reg[951] ;
 wire \rf_reg[952] ;
 wire \rf_reg[953] ;
 wire \rf_reg[954] ;
 wire \rf_reg[955] ;
 wire \rf_reg[956] ;
 wire \rf_reg[957] ;
 wire \rf_reg[958] ;
 wire \rf_reg[959] ;
 wire \rf_reg[95] ;
 wire \rf_reg[960] ;
 wire \rf_reg[961] ;
 wire \rf_reg[962] ;
 wire \rf_reg[963] ;
 wire \rf_reg[964] ;
 wire \rf_reg[965] ;
 wire \rf_reg[966] ;
 wire \rf_reg[967] ;
 wire \rf_reg[968] ;
 wire \rf_reg[969] ;
 wire \rf_reg[96] ;
 wire \rf_reg[970] ;
 wire \rf_reg[971] ;
 wire \rf_reg[972] ;
 wire \rf_reg[973] ;
 wire \rf_reg[974] ;
 wire \rf_reg[975] ;
 wire \rf_reg[976] ;
 wire \rf_reg[977] ;
 wire \rf_reg[978] ;
 wire \rf_reg[979] ;
 wire \rf_reg[97] ;
 wire \rf_reg[980] ;
 wire \rf_reg[981] ;
 wire \rf_reg[982] ;
 wire \rf_reg[983] ;
 wire \rf_reg[984] ;
 wire \rf_reg[985] ;
 wire \rf_reg[986] ;
 wire \rf_reg[987] ;
 wire \rf_reg[988] ;
 wire \rf_reg[989] ;
 wire \rf_reg[98] ;
 wire \rf_reg[990] ;
 wire \rf_reg[991] ;
 wire \rf_reg[992] ;
 wire \rf_reg[993] ;
 wire \rf_reg[994] ;
 wire \rf_reg[995] ;
 wire \rf_reg[996] ;
 wire \rf_reg[997] ;
 wire \rf_reg[998] ;
 wire \rf_reg[999] ;
 wire \rf_reg[99] ;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_leaf_39_clk_i;
 wire clknet_leaf_40_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_42_clk_i;
 wire clknet_leaf_43_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_45_clk_i;
 wire clknet_leaf_46_clk_i;
 wire clknet_leaf_47_clk_i;
 wire clknet_leaf_48_clk_i;
 wire clknet_leaf_49_clk_i;
 wire clknet_leaf_50_clk_i;
 wire clknet_leaf_51_clk_i;
 wire clknet_leaf_52_clk_i;
 wire clknet_leaf_53_clk_i;
 wire clknet_leaf_54_clk_i;
 wire clknet_leaf_55_clk_i;
 wire clknet_leaf_56_clk_i;
 wire clknet_leaf_57_clk_i;
 wire clknet_leaf_58_clk_i;
 wire clknet_leaf_59_clk_i;
 wire clknet_leaf_60_clk_i;
 wire clknet_leaf_61_clk_i;
 wire clknet_leaf_62_clk_i;
 wire clknet_leaf_63_clk_i;
 wire clknet_leaf_64_clk_i;
 wire clknet_leaf_65_clk_i;
 wire clknet_leaf_66_clk_i;
 wire clknet_leaf_67_clk_i;
 wire clknet_leaf_68_clk_i;
 wire clknet_leaf_69_clk_i;
 wire clknet_leaf_70_clk_i;
 wire clknet_leaf_71_clk_i;
 wire clknet_leaf_72_clk_i;
 wire clknet_leaf_73_clk_i;
 wire clknet_leaf_74_clk_i;
 wire clknet_leaf_75_clk_i;
 wire clknet_leaf_76_clk_i;
 wire clknet_leaf_77_clk_i;
 wire clknet_leaf_78_clk_i;
 wire clknet_leaf_79_clk_i;
 wire clknet_leaf_80_clk_i;
 wire clknet_leaf_81_clk_i;
 wire clknet_leaf_82_clk_i;
 wire clknet_leaf_83_clk_i;
 wire clknet_leaf_84_clk_i;
 wire clknet_leaf_85_clk_i;
 wire clknet_leaf_86_clk_i;
 wire clknet_leaf_87_clk_i;
 wire clknet_leaf_88_clk_i;
 wire clknet_leaf_89_clk_i;
 wire clknet_leaf_90_clk_i;
 wire clknet_leaf_91_clk_i;
 wire clknet_leaf_92_clk_i;
 wire clknet_leaf_93_clk_i;
 wire clknet_leaf_94_clk_i;
 wire clknet_leaf_95_clk_i;
 wire clknet_leaf_96_clk_i;
 wire clknet_leaf_97_clk_i;
 wire clknet_leaf_98_clk_i;
 wire clknet_leaf_99_clk_i;
 wire clknet_leaf_100_clk_i;
 wire clknet_leaf_101_clk_i;
 wire clknet_leaf_102_clk_i;
 wire clknet_leaf_103_clk_i;
 wire clknet_leaf_104_clk_i;
 wire clknet_leaf_105_clk_i;
 wire clknet_leaf_106_clk_i;
 wire clknet_leaf_107_clk_i;
 wire clknet_0_clk_i;
 wire clknet_3_0__leaf_clk_i;
 wire clknet_3_1__leaf_clk_i;
 wire clknet_3_2__leaf_clk_i;
 wire clknet_3_3__leaf_clk_i;
 wire clknet_3_4__leaf_clk_i;
 wire clknet_3_5__leaf_clk_i;
 wire clknet_3_6__leaf_clk_i;
 wire clknet_3_7__leaf_clk_i;

 sky130_fd_sc_hd__clkbuf_4 _2326_ (.A(net6),
    .X(_0992_));
 sky130_fd_sc_hd__buf_6 _2327_ (.A(net4),
    .X(_0993_));
 sky130_fd_sc_hd__buf_6 _2328_ (.A(net3),
    .X(_0994_));
 sky130_fd_sc_hd__nor2b_4 _2329_ (.A(_0993_),
    .B_N(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__buf_6 _2330_ (.A(waddr_a_i[3]),
    .X(_0996_));
 sky130_fd_sc_hd__buf_6 _2331_ (.A(waddr_a_i[2]),
    .X(_0997_));
 sky130_fd_sc_hd__nand2b_2 _2332_ (.A_N(net5),
    .B(net46),
    .Y(_0998_));
 sky130_fd_sc_hd__nor3_4 _2333_ (.A(_0996_),
    .B(_0997_),
    .C(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2_8 _2334_ (.A(_0995_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__buf_8 _2335_ (.A(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _2336_ (.A0(_0992_),
    .A1(\rf_reg[32] ),
    .S(_1001_),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _2337_ (.A(net40),
    .X(_1002_));
 sky130_fd_sc_hd__nor2_8 _2338_ (.A(_0993_),
    .B(_0994_),
    .Y(_1003_));
 sky130_fd_sc_hd__nor3b_4 _2339_ (.A(_0998_),
    .B(_0996_),
    .C_N(_0997_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand2_8 _2340_ (.A(_1003_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__buf_8 _2341_ (.A(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(_1002_),
    .A1(\rf_reg[132] ),
    .S(_1006_),
    .X(_0001_));
 sky130_fd_sc_hd__clkbuf_4 _2343_ (.A(net41),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _2344_ (.A0(_1007_),
    .A1(\rf_reg[133] ),
    .S(_1006_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _2345_ (.A(net42),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(_1008_),
    .A1(\rf_reg[134] ),
    .S(_1006_),
    .X(_0003_));
 sky130_fd_sc_hd__clkbuf_4 _2347_ (.A(net43),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _2348_ (.A0(_1009_),
    .A1(\rf_reg[135] ),
    .S(_1006_),
    .X(_0004_));
 sky130_fd_sc_hd__buf_2 _2349_ (.A(net44),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _2350_ (.A0(_1010_),
    .A1(\rf_reg[136] ),
    .S(_1006_),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_4 _2351_ (.A(net45),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_1 _2352_ (.A0(_1011_),
    .A1(\rf_reg[137] ),
    .S(_1006_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_4 _2353_ (.A(net7),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(_1012_),
    .A1(\rf_reg[138] ),
    .S(_1006_),
    .X(_0007_));
 sky130_fd_sc_hd__clkbuf_4 _2355_ (.A(net16),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _2356_ (.A0(_1013_),
    .A1(\rf_reg[139] ),
    .S(_1006_),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_4 _2357_ (.A(net17),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _2358_ (.A0(_1014_),
    .A1(\rf_reg[140] ),
    .S(_1006_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _2359_ (.A(net18),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_1 _2360_ (.A0(_1015_),
    .A1(\rf_reg[141] ),
    .S(_1006_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2361_ (.A0(_1012_),
    .A1(\rf_reg[42] ),
    .S(_1001_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_2 _2362_ (.A(net19),
    .X(_1016_));
 sky130_fd_sc_hd__buf_8 _2363_ (.A(_1005_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _2364_ (.A0(_1016_),
    .A1(\rf_reg[142] ),
    .S(_1017_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_4 _2365_ (.A(net20),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(_1018_),
    .A1(\rf_reg[143] ),
    .S(_1017_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _2367_ (.A(net21),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(_1019_),
    .A1(\rf_reg[144] ),
    .S(_1017_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _2369_ (.A(net22),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _2370_ (.A0(_1020_),
    .A1(\rf_reg[145] ),
    .S(_1017_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_4 _2371_ (.A(net23),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _2372_ (.A0(_1021_),
    .A1(\rf_reg[146] ),
    .S(_1017_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_4 _2373_ (.A(net24),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(_1022_),
    .A1(\rf_reg[147] ),
    .S(_1017_),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_4 _2375_ (.A(net26),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(_1023_),
    .A1(\rf_reg[148] ),
    .S(_1017_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _2377_ (.A(net27),
    .X(_1024_));
 sky130_fd_sc_hd__mux2_1 _2378_ (.A0(_1024_),
    .A1(\rf_reg[149] ),
    .S(_1017_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _2379_ (.A(net28),
    .X(_1025_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(_1025_),
    .A1(\rf_reg[150] ),
    .S(_1017_),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_4 _2381_ (.A(net29),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(_1026_),
    .A1(\rf_reg[151] ),
    .S(_1017_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(_1013_),
    .A1(\rf_reg[43] ),
    .S(_1001_),
    .X(_0022_));
 sky130_fd_sc_hd__buf_4 _2384_ (.A(net30),
    .X(_1027_));
 sky130_fd_sc_hd__buf_8 _2385_ (.A(_1005_),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(_1027_),
    .A1(\rf_reg[152] ),
    .S(_1028_),
    .X(_0023_));
 sky130_fd_sc_hd__buf_4 _2387_ (.A(net31),
    .X(_1029_));
 sky130_fd_sc_hd__mux2_1 _2388_ (.A0(_1029_),
    .A1(\rf_reg[153] ),
    .S(_1028_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_4 _2389_ (.A(net32),
    .X(_1030_));
 sky130_fd_sc_hd__mux2_1 _2390_ (.A0(_1030_),
    .A1(\rf_reg[154] ),
    .S(_1028_),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_4 _2391_ (.A(net33),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_1 _2392_ (.A0(_1031_),
    .A1(\rf_reg[155] ),
    .S(_1028_),
    .X(_0026_));
 sky130_fd_sc_hd__clkbuf_4 _2393_ (.A(net34),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _2394_ (.A0(_1032_),
    .A1(\rf_reg[156] ),
    .S(_1028_),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_4 _2395_ (.A(net35),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(_1033_),
    .A1(\rf_reg[157] ),
    .S(_1028_),
    .X(_0028_));
 sky130_fd_sc_hd__clkbuf_4 _2397_ (.A(net37),
    .X(_1034_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(_1034_),
    .A1(\rf_reg[158] ),
    .S(_1028_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_4 _2399_ (.A(net38),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _2400_ (.A0(_1035_),
    .A1(\rf_reg[159] ),
    .S(_1028_),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_4 _2401_ (.A(_0995_),
    .B(_1004_),
    .Y(_1036_));
 sky130_fd_sc_hd__buf_8 _2402_ (.A(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(_0992_),
    .A1(\rf_reg[160] ),
    .S(_1037_),
    .X(_0031_));
 sky130_fd_sc_hd__buf_2 _2404_ (.A(net25),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(_1038_),
    .A1(\rf_reg[161] ),
    .S(_1037_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2406_ (.A0(_1014_),
    .A1(\rf_reg[44] ),
    .S(_1001_),
    .X(_0033_));
 sky130_fd_sc_hd__buf_2 _2407_ (.A(net36),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _2408_ (.A0(_1039_),
    .A1(\rf_reg[162] ),
    .S(_1037_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_4 _2409_ (.A(net39),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _2410_ (.A0(_1040_),
    .A1(\rf_reg[163] ),
    .S(_1037_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(_1002_),
    .A1(\rf_reg[164] ),
    .S(_1037_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2412_ (.A0(_1007_),
    .A1(\rf_reg[165] ),
    .S(_1037_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(_1008_),
    .A1(\rf_reg[166] ),
    .S(_1037_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2414_ (.A0(_1009_),
    .A1(\rf_reg[167] ),
    .S(_1037_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(_1010_),
    .A1(\rf_reg[168] ),
    .S(_1037_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(_1011_),
    .A1(\rf_reg[169] ),
    .S(_1037_),
    .X(_0041_));
 sky130_fd_sc_hd__clkbuf_16 _2417_ (.A(_1036_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _2418_ (.A0(_1012_),
    .A1(\rf_reg[170] ),
    .S(_1041_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(_1013_),
    .A1(\rf_reg[171] ),
    .S(_1041_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(_1015_),
    .A1(\rf_reg[45] ),
    .S(_1001_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(_1014_),
    .A1(\rf_reg[172] ),
    .S(_1041_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(_1015_),
    .A1(\rf_reg[173] ),
    .S(_1041_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(_1016_),
    .A1(\rf_reg[174] ),
    .S(_1041_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2424_ (.A0(_1018_),
    .A1(\rf_reg[175] ),
    .S(_1041_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(_1019_),
    .A1(\rf_reg[176] ),
    .S(_1041_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(_1020_),
    .A1(\rf_reg[177] ),
    .S(_1041_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(_1021_),
    .A1(\rf_reg[178] ),
    .S(_1041_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2428_ (.A0(_1022_),
    .A1(\rf_reg[179] ),
    .S(_1041_),
    .X(_0052_));
 sky130_fd_sc_hd__buf_8 _2429_ (.A(_1036_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _2430_ (.A0(_1023_),
    .A1(\rf_reg[180] ),
    .S(_1042_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(_1024_),
    .A1(\rf_reg[181] ),
    .S(_1042_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2432_ (.A0(_1016_),
    .A1(\rf_reg[46] ),
    .S(_1001_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2433_ (.A0(_1025_),
    .A1(\rf_reg[182] ),
    .S(_1042_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(_1026_),
    .A1(\rf_reg[183] ),
    .S(_1042_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(_1027_),
    .A1(\rf_reg[184] ),
    .S(_1042_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(_1029_),
    .A1(\rf_reg[185] ),
    .S(_1042_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2437_ (.A0(_1030_),
    .A1(\rf_reg[186] ),
    .S(_1042_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(_1031_),
    .A1(\rf_reg[187] ),
    .S(_1042_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(_1032_),
    .A1(\rf_reg[188] ),
    .S(_1042_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(_1033_),
    .A1(\rf_reg[189] ),
    .S(_1042_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2441_ (.A0(_1034_),
    .A1(\rf_reg[190] ),
    .S(_1036_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2442_ (.A0(_1035_),
    .A1(\rf_reg[191] ),
    .S(_1036_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2443_ (.A0(_1018_),
    .A1(\rf_reg[47] ),
    .S(_1001_),
    .X(_0066_));
 sky130_fd_sc_hd__nor2b_4 _2444_ (.A(_0994_),
    .B_N(_0993_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_4 _2445_ (.A(_1004_),
    .B(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__buf_8 _2446_ (.A(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(_0992_),
    .A1(\rf_reg[192] ),
    .S(_1045_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2448_ (.A0(_1038_),
    .A1(\rf_reg[193] ),
    .S(_1045_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2449_ (.A0(_1039_),
    .A1(\rf_reg[194] ),
    .S(_1045_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(_1040_),
    .A1(\rf_reg[195] ),
    .S(_1045_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2451_ (.A0(_1002_),
    .A1(\rf_reg[196] ),
    .S(_1045_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2452_ (.A0(_1007_),
    .A1(\rf_reg[197] ),
    .S(_1045_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(_1008_),
    .A1(\rf_reg[198] ),
    .S(_1045_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2454_ (.A0(_1009_),
    .A1(\rf_reg[199] ),
    .S(_1045_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(_1010_),
    .A1(\rf_reg[200] ),
    .S(_1045_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2456_ (.A0(_1011_),
    .A1(\rf_reg[201] ),
    .S(_1045_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2457_ (.A0(_1019_),
    .A1(\rf_reg[48] ),
    .S(_1001_),
    .X(_0077_));
 sky130_fd_sc_hd__buf_8 _2458_ (.A(_1044_),
    .X(_1046_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(_1012_),
    .A1(\rf_reg[202] ),
    .S(_1046_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2460_ (.A0(_1013_),
    .A1(\rf_reg[203] ),
    .S(_1046_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2461_ (.A0(_1014_),
    .A1(\rf_reg[204] ),
    .S(_1046_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(_1015_),
    .A1(\rf_reg[205] ),
    .S(_1046_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2463_ (.A0(_1016_),
    .A1(\rf_reg[206] ),
    .S(_1046_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2464_ (.A0(_1018_),
    .A1(\rf_reg[207] ),
    .S(_1046_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2465_ (.A0(_1019_),
    .A1(\rf_reg[208] ),
    .S(_1046_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2466_ (.A0(_1020_),
    .A1(\rf_reg[209] ),
    .S(_1046_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(_1021_),
    .A1(\rf_reg[210] ),
    .S(_1046_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2468_ (.A0(_1022_),
    .A1(\rf_reg[211] ),
    .S(_1046_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(_1020_),
    .A1(\rf_reg[49] ),
    .S(_1001_),
    .X(_0088_));
 sky130_fd_sc_hd__buf_8 _2470_ (.A(_1044_),
    .X(_1047_));
 sky130_fd_sc_hd__mux2_1 _2471_ (.A0(_1023_),
    .A1(\rf_reg[212] ),
    .S(_1047_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2472_ (.A0(_1024_),
    .A1(\rf_reg[213] ),
    .S(_1047_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2473_ (.A0(_1025_),
    .A1(\rf_reg[214] ),
    .S(_1047_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(_1026_),
    .A1(\rf_reg[215] ),
    .S(_1047_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2475_ (.A0(_1027_),
    .A1(\rf_reg[216] ),
    .S(_1047_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(_1029_),
    .A1(\rf_reg[217] ),
    .S(_1047_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(_1030_),
    .A1(\rf_reg[218] ),
    .S(_1047_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(_1031_),
    .A1(\rf_reg[219] ),
    .S(_1047_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2479_ (.A0(_1032_),
    .A1(\rf_reg[220] ),
    .S(_1047_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2480_ (.A0(_1033_),
    .A1(\rf_reg[221] ),
    .S(_1047_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2481_ (.A0(_1021_),
    .A1(\rf_reg[50] ),
    .S(_1001_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(_1034_),
    .A1(\rf_reg[222] ),
    .S(_1044_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(_1035_),
    .A1(\rf_reg[223] ),
    .S(_1044_),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_4 _2484_ (.A(net6),
    .X(_1048_));
 sky130_fd_sc_hd__and3_1 _2485_ (.A(_0993_),
    .B(_0994_),
    .C(_1004_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_4 _2486_ (.A(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__buf_8 _2487_ (.A(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _2488_ (.A0(\rf_reg[224] ),
    .A1(_1048_),
    .S(_1051_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_4 _2489_ (.A(net25),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(\rf_reg[225] ),
    .A1(_1052_),
    .S(_1051_),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_4 _2491_ (.A(net36),
    .X(_1053_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(\rf_reg[226] ),
    .A1(_1053_),
    .S(_1051_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_4 _2493_ (.A(net39),
    .X(_1054_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(\rf_reg[227] ),
    .A1(_1054_),
    .S(_1051_),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_4 _2495_ (.A(net40),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(\rf_reg[228] ),
    .A1(_1055_),
    .S(_1051_),
    .X(_0106_));
 sky130_fd_sc_hd__buf_2 _2497_ (.A(net41),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(\rf_reg[229] ),
    .A1(_1056_),
    .S(_1051_),
    .X(_0107_));
 sky130_fd_sc_hd__buf_2 _2499_ (.A(net42),
    .X(_1057_));
 sky130_fd_sc_hd__mux2_1 _2500_ (.A0(\rf_reg[230] ),
    .A1(_1057_),
    .S(_1051_),
    .X(_0108_));
 sky130_fd_sc_hd__buf_2 _2501_ (.A(net43),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(\rf_reg[231] ),
    .A1(_1058_),
    .S(_1051_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_6 _2503_ (.A(_1000_),
    .X(_1059_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(_1022_),
    .A1(\rf_reg[51] ),
    .S(_1059_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(_1038_),
    .A1(\rf_reg[33] ),
    .S(_1059_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_4 _2506_ (.A(net44),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _2507_ (.A0(\rf_reg[232] ),
    .A1(_1060_),
    .S(_1051_),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_4 _2508_ (.A(net45),
    .X(_1061_));
 sky130_fd_sc_hd__mux2_1 _2509_ (.A0(\rf_reg[233] ),
    .A1(_1061_),
    .S(_1051_),
    .X(_0113_));
 sky130_fd_sc_hd__buf_4 _2510_ (.A(net7),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_16 _2511_ (.A(_1050_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(\rf_reg[234] ),
    .A1(_1062_),
    .S(_1063_),
    .X(_0114_));
 sky130_fd_sc_hd__buf_4 _2513_ (.A(net16),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(\rf_reg[235] ),
    .A1(_1064_),
    .S(_1063_),
    .X(_0115_));
 sky130_fd_sc_hd__buf_4 _2515_ (.A(net17),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(\rf_reg[236] ),
    .A1(_1065_),
    .S(_1063_),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_4 _2517_ (.A(net18),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(\rf_reg[237] ),
    .A1(_1066_),
    .S(_1063_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_4 _2519_ (.A(net19),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(\rf_reg[238] ),
    .A1(_1067_),
    .S(_1063_),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_4 _2521_ (.A(net20),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(\rf_reg[239] ),
    .A1(_1068_),
    .S(_1063_),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_4 _2523_ (.A(net21),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(\rf_reg[240] ),
    .A1(_1069_),
    .S(_1063_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_4 _2525_ (.A(net22),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\rf_reg[241] ),
    .A1(_1070_),
    .S(_1063_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(_1023_),
    .A1(\rf_reg[52] ),
    .S(_1059_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_4 _2528_ (.A(net23),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(\rf_reg[242] ),
    .A1(_1071_),
    .S(_1063_),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_4 _2530_ (.A(net24),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(\rf_reg[243] ),
    .A1(_1072_),
    .S(_1063_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_4 _2532_ (.A(net26),
    .X(_1073_));
 sky130_fd_sc_hd__buf_8 _2533_ (.A(_1050_),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(\rf_reg[244] ),
    .A1(_1073_),
    .S(_1074_),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_4 _2535_ (.A(net27),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(\rf_reg[245] ),
    .A1(_1075_),
    .S(_1074_),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_4 _2537_ (.A(net28),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\rf_reg[246] ),
    .A1(_1076_),
    .S(_1074_),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_4 _2539_ (.A(net29),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(\rf_reg[247] ),
    .A1(_1077_),
    .S(_1074_),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_4 _2541_ (.A(net30),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(\rf_reg[248] ),
    .A1(_1078_),
    .S(_1074_),
    .X(_0129_));
 sky130_fd_sc_hd__buf_4 _2543_ (.A(net31),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(\rf_reg[249] ),
    .A1(_1079_),
    .S(_1074_),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_4 _2545_ (.A(net32),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(\rf_reg[250] ),
    .A1(_1080_),
    .S(_1074_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_4 _2547_ (.A(net33),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(\rf_reg[251] ),
    .A1(_1081_),
    .S(_1074_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2549_ (.A0(_1024_),
    .A1(\rf_reg[53] ),
    .S(_1059_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_4 _2550_ (.A(net34),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(\rf_reg[252] ),
    .A1(_1082_),
    .S(_1074_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_4 _2552_ (.A(net35),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(\rf_reg[253] ),
    .A1(_1083_),
    .S(_1074_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_4 _2554_ (.A(net37),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(\rf_reg[254] ),
    .A1(_1084_),
    .S(_1050_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_4 _2556_ (.A(net38),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(\rf_reg[255] ),
    .A1(_1085_),
    .S(_1050_),
    .X(_0137_));
 sky130_fd_sc_hd__nor3b_4 _2558_ (.A(_0997_),
    .B(_0998_),
    .C_N(_0996_),
    .Y(_1086_));
 sky130_fd_sc_hd__nand2_8 _2559_ (.A(_1003_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__buf_16 _2560_ (.A(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(_0992_),
    .A1(\rf_reg[256] ),
    .S(_1088_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(_1038_),
    .A1(\rf_reg[257] ),
    .S(_1088_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(_1039_),
    .A1(\rf_reg[258] ),
    .S(_1088_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2564_ (.A0(_1040_),
    .A1(\rf_reg[259] ),
    .S(_1088_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(_1002_),
    .A1(\rf_reg[260] ),
    .S(_1088_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(_1007_),
    .A1(\rf_reg[261] ),
    .S(_1088_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(_1025_),
    .A1(\rf_reg[54] ),
    .S(_1059_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2568_ (.A0(_1008_),
    .A1(\rf_reg[262] ),
    .S(_1088_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(_1009_),
    .A1(\rf_reg[263] ),
    .S(_1088_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(_1010_),
    .A1(\rf_reg[264] ),
    .S(_1088_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(_1011_),
    .A1(\rf_reg[265] ),
    .S(_1088_),
    .X(_0148_));
 sky130_fd_sc_hd__buf_16 _2572_ (.A(_1087_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(_1012_),
    .A1(\rf_reg[266] ),
    .S(_1089_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(_1013_),
    .A1(\rf_reg[267] ),
    .S(_1089_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(_1014_),
    .A1(\rf_reg[268] ),
    .S(_1089_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(_1015_),
    .A1(\rf_reg[269] ),
    .S(_1089_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2577_ (.A0(_1016_),
    .A1(\rf_reg[270] ),
    .S(_1089_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(_1018_),
    .A1(\rf_reg[271] ),
    .S(_1089_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(_1026_),
    .A1(\rf_reg[55] ),
    .S(_1059_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(_1019_),
    .A1(\rf_reg[272] ),
    .S(_1089_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2581_ (.A0(_1020_),
    .A1(\rf_reg[273] ),
    .S(_1089_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(_1021_),
    .A1(\rf_reg[274] ),
    .S(_1089_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(_1022_),
    .A1(\rf_reg[275] ),
    .S(_1089_),
    .X(_0159_));
 sky130_fd_sc_hd__buf_8 _2584_ (.A(_1087_),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(_1023_),
    .A1(\rf_reg[276] ),
    .S(_1090_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(_1024_),
    .A1(\rf_reg[277] ),
    .S(_1090_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(_1025_),
    .A1(\rf_reg[278] ),
    .S(_1090_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(_1026_),
    .A1(\rf_reg[279] ),
    .S(_1090_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(_1027_),
    .A1(\rf_reg[280] ),
    .S(_1090_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(_1029_),
    .A1(\rf_reg[281] ),
    .S(_1090_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(_1027_),
    .A1(\rf_reg[56] ),
    .S(_1059_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(_1030_),
    .A1(\rf_reg[282] ),
    .S(_1090_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(_1031_),
    .A1(\rf_reg[283] ),
    .S(_1090_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2594_ (.A0(_1032_),
    .A1(\rf_reg[284] ),
    .S(_1090_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(_1033_),
    .A1(\rf_reg[285] ),
    .S(_1090_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(_1034_),
    .A1(\rf_reg[286] ),
    .S(_1087_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(_1035_),
    .A1(\rf_reg[287] ),
    .S(_1087_),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_4 _2598_ (.A(_0995_),
    .B(_1086_),
    .Y(_1091_));
 sky130_fd_sc_hd__clkbuf_16 _2599_ (.A(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(_0992_),
    .A1(\rf_reg[288] ),
    .S(_1092_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(_1038_),
    .A1(\rf_reg[289] ),
    .S(_1092_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(_1039_),
    .A1(\rf_reg[290] ),
    .S(_1092_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(_1040_),
    .A1(\rf_reg[291] ),
    .S(_1092_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(_1029_),
    .A1(\rf_reg[57] ),
    .S(_1059_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2605_ (.A0(_1002_),
    .A1(\rf_reg[292] ),
    .S(_1092_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2606_ (.A0(_1007_),
    .A1(\rf_reg[293] ),
    .S(_1092_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(_1008_),
    .A1(\rf_reg[294] ),
    .S(_1092_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2608_ (.A0(_1009_),
    .A1(\rf_reg[295] ),
    .S(_1092_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(_1010_),
    .A1(\rf_reg[296] ),
    .S(_1092_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(_1011_),
    .A1(\rf_reg[297] ),
    .S(_1092_),
    .X(_0183_));
 sky130_fd_sc_hd__buf_12 _2611_ (.A(_1091_),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(_1012_),
    .A1(\rf_reg[298] ),
    .S(_1093_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(_1013_),
    .A1(\rf_reg[299] ),
    .S(_1093_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2614_ (.A0(_1014_),
    .A1(\rf_reg[300] ),
    .S(_1093_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(_1015_),
    .A1(\rf_reg[301] ),
    .S(_1093_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2616_ (.A0(_1030_),
    .A1(\rf_reg[58] ),
    .S(_1059_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(_1016_),
    .A1(\rf_reg[302] ),
    .S(_1093_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2618_ (.A0(_1018_),
    .A1(\rf_reg[303] ),
    .S(_1093_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(_1019_),
    .A1(\rf_reg[304] ),
    .S(_1093_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2620_ (.A0(_1020_),
    .A1(\rf_reg[305] ),
    .S(_1093_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2621_ (.A0(_1021_),
    .A1(\rf_reg[306] ),
    .S(_1093_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2622_ (.A0(_1022_),
    .A1(\rf_reg[307] ),
    .S(_1093_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_16 _2623_ (.A(_1091_),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(_1023_),
    .A1(\rf_reg[308] ),
    .S(_1094_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(_1024_),
    .A1(\rf_reg[309] ),
    .S(_1094_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(_1025_),
    .A1(\rf_reg[310] ),
    .S(_1094_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(_1026_),
    .A1(\rf_reg[311] ),
    .S(_1094_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(_1031_),
    .A1(\rf_reg[59] ),
    .S(_1059_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2629_ (.A0(_1027_),
    .A1(\rf_reg[312] ),
    .S(_1094_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(_1029_),
    .A1(\rf_reg[313] ),
    .S(_1094_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(_1030_),
    .A1(\rf_reg[314] ),
    .S(_1094_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(_1031_),
    .A1(\rf_reg[315] ),
    .S(_1094_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2633_ (.A0(_1032_),
    .A1(\rf_reg[316] ),
    .S(_1094_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(_1033_),
    .A1(\rf_reg[317] ),
    .S(_1094_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2635_ (.A0(_1034_),
    .A1(\rf_reg[318] ),
    .S(_1091_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(_1035_),
    .A1(\rf_reg[319] ),
    .S(_1091_),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_8 _2637_ (.A(_1043_),
    .B(_1086_),
    .Y(_1095_));
 sky130_fd_sc_hd__buf_8 _2638_ (.A(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(_0992_),
    .A1(\rf_reg[320] ),
    .S(_1096_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(_1038_),
    .A1(\rf_reg[321] ),
    .S(_1096_),
    .X(_0209_));
 sky130_fd_sc_hd__buf_6 _2641_ (.A(_1000_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(_1032_),
    .A1(\rf_reg[60] ),
    .S(_1097_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(_1039_),
    .A1(\rf_reg[322] ),
    .S(_1096_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(_1040_),
    .A1(\rf_reg[323] ),
    .S(_1096_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(_1002_),
    .A1(\rf_reg[324] ),
    .S(_1096_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(_1007_),
    .A1(\rf_reg[325] ),
    .S(_1096_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(_1008_),
    .A1(\rf_reg[326] ),
    .S(_1096_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(_1009_),
    .A1(\rf_reg[327] ),
    .S(_1096_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(_1010_),
    .A1(\rf_reg[328] ),
    .S(_1096_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(_1011_),
    .A1(\rf_reg[329] ),
    .S(_1096_),
    .X(_0218_));
 sky130_fd_sc_hd__buf_12 _2651_ (.A(_1095_),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(_1012_),
    .A1(\rf_reg[330] ),
    .S(_1098_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(_1013_),
    .A1(\rf_reg[331] ),
    .S(_1098_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2654_ (.A0(_1033_),
    .A1(\rf_reg[61] ),
    .S(_1097_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(_1039_),
    .A1(\rf_reg[34] ),
    .S(_1097_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(_1014_),
    .A1(\rf_reg[332] ),
    .S(_1098_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(_1015_),
    .A1(\rf_reg[333] ),
    .S(_1098_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(_1016_),
    .A1(\rf_reg[334] ),
    .S(_1098_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(_1018_),
    .A1(\rf_reg[335] ),
    .S(_1098_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(_1019_),
    .A1(\rf_reg[336] ),
    .S(_1098_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(_1020_),
    .A1(\rf_reg[337] ),
    .S(_1098_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(_1021_),
    .A1(\rf_reg[338] ),
    .S(_1098_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(_1022_),
    .A1(\rf_reg[339] ),
    .S(_1098_),
    .X(_0230_));
 sky130_fd_sc_hd__buf_8 _2664_ (.A(_1095_),
    .X(_1099_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(_1023_),
    .A1(\rf_reg[340] ),
    .S(_1099_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(_1024_),
    .A1(\rf_reg[341] ),
    .S(_1099_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(_1034_),
    .A1(\rf_reg[62] ),
    .S(_1097_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2668_ (.A0(_1025_),
    .A1(\rf_reg[342] ),
    .S(_1099_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2669_ (.A0(_1026_),
    .A1(\rf_reg[343] ),
    .S(_1099_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(_1027_),
    .A1(\rf_reg[344] ),
    .S(_1099_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2671_ (.A0(_1029_),
    .A1(\rf_reg[345] ),
    .S(_1099_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(_1030_),
    .A1(\rf_reg[346] ),
    .S(_1099_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2673_ (.A0(_1031_),
    .A1(\rf_reg[347] ),
    .S(_1099_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(_1032_),
    .A1(\rf_reg[348] ),
    .S(_1099_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(_1033_),
    .A1(\rf_reg[349] ),
    .S(_1099_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(_1034_),
    .A1(\rf_reg[350] ),
    .S(_1095_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2677_ (.A0(_1035_),
    .A1(\rf_reg[351] ),
    .S(_1095_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2678_ (.A0(_1035_),
    .A1(\rf_reg[63] ),
    .S(_1097_),
    .X(_0244_));
 sky130_fd_sc_hd__nand2_8 _2679_ (.A(net4),
    .B(net3),
    .Y(_1100_));
 sky130_fd_sc_hd__nor2b_1 _2680_ (.A(_1100_),
    .B_N(_1086_),
    .Y(_1101_));
 sky130_fd_sc_hd__buf_6 _2681_ (.A(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__buf_16 _2682_ (.A(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _2683_ (.A0(\rf_reg[352] ),
    .A1(_1048_),
    .S(_1103_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(\rf_reg[353] ),
    .A1(_1052_),
    .S(_1103_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2685_ (.A0(\rf_reg[354] ),
    .A1(_1053_),
    .S(_1103_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(\rf_reg[355] ),
    .A1(_1054_),
    .S(_1103_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _2687_ (.A0(\rf_reg[356] ),
    .A1(_1055_),
    .S(_1103_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(\rf_reg[357] ),
    .A1(_1056_),
    .S(_1103_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _2689_ (.A0(\rf_reg[358] ),
    .A1(_1057_),
    .S(_1103_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(\rf_reg[359] ),
    .A1(_1058_),
    .S(_1103_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _2691_ (.A0(\rf_reg[360] ),
    .A1(_1060_),
    .S(_1103_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(\rf_reg[361] ),
    .A1(_1061_),
    .S(_1103_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_4 _2693_ (.A(_0999_),
    .B(_1043_),
    .Y(_1104_));
 sky130_fd_sc_hd__buf_8 _2694_ (.A(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _2695_ (.A0(_0992_),
    .A1(\rf_reg[64] ),
    .S(_1105_),
    .X(_0255_));
 sky130_fd_sc_hd__buf_16 _2696_ (.A(_1102_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _2697_ (.A0(\rf_reg[362] ),
    .A1(_1062_),
    .S(_1106_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(\rf_reg[363] ),
    .A1(_1064_),
    .S(_1106_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(\rf_reg[364] ),
    .A1(_1065_),
    .S(_1106_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(\rf_reg[365] ),
    .A1(_1066_),
    .S(_1106_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(\rf_reg[366] ),
    .A1(_1067_),
    .S(_1106_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2702_ (.A0(\rf_reg[367] ),
    .A1(_1068_),
    .S(_1106_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(\rf_reg[368] ),
    .A1(_1069_),
    .S(_1106_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _2704_ (.A0(\rf_reg[369] ),
    .A1(_1070_),
    .S(_1106_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(\rf_reg[370] ),
    .A1(_1071_),
    .S(_1106_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _2706_ (.A0(\rf_reg[371] ),
    .A1(_1072_),
    .S(_1106_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _2707_ (.A0(_1038_),
    .A1(\rf_reg[65] ),
    .S(_1105_),
    .X(_0266_));
 sky130_fd_sc_hd__buf_16 _2708_ (.A(_1102_),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(\rf_reg[372] ),
    .A1(_1073_),
    .S(_1107_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _2710_ (.A0(\rf_reg[373] ),
    .A1(_1075_),
    .S(_1107_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(\rf_reg[374] ),
    .A1(_1076_),
    .S(_1107_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _2712_ (.A0(\rf_reg[375] ),
    .A1(_1077_),
    .S(_1107_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(\rf_reg[376] ),
    .A1(_1078_),
    .S(_1107_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _2714_ (.A0(\rf_reg[377] ),
    .A1(_1079_),
    .S(_1107_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(\rf_reg[378] ),
    .A1(_1080_),
    .S(_1107_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(\rf_reg[379] ),
    .A1(_1081_),
    .S(_1107_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(\rf_reg[380] ),
    .A1(_1082_),
    .S(_1107_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(\rf_reg[381] ),
    .A1(_1083_),
    .S(_1107_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(_1039_),
    .A1(\rf_reg[66] ),
    .S(_1105_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2720_ (.A0(\rf_reg[382] ),
    .A1(_1084_),
    .S(_1102_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(\rf_reg[383] ),
    .A1(_1085_),
    .S(_1102_),
    .X(_0279_));
 sky130_fd_sc_hd__nand4b_4 _2722_ (.A_N(net5),
    .B(net46),
    .C(_0996_),
    .D(_0997_),
    .Y(_1108_));
 sky130_fd_sc_hd__or3_1 _2723_ (.A(_0993_),
    .B(_0994_),
    .C(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__buf_4 _2724_ (.A(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_16 _2725_ (.A(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(_0992_),
    .A1(\rf_reg[384] ),
    .S(_1111_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(_1038_),
    .A1(\rf_reg[385] ),
    .S(_1111_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(_1039_),
    .A1(\rf_reg[386] ),
    .S(_1111_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(_1040_),
    .A1(\rf_reg[387] ),
    .S(_1111_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(_1002_),
    .A1(\rf_reg[388] ),
    .S(_1111_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2731_ (.A0(_1007_),
    .A1(\rf_reg[389] ),
    .S(_1111_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(_1008_),
    .A1(\rf_reg[390] ),
    .S(_1111_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(_1009_),
    .A1(\rf_reg[391] ),
    .S(_1111_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(_1040_),
    .A1(\rf_reg[67] ),
    .S(_1105_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(_1010_),
    .A1(\rf_reg[392] ),
    .S(_1111_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(_1011_),
    .A1(\rf_reg[393] ),
    .S(_1111_),
    .X(_0290_));
 sky130_fd_sc_hd__buf_12 _2737_ (.A(_1110_),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(_1012_),
    .A1(\rf_reg[394] ),
    .S(_1112_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(_1013_),
    .A1(\rf_reg[395] ),
    .S(_1112_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(_1014_),
    .A1(\rf_reg[396] ),
    .S(_1112_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(_1015_),
    .A1(\rf_reg[397] ),
    .S(_1112_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(_1016_),
    .A1(\rf_reg[398] ),
    .S(_1112_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _2743_ (.A0(_1018_),
    .A1(\rf_reg[399] ),
    .S(_1112_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(_1019_),
    .A1(\rf_reg[400] ),
    .S(_1112_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(_1020_),
    .A1(\rf_reg[401] ),
    .S(_1112_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(_1002_),
    .A1(\rf_reg[68] ),
    .S(_1105_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(_1021_),
    .A1(\rf_reg[402] ),
    .S(_1112_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(_1022_),
    .A1(\rf_reg[403] ),
    .S(_1112_),
    .X(_0301_));
 sky130_fd_sc_hd__buf_16 _2749_ (.A(_1110_),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _2750_ (.A0(_1023_),
    .A1(\rf_reg[404] ),
    .S(_1113_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(_1024_),
    .A1(\rf_reg[405] ),
    .S(_1113_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(_1025_),
    .A1(\rf_reg[406] ),
    .S(_1113_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(_1026_),
    .A1(\rf_reg[407] ),
    .S(_1113_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(_1027_),
    .A1(\rf_reg[408] ),
    .S(_1113_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(_1029_),
    .A1(\rf_reg[409] ),
    .S(_1113_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _2756_ (.A0(_1030_),
    .A1(\rf_reg[410] ),
    .S(_1113_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(_1031_),
    .A1(\rf_reg[411] ),
    .S(_1113_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2758_ (.A0(_1007_),
    .A1(\rf_reg[69] ),
    .S(_1105_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(_1032_),
    .A1(\rf_reg[412] ),
    .S(_1113_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2760_ (.A0(_1033_),
    .A1(\rf_reg[413] ),
    .S(_1113_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(_1034_),
    .A1(\rf_reg[414] ),
    .S(_1110_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2762_ (.A0(_1035_),
    .A1(\rf_reg[415] ),
    .S(_1110_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2b_4 _2763_ (.A_N(_0993_),
    .B(_0994_),
    .Y(_1114_));
 sky130_fd_sc_hd__nor2_8 _2764_ (.A(_1114_),
    .B(_1108_),
    .Y(_1115_));
 sky130_fd_sc_hd__buf_12 _2765_ (.A(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(\rf_reg[416] ),
    .A1(_1048_),
    .S(_1116_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _2767_ (.A0(\rf_reg[417] ),
    .A1(_1052_),
    .S(_1116_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2768_ (.A0(\rf_reg[418] ),
    .A1(_1053_),
    .S(_1116_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(\rf_reg[419] ),
    .A1(_1054_),
    .S(_1116_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2770_ (.A0(\rf_reg[420] ),
    .A1(_1055_),
    .S(_1116_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2771_ (.A0(\rf_reg[421] ),
    .A1(_1056_),
    .S(_1116_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(_1008_),
    .A1(\rf_reg[70] ),
    .S(_1105_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(\rf_reg[422] ),
    .A1(_1057_),
    .S(_1116_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2774_ (.A0(\rf_reg[423] ),
    .A1(_1058_),
    .S(_1116_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(\rf_reg[424] ),
    .A1(_1060_),
    .S(_1116_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _2776_ (.A0(\rf_reg[425] ),
    .A1(_1061_),
    .S(_1116_),
    .X(_0325_));
 sky130_fd_sc_hd__buf_12 _2777_ (.A(_1115_),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _2778_ (.A0(\rf_reg[426] ),
    .A1(_1062_),
    .S(_1117_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(\rf_reg[427] ),
    .A1(_1064_),
    .S(_1117_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _2780_ (.A0(\rf_reg[428] ),
    .A1(_1065_),
    .S(_1117_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\rf_reg[429] ),
    .A1(_1066_),
    .S(_1117_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2782_ (.A0(\rf_reg[430] ),
    .A1(_1067_),
    .S(_1117_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(\rf_reg[431] ),
    .A1(_1068_),
    .S(_1117_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(_1009_),
    .A1(\rf_reg[71] ),
    .S(_1105_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(_1040_),
    .A1(\rf_reg[35] ),
    .S(_1097_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _2786_ (.A0(\rf_reg[432] ),
    .A1(_1069_),
    .S(_1117_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _2787_ (.A0(\rf_reg[433] ),
    .A1(_1070_),
    .S(_1117_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _2788_ (.A0(\rf_reg[434] ),
    .A1(_1071_),
    .S(_1117_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(\rf_reg[435] ),
    .A1(_1072_),
    .S(_1117_),
    .X(_0337_));
 sky130_fd_sc_hd__buf_16 _2790_ (.A(_1115_),
    .X(_1118_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(\rf_reg[436] ),
    .A1(_1073_),
    .S(_1118_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(\rf_reg[437] ),
    .A1(_1075_),
    .S(_1118_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _2793_ (.A0(\rf_reg[438] ),
    .A1(_1076_),
    .S(_1118_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(\rf_reg[439] ),
    .A1(_1077_),
    .S(_1118_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _2795_ (.A0(\rf_reg[440] ),
    .A1(_1078_),
    .S(_1118_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(\rf_reg[441] ),
    .A1(_1079_),
    .S(_1118_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(_1010_),
    .A1(\rf_reg[72] ),
    .S(_1105_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _2798_ (.A0(\rf_reg[442] ),
    .A1(_1080_),
    .S(_1118_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _2799_ (.A0(\rf_reg[443] ),
    .A1(_1081_),
    .S(_1118_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(\rf_reg[444] ),
    .A1(_1082_),
    .S(_1118_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _2801_ (.A0(\rf_reg[445] ),
    .A1(_1083_),
    .S(_1118_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(\rf_reg[446] ),
    .A1(_1084_),
    .S(_1115_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(\rf_reg[447] ),
    .A1(_1085_),
    .S(_1115_),
    .X(_0350_));
 sky130_fd_sc_hd__nand2b_4 _2804_ (.A_N(_0994_),
    .B(_0993_),
    .Y(_1119_));
 sky130_fd_sc_hd__nor2_8 _2805_ (.A(_1119_),
    .B(_1108_),
    .Y(_1120_));
 sky130_fd_sc_hd__buf_16 _2806_ (.A(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__mux2_1 _2807_ (.A0(\rf_reg[448] ),
    .A1(_1048_),
    .S(_1121_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(\rf_reg[449] ),
    .A1(_1052_),
    .S(_1121_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(\rf_reg[450] ),
    .A1(_1053_),
    .S(_1121_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(\rf_reg[451] ),
    .A1(_1054_),
    .S(_1121_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(_1011_),
    .A1(\rf_reg[73] ),
    .S(_1105_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(\rf_reg[452] ),
    .A1(_1055_),
    .S(_1121_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(\rf_reg[453] ),
    .A1(_1056_),
    .S(_1121_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _2814_ (.A0(\rf_reg[454] ),
    .A1(_1057_),
    .S(_1121_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(\rf_reg[455] ),
    .A1(_1058_),
    .S(_1121_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _2816_ (.A0(\rf_reg[456] ),
    .A1(_1060_),
    .S(_1121_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(\rf_reg[457] ),
    .A1(_1061_),
    .S(_1121_),
    .X(_0361_));
 sky130_fd_sc_hd__buf_12 _2818_ (.A(_1120_),
    .X(_1122_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(\rf_reg[458] ),
    .A1(_1062_),
    .S(_1122_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _2820_ (.A0(\rf_reg[459] ),
    .A1(_1064_),
    .S(_1122_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(\rf_reg[460] ),
    .A1(_1065_),
    .S(_1122_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _2822_ (.A0(\rf_reg[461] ),
    .A1(_1066_),
    .S(_1122_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_8 _2823_ (.A(_1104_),
    .X(_1123_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(_1012_),
    .A1(\rf_reg[74] ),
    .S(_1123_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _2825_ (.A0(\rf_reg[462] ),
    .A1(_1067_),
    .S(_1122_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(\rf_reg[463] ),
    .A1(_1068_),
    .S(_1122_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(\rf_reg[464] ),
    .A1(_1069_),
    .S(_1122_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(\rf_reg[465] ),
    .A1(_1070_),
    .S(_1122_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _2829_ (.A0(\rf_reg[466] ),
    .A1(_1071_),
    .S(_1122_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _2830_ (.A0(\rf_reg[467] ),
    .A1(_1072_),
    .S(_1122_),
    .X(_0372_));
 sky130_fd_sc_hd__buf_8 _2831_ (.A(_1120_),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_1 _2832_ (.A0(\rf_reg[468] ),
    .A1(_1073_),
    .S(_1124_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _2833_ (.A0(\rf_reg[469] ),
    .A1(_1075_),
    .S(_1124_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _2834_ (.A0(\rf_reg[470] ),
    .A1(_1076_),
    .S(_1124_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(\rf_reg[471] ),
    .A1(_1077_),
    .S(_1124_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(_1013_),
    .A1(\rf_reg[75] ),
    .S(_1123_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(\rf_reg[472] ),
    .A1(_1078_),
    .S(_1124_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(\rf_reg[473] ),
    .A1(_1079_),
    .S(_1124_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(\rf_reg[474] ),
    .A1(_1080_),
    .S(_1124_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _2840_ (.A0(\rf_reg[475] ),
    .A1(_1081_),
    .S(_1124_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(\rf_reg[476] ),
    .A1(_1082_),
    .S(_1124_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(\rf_reg[477] ),
    .A1(_1083_),
    .S(_1124_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _2843_ (.A0(\rf_reg[478] ),
    .A1(_1084_),
    .S(_1120_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(\rf_reg[479] ),
    .A1(_1085_),
    .S(_1120_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_8 _2845_ (.A(_1100_),
    .B(_1108_),
    .Y(_1125_));
 sky130_fd_sc_hd__buf_16 _2846_ (.A(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_1 _2847_ (.A0(\rf_reg[480] ),
    .A1(_1048_),
    .S(_1126_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(\rf_reg[481] ),
    .A1(_1052_),
    .S(_1126_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(_1014_),
    .A1(\rf_reg[76] ),
    .S(_1123_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _2850_ (.A0(\rf_reg[482] ),
    .A1(_1053_),
    .S(_1126_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\rf_reg[483] ),
    .A1(_1054_),
    .S(_1126_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(\rf_reg[484] ),
    .A1(_1055_),
    .S(_1126_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(\rf_reg[485] ),
    .A1(_1056_),
    .S(_1126_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _2854_ (.A0(\rf_reg[486] ),
    .A1(_1057_),
    .S(_1126_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(\rf_reg[487] ),
    .A1(_1058_),
    .S(_1126_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(\rf_reg[488] ),
    .A1(_1060_),
    .S(_1126_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\rf_reg[489] ),
    .A1(_1061_),
    .S(_1126_),
    .X(_0396_));
 sky130_fd_sc_hd__buf_12 _2858_ (.A(_1125_),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(\rf_reg[490] ),
    .A1(_1062_),
    .S(_1127_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(\rf_reg[491] ),
    .A1(_1064_),
    .S(_1127_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _2861_ (.A0(_1015_),
    .A1(\rf_reg[77] ),
    .S(_1123_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(\rf_reg[492] ),
    .A1(_1065_),
    .S(_1127_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(\rf_reg[493] ),
    .A1(_1066_),
    .S(_1127_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(\rf_reg[494] ),
    .A1(_1067_),
    .S(_1127_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(\rf_reg[495] ),
    .A1(_1068_),
    .S(_1127_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _2866_ (.A0(\rf_reg[496] ),
    .A1(_1069_),
    .S(_1127_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(\rf_reg[497] ),
    .A1(_1070_),
    .S(_1127_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(\rf_reg[498] ),
    .A1(_1071_),
    .S(_1127_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _2869_ (.A0(\rf_reg[499] ),
    .A1(_1072_),
    .S(_1127_),
    .X(_0407_));
 sky130_fd_sc_hd__buf_16 _2870_ (.A(_1125_),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(\rf_reg[500] ),
    .A1(_1073_),
    .S(_1128_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(\rf_reg[501] ),
    .A1(_1075_),
    .S(_1128_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _2873_ (.A0(_1016_),
    .A1(\rf_reg[78] ),
    .S(_1123_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\rf_reg[502] ),
    .A1(_1076_),
    .S(_1128_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _2875_ (.A0(\rf_reg[503] ),
    .A1(_1077_),
    .S(_1128_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\rf_reg[504] ),
    .A1(_1078_),
    .S(_1128_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _2877_ (.A0(\rf_reg[505] ),
    .A1(_1079_),
    .S(_1128_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(\rf_reg[506] ),
    .A1(_1080_),
    .S(_1128_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _2879_ (.A0(\rf_reg[507] ),
    .A1(_1081_),
    .S(_1128_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _2880_ (.A0(\rf_reg[508] ),
    .A1(_1082_),
    .S(_1128_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _2881_ (.A0(\rf_reg[509] ),
    .A1(_1083_),
    .S(_1128_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(\rf_reg[510] ),
    .A1(_1084_),
    .S(_1125_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _2883_ (.A0(\rf_reg[511] ),
    .A1(_1085_),
    .S(_1125_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(_1018_),
    .A1(\rf_reg[79] ),
    .S(_1123_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_2 _2885_ (.A(net5),
    .B(net46),
    .Y(_1129_));
 sky130_fd_sc_hd__nor3_4 _2886_ (.A(_0996_),
    .B(_0997_),
    .C(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand2_8 _2887_ (.A(_1003_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__clkbuf_16 _2888_ (.A(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(_0992_),
    .A1(\rf_reg[512] ),
    .S(_1132_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(_1038_),
    .A1(\rf_reg[513] ),
    .S(_1132_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(_1039_),
    .A1(\rf_reg[514] ),
    .S(_1132_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _2892_ (.A0(_1040_),
    .A1(\rf_reg[515] ),
    .S(_1132_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _2893_ (.A0(_1002_),
    .A1(\rf_reg[516] ),
    .S(_1132_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(_1007_),
    .A1(\rf_reg[517] ),
    .S(_1132_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _2895_ (.A0(_1008_),
    .A1(\rf_reg[518] ),
    .S(_1132_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(_1009_),
    .A1(\rf_reg[519] ),
    .S(_1132_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(_1010_),
    .A1(\rf_reg[520] ),
    .S(_1132_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(_1011_),
    .A1(\rf_reg[521] ),
    .S(_1132_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(_1019_),
    .A1(\rf_reg[80] ),
    .S(_1123_),
    .X(_0432_));
 sky130_fd_sc_hd__buf_8 _2900_ (.A(_1131_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(_1012_),
    .A1(\rf_reg[522] ),
    .S(_1133_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(_1013_),
    .A1(\rf_reg[523] ),
    .S(_1133_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(_1014_),
    .A1(\rf_reg[524] ),
    .S(_1133_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _2904_ (.A0(_1015_),
    .A1(\rf_reg[525] ),
    .S(_1133_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(_1016_),
    .A1(\rf_reg[526] ),
    .S(_1133_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _2906_ (.A0(_1018_),
    .A1(\rf_reg[527] ),
    .S(_1133_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(_1019_),
    .A1(\rf_reg[528] ),
    .S(_1133_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _2908_ (.A0(_1020_),
    .A1(\rf_reg[529] ),
    .S(_1133_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(_1021_),
    .A1(\rf_reg[530] ),
    .S(_1133_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _2910_ (.A0(_1022_),
    .A1(\rf_reg[531] ),
    .S(_1133_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(_1020_),
    .A1(\rf_reg[81] ),
    .S(_1123_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _2912_ (.A0(_1002_),
    .A1(\rf_reg[36] ),
    .S(_1097_),
    .X(_0444_));
 sky130_fd_sc_hd__buf_16 _2913_ (.A(_1131_),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _2914_ (.A0(_1023_),
    .A1(\rf_reg[532] ),
    .S(_1134_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(_1024_),
    .A1(\rf_reg[533] ),
    .S(_1134_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(_1025_),
    .A1(\rf_reg[534] ),
    .S(_1134_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _2917_ (.A0(_1026_),
    .A1(\rf_reg[535] ),
    .S(_1134_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(_1027_),
    .A1(\rf_reg[536] ),
    .S(_1134_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _2919_ (.A0(_1029_),
    .A1(\rf_reg[537] ),
    .S(_1134_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(_1030_),
    .A1(\rf_reg[538] ),
    .S(_1134_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(_1031_),
    .A1(\rf_reg[539] ),
    .S(_1134_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(_1032_),
    .A1(\rf_reg[540] ),
    .S(_1134_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(_1033_),
    .A1(\rf_reg[541] ),
    .S(_1134_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _2924_ (.A0(_1021_),
    .A1(\rf_reg[82] ),
    .S(_1123_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _2925_ (.A0(_1034_),
    .A1(\rf_reg[542] ),
    .S(_1131_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _2926_ (.A0(_1035_),
    .A1(\rf_reg[543] ),
    .S(_1131_),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_8 _2927_ (.A(_0995_),
    .B(_1130_),
    .Y(_1135_));
 sky130_fd_sc_hd__clkbuf_16 _2928_ (.A(_1135_),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(_0992_),
    .A1(\rf_reg[544] ),
    .S(_1136_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _2930_ (.A0(_1038_),
    .A1(\rf_reg[545] ),
    .S(_1136_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _2931_ (.A0(_1039_),
    .A1(\rf_reg[546] ),
    .S(_1136_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(_1040_),
    .A1(\rf_reg[547] ),
    .S(_1136_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _2933_ (.A0(_1055_),
    .A1(\rf_reg[548] ),
    .S(_1136_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _2934_ (.A0(_1007_),
    .A1(\rf_reg[549] ),
    .S(_1136_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _2935_ (.A0(_1008_),
    .A1(\rf_reg[550] ),
    .S(_1136_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _2936_ (.A0(_1009_),
    .A1(\rf_reg[551] ),
    .S(_1136_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _2937_ (.A0(_1022_),
    .A1(\rf_reg[83] ),
    .S(_1123_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(_1010_),
    .A1(\rf_reg[552] ),
    .S(_1136_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _2939_ (.A0(_1011_),
    .A1(\rf_reg[553] ),
    .S(_1136_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_8 _2940_ (.A(_1135_),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(_1062_),
    .A1(\rf_reg[554] ),
    .S(_1137_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(_1064_),
    .A1(\rf_reg[555] ),
    .S(_1137_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _2943_ (.A0(_1065_),
    .A1(\rf_reg[556] ),
    .S(_1137_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _2944_ (.A0(_1066_),
    .A1(\rf_reg[557] ),
    .S(_1137_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _2945_ (.A0(_1067_),
    .A1(\rf_reg[558] ),
    .S(_1137_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _2946_ (.A0(_1068_),
    .A1(\rf_reg[559] ),
    .S(_1137_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(_1069_),
    .A1(\rf_reg[560] ),
    .S(_1137_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _2948_ (.A0(_1070_),
    .A1(\rf_reg[561] ),
    .S(_1137_),
    .X(_0476_));
 sky130_fd_sc_hd__buf_8 _2949_ (.A(_1104_),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(_1023_),
    .A1(\rf_reg[84] ),
    .S(_1138_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(_1071_),
    .A1(\rf_reg[562] ),
    .S(_1137_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _2952_ (.A0(_1072_),
    .A1(\rf_reg[563] ),
    .S(_1137_),
    .X(_0479_));
 sky130_fd_sc_hd__buf_16 _2953_ (.A(_1135_),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _2954_ (.A0(_1073_),
    .A1(\rf_reg[564] ),
    .S(_1139_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _2955_ (.A0(_1024_),
    .A1(\rf_reg[565] ),
    .S(_1139_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(_1025_),
    .A1(\rf_reg[566] ),
    .S(_1139_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(_1026_),
    .A1(\rf_reg[567] ),
    .S(_1139_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(_1027_),
    .A1(\rf_reg[568] ),
    .S(_1139_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(_1029_),
    .A1(\rf_reg[569] ),
    .S(_1139_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _2960_ (.A0(_1030_),
    .A1(\rf_reg[570] ),
    .S(_1139_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(_1031_),
    .A1(\rf_reg[571] ),
    .S(_1139_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(_1075_),
    .A1(\rf_reg[85] ),
    .S(_1138_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _2963_ (.A0(_1032_),
    .A1(\rf_reg[572] ),
    .S(_1139_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(_1033_),
    .A1(\rf_reg[573] ),
    .S(_1139_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(_1034_),
    .A1(\rf_reg[574] ),
    .S(_1135_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(_1035_),
    .A1(\rf_reg[575] ),
    .S(_1135_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_8 _2967_ (.A(_1043_),
    .B(_1130_),
    .Y(_1140_));
 sky130_fd_sc_hd__buf_16 _2968_ (.A(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(_1048_),
    .A1(\rf_reg[576] ),
    .S(_1141_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(_1052_),
    .A1(\rf_reg[577] ),
    .S(_1141_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(_1053_),
    .A1(\rf_reg[578] ),
    .S(_1141_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _2972_ (.A0(_1054_),
    .A1(\rf_reg[579] ),
    .S(_1141_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(_1055_),
    .A1(\rf_reg[580] ),
    .S(_1141_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(_1056_),
    .A1(\rf_reg[581] ),
    .S(_1141_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _2975_ (.A0(_1076_),
    .A1(\rf_reg[86] ),
    .S(_1138_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(_1057_),
    .A1(\rf_reg[582] ),
    .S(_1141_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _2977_ (.A0(_1058_),
    .A1(\rf_reg[583] ),
    .S(_1141_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(_1060_),
    .A1(\rf_reg[584] ),
    .S(_1141_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _2979_ (.A0(_1061_),
    .A1(\rf_reg[585] ),
    .S(_1141_),
    .X(_0503_));
 sky130_fd_sc_hd__buf_8 _2980_ (.A(_1140_),
    .X(_1142_));
 sky130_fd_sc_hd__mux2_1 _2981_ (.A0(_1062_),
    .A1(\rf_reg[586] ),
    .S(_1142_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(_1064_),
    .A1(\rf_reg[587] ),
    .S(_1142_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(_1065_),
    .A1(\rf_reg[588] ),
    .S(_1142_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(_1066_),
    .A1(\rf_reg[589] ),
    .S(_1142_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(_1067_),
    .A1(\rf_reg[590] ),
    .S(_1142_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(_1068_),
    .A1(\rf_reg[591] ),
    .S(_1142_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(_1077_),
    .A1(\rf_reg[87] ),
    .S(_1138_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(_1069_),
    .A1(\rf_reg[592] ),
    .S(_1142_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(_1070_),
    .A1(\rf_reg[593] ),
    .S(_1142_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(_1071_),
    .A1(\rf_reg[594] ),
    .S(_1142_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(_1072_),
    .A1(\rf_reg[595] ),
    .S(_1142_),
    .X(_0514_));
 sky130_fd_sc_hd__buf_8 _2992_ (.A(_1140_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(_1073_),
    .A1(\rf_reg[596] ),
    .S(_1143_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(_1075_),
    .A1(\rf_reg[597] ),
    .S(_1143_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _2995_ (.A0(_1076_),
    .A1(\rf_reg[598] ),
    .S(_1143_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(_1077_),
    .A1(\rf_reg[599] ),
    .S(_1143_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(_1078_),
    .A1(\rf_reg[600] ),
    .S(_1143_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(_1079_),
    .A1(\rf_reg[601] ),
    .S(_1143_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(_1078_),
    .A1(\rf_reg[88] ),
    .S(_1138_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _3000_ (.A0(_1080_),
    .A1(\rf_reg[602] ),
    .S(_1143_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(_1081_),
    .A1(\rf_reg[603] ),
    .S(_1143_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(_1082_),
    .A1(\rf_reg[604] ),
    .S(_1143_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(_1083_),
    .A1(\rf_reg[605] ),
    .S(_1143_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3004_ (.A0(_1084_),
    .A1(\rf_reg[606] ),
    .S(_1140_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(_1085_),
    .A1(\rf_reg[607] ),
    .S(_1140_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _3006_ (.A(net6),
    .X(_1144_));
 sky130_fd_sc_hd__nor4_4 _3007_ (.A(_0996_),
    .B(_0997_),
    .C(_1100_),
    .D(_1129_),
    .Y(_1145_));
 sky130_fd_sc_hd__clkbuf_16 _3008_ (.A(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(\rf_reg[608] ),
    .A1(_1144_),
    .S(_1146_),
    .X(_0528_));
 sky130_fd_sc_hd__buf_2 _3010_ (.A(net25),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(\rf_reg[609] ),
    .A1(_1147_),
    .S(_1146_),
    .X(_0529_));
 sky130_fd_sc_hd__buf_2 _3012_ (.A(net36),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(\rf_reg[610] ),
    .A1(_1148_),
    .S(_1146_),
    .X(_0530_));
 sky130_fd_sc_hd__buf_2 _3014_ (.A(net39),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _3015_ (.A0(\rf_reg[611] ),
    .A1(_1149_),
    .S(_1146_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(_1079_),
    .A1(\rf_reg[89] ),
    .S(_1138_),
    .X(_0532_));
 sky130_fd_sc_hd__buf_2 _3017_ (.A(net40),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(\rf_reg[612] ),
    .A1(_1150_),
    .S(_1146_),
    .X(_0533_));
 sky130_fd_sc_hd__buf_2 _3019_ (.A(net41),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(\rf_reg[613] ),
    .A1(_1151_),
    .S(_1146_),
    .X(_0534_));
 sky130_fd_sc_hd__buf_2 _3021_ (.A(net42),
    .X(_1152_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(\rf_reg[614] ),
    .A1(_1152_),
    .S(_1146_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_2 _3023_ (.A(net43),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(\rf_reg[615] ),
    .A1(_1153_),
    .S(_1146_),
    .X(_0536_));
 sky130_fd_sc_hd__buf_2 _3025_ (.A(net44),
    .X(_1154_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(\rf_reg[616] ),
    .A1(_1154_),
    .S(_1146_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_2 _3027_ (.A(net45),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(\rf_reg[617] ),
    .A1(_1155_),
    .S(_1146_),
    .X(_0538_));
 sky130_fd_sc_hd__buf_2 _3029_ (.A(net7),
    .X(_1156_));
 sky130_fd_sc_hd__buf_6 _3030_ (.A(_1145_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _3031_ (.A0(\rf_reg[618] ),
    .A1(_1156_),
    .S(_1157_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_4 _3032_ (.A(net16),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _3033_ (.A0(\rf_reg[619] ),
    .A1(_1158_),
    .S(_1157_),
    .X(_0540_));
 sky130_fd_sc_hd__clkbuf_4 _3034_ (.A(net17),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_1 _3035_ (.A0(\rf_reg[620] ),
    .A1(_1159_),
    .S(_1157_),
    .X(_0541_));
 sky130_fd_sc_hd__buf_2 _3036_ (.A(net18),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(\rf_reg[621] ),
    .A1(_1160_),
    .S(_1157_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(_1080_),
    .A1(\rf_reg[90] ),
    .S(_1138_),
    .X(_0543_));
 sky130_fd_sc_hd__buf_2 _3039_ (.A(net19),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(\rf_reg[622] ),
    .A1(_1161_),
    .S(_1157_),
    .X(_0544_));
 sky130_fd_sc_hd__clkbuf_4 _3041_ (.A(net20),
    .X(_1162_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(\rf_reg[623] ),
    .A1(_1162_),
    .S(_1157_),
    .X(_0545_));
 sky130_fd_sc_hd__buf_2 _3043_ (.A(net21),
    .X(_1163_));
 sky130_fd_sc_hd__mux2_1 _3044_ (.A0(\rf_reg[624] ),
    .A1(_1163_),
    .S(_1157_),
    .X(_0546_));
 sky130_fd_sc_hd__buf_2 _3045_ (.A(net22),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _3046_ (.A0(\rf_reg[625] ),
    .A1(_1164_),
    .S(_1157_),
    .X(_0547_));
 sky130_fd_sc_hd__buf_2 _3047_ (.A(net23),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(\rf_reg[626] ),
    .A1(_1165_),
    .S(_1157_),
    .X(_0548_));
 sky130_fd_sc_hd__buf_2 _3049_ (.A(net24),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(\rf_reg[627] ),
    .A1(_1166_),
    .S(_1157_),
    .X(_0549_));
 sky130_fd_sc_hd__buf_2 _3051_ (.A(net26),
    .X(_1167_));
 sky130_fd_sc_hd__buf_16 _3052_ (.A(_1145_),
    .X(_1168_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(\rf_reg[628] ),
    .A1(_1167_),
    .S(_1168_),
    .X(_0550_));
 sky130_fd_sc_hd__buf_2 _3054_ (.A(net27),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(\rf_reg[629] ),
    .A1(_1169_),
    .S(_1168_),
    .X(_0551_));
 sky130_fd_sc_hd__buf_2 _3056_ (.A(net28),
    .X(_1170_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(\rf_reg[630] ),
    .A1(_1170_),
    .S(_1168_),
    .X(_0552_));
 sky130_fd_sc_hd__buf_2 _3058_ (.A(net29),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(\rf_reg[631] ),
    .A1(_1171_),
    .S(_1168_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(_1081_),
    .A1(\rf_reg[91] ),
    .S(_1138_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(_1056_),
    .A1(\rf_reg[37] ),
    .S(_1097_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _3062_ (.A(net30),
    .X(_1172_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(\rf_reg[632] ),
    .A1(_1172_),
    .S(_1168_),
    .X(_0556_));
 sky130_fd_sc_hd__buf_2 _3064_ (.A(net31),
    .X(_1173_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(\rf_reg[633] ),
    .A1(_1173_),
    .S(_1168_),
    .X(_0557_));
 sky130_fd_sc_hd__buf_2 _3066_ (.A(net32),
    .X(_1174_));
 sky130_fd_sc_hd__mux2_1 _3067_ (.A0(\rf_reg[634] ),
    .A1(_1174_),
    .S(_1168_),
    .X(_0558_));
 sky130_fd_sc_hd__buf_2 _3068_ (.A(net33),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(\rf_reg[635] ),
    .A1(_1175_),
    .S(_1168_),
    .X(_0559_));
 sky130_fd_sc_hd__buf_2 _3070_ (.A(net34),
    .X(_1176_));
 sky130_fd_sc_hd__mux2_1 _3071_ (.A0(\rf_reg[636] ),
    .A1(_1176_),
    .S(_1168_),
    .X(_0560_));
 sky130_fd_sc_hd__buf_2 _3072_ (.A(net35),
    .X(_1177_));
 sky130_fd_sc_hd__mux2_1 _3073_ (.A0(\rf_reg[637] ),
    .A1(_1177_),
    .S(_1168_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_4 _3074_ (.A(net37),
    .X(_1178_));
 sky130_fd_sc_hd__mux2_1 _3075_ (.A0(\rf_reg[638] ),
    .A1(_1178_),
    .S(_1145_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_4 _3076_ (.A(net38),
    .X(_1179_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(\rf_reg[639] ),
    .A1(_1179_),
    .S(_1145_),
    .X(_0563_));
 sky130_fd_sc_hd__nand4b_4 _3078_ (.A_N(_0996_),
    .B(_0997_),
    .C(net5),
    .D(net46),
    .Y(_1180_));
 sky130_fd_sc_hd__or3_1 _3079_ (.A(_0993_),
    .B(_0994_),
    .C(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__buf_6 _3080_ (.A(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__buf_16 _3081_ (.A(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(_1048_),
    .A1(\rf_reg[640] ),
    .S(_1183_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(_1052_),
    .A1(\rf_reg[641] ),
    .S(_1183_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(_1082_),
    .A1(\rf_reg[92] ),
    .S(_1138_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(_1053_),
    .A1(\rf_reg[642] ),
    .S(_1183_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(_1054_),
    .A1(\rf_reg[643] ),
    .S(_1183_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(_1055_),
    .A1(\rf_reg[644] ),
    .S(_1183_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _3088_ (.A0(_1056_),
    .A1(\rf_reg[645] ),
    .S(_1183_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(_1057_),
    .A1(\rf_reg[646] ),
    .S(_1183_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(_1058_),
    .A1(\rf_reg[647] ),
    .S(_1183_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(_1060_),
    .A1(\rf_reg[648] ),
    .S(_1183_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _3092_ (.A0(_1061_),
    .A1(\rf_reg[649] ),
    .S(_1183_),
    .X(_0574_));
 sky130_fd_sc_hd__buf_8 _3093_ (.A(_1182_),
    .X(_1184_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(_1062_),
    .A1(\rf_reg[650] ),
    .S(_1184_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(_1064_),
    .A1(\rf_reg[651] ),
    .S(_1184_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(_1083_),
    .A1(\rf_reg[93] ),
    .S(_1138_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(_1065_),
    .A1(\rf_reg[652] ),
    .S(_1184_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _3098_ (.A0(_1066_),
    .A1(\rf_reg[653] ),
    .S(_1184_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_1067_),
    .A1(\rf_reg[654] ),
    .S(_1184_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(_1068_),
    .A1(\rf_reg[655] ),
    .S(_1184_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1069_),
    .A1(\rf_reg[656] ),
    .S(_1184_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _3102_ (.A0(_1070_),
    .A1(\rf_reg[657] ),
    .S(_1184_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_1071_),
    .A1(\rf_reg[658] ),
    .S(_1184_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(_1072_),
    .A1(\rf_reg[659] ),
    .S(_1184_),
    .X(_0585_));
 sky130_fd_sc_hd__buf_16 _3105_ (.A(_1182_),
    .X(_1185_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(_1073_),
    .A1(\rf_reg[660] ),
    .S(_1185_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(_1075_),
    .A1(\rf_reg[661] ),
    .S(_1185_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(_1084_),
    .A1(\rf_reg[94] ),
    .S(_1104_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(_1076_),
    .A1(\rf_reg[662] ),
    .S(_1185_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(_1077_),
    .A1(\rf_reg[663] ),
    .S(_1185_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(_1078_),
    .A1(\rf_reg[664] ),
    .S(_1185_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(_1079_),
    .A1(\rf_reg[665] ),
    .S(_1185_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _3113_ (.A0(_1080_),
    .A1(\rf_reg[666] ),
    .S(_1185_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(_1081_),
    .A1(\rf_reg[667] ),
    .S(_1185_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(_1082_),
    .A1(\rf_reg[668] ),
    .S(_1185_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(_1083_),
    .A1(\rf_reg[669] ),
    .S(_1185_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(_1084_),
    .A1(\rf_reg[670] ),
    .S(_1182_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(_1085_),
    .A1(\rf_reg[671] ),
    .S(_1182_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(_1085_),
    .A1(\rf_reg[95] ),
    .S(_1104_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_8 _3120_ (.A(_1114_),
    .B(_1180_),
    .Y(_1186_));
 sky130_fd_sc_hd__buf_16 _3121_ (.A(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(\rf_reg[672] ),
    .A1(_1144_),
    .S(_1187_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(\rf_reg[673] ),
    .A1(_1147_),
    .S(_1187_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _3124_ (.A0(\rf_reg[674] ),
    .A1(_1148_),
    .S(_1187_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(\rf_reg[675] ),
    .A1(_1149_),
    .S(_1187_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(\rf_reg[676] ),
    .A1(_1150_),
    .S(_1187_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(\rf_reg[677] ),
    .A1(_1151_),
    .S(_1187_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(\rf_reg[678] ),
    .A1(_1152_),
    .S(_1187_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(\rf_reg[679] ),
    .A1(_1153_),
    .S(_1187_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(\rf_reg[680] ),
    .A1(_1154_),
    .S(_1187_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _3131_ (.A0(\rf_reg[681] ),
    .A1(_1155_),
    .S(_1187_),
    .X(_0609_));
 sky130_fd_sc_hd__nand3_4 _3132_ (.A(_0993_),
    .B(_0994_),
    .C(_0999_),
    .Y(_1188_));
 sky130_fd_sc_hd__buf_8 _3133_ (.A(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(_1048_),
    .A1(\rf_reg[96] ),
    .S(_1189_),
    .X(_0610_));
 sky130_fd_sc_hd__buf_8 _3135_ (.A(_1186_),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_1 _3136_ (.A0(\rf_reg[682] ),
    .A1(_1156_),
    .S(_1190_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(\rf_reg[683] ),
    .A1(_1158_),
    .S(_1190_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _3138_ (.A0(\rf_reg[684] ),
    .A1(_1159_),
    .S(_1190_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(\rf_reg[685] ),
    .A1(_1160_),
    .S(_1190_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _3140_ (.A0(\rf_reg[686] ),
    .A1(_1161_),
    .S(_1190_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _3141_ (.A0(\rf_reg[687] ),
    .A1(_1162_),
    .S(_1190_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _3142_ (.A0(\rf_reg[688] ),
    .A1(_1163_),
    .S(_1190_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _3143_ (.A0(\rf_reg[689] ),
    .A1(_1164_),
    .S(_1190_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(\rf_reg[690] ),
    .A1(_1165_),
    .S(_1190_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(\rf_reg[691] ),
    .A1(_1166_),
    .S(_1190_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(_1052_),
    .A1(\rf_reg[97] ),
    .S(_1189_),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_16 _3147_ (.A(_1186_),
    .X(_1191_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(\rf_reg[692] ),
    .A1(_1167_),
    .S(_1191_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(\rf_reg[693] ),
    .A1(_1169_),
    .S(_1191_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(\rf_reg[694] ),
    .A1(_1170_),
    .S(_1191_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _3151_ (.A0(\rf_reg[695] ),
    .A1(_1171_),
    .S(_1191_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(\rf_reg[696] ),
    .A1(_1172_),
    .S(_1191_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(\rf_reg[697] ),
    .A1(_1173_),
    .S(_1191_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(\rf_reg[698] ),
    .A1(_1174_),
    .S(_1191_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(\rf_reg[699] ),
    .A1(_1175_),
    .S(_1191_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(\rf_reg[700] ),
    .A1(_1176_),
    .S(_1191_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(\rf_reg[701] ),
    .A1(_1177_),
    .S(_1191_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(_1053_),
    .A1(\rf_reg[98] ),
    .S(_1189_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(\rf_reg[702] ),
    .A1(_1178_),
    .S(_1186_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(\rf_reg[703] ),
    .A1(_1179_),
    .S(_1186_),
    .X(_0634_));
 sky130_fd_sc_hd__nor2_8 _3161_ (.A(_1119_),
    .B(_1180_),
    .Y(_1192_));
 sky130_fd_sc_hd__buf_16 _3162_ (.A(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(\rf_reg[704] ),
    .A1(_1144_),
    .S(_1193_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(\rf_reg[705] ),
    .A1(_1147_),
    .S(_1193_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(\rf_reg[706] ),
    .A1(_1148_),
    .S(_1193_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _3166_ (.A0(\rf_reg[707] ),
    .A1(_1149_),
    .S(_1193_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(\rf_reg[708] ),
    .A1(_1150_),
    .S(_1193_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _3168_ (.A0(\rf_reg[709] ),
    .A1(_1151_),
    .S(_1193_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(\rf_reg[710] ),
    .A1(_1152_),
    .S(_1193_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _3170_ (.A0(\rf_reg[711] ),
    .A1(_1153_),
    .S(_1193_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(_1054_),
    .A1(\rf_reg[99] ),
    .S(_1189_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _3172_ (.A0(\rf_reg[712] ),
    .A1(_1154_),
    .S(_1193_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(\rf_reg[713] ),
    .A1(_1155_),
    .S(_1193_),
    .X(_0645_));
 sky130_fd_sc_hd__buf_8 _3174_ (.A(_1192_),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(\rf_reg[714] ),
    .A1(_1156_),
    .S(_1194_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _3176_ (.A0(\rf_reg[715] ),
    .A1(_1158_),
    .S(_1194_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(\rf_reg[716] ),
    .A1(_1159_),
    .S(_1194_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(\rf_reg[717] ),
    .A1(_1160_),
    .S(_1194_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(\rf_reg[718] ),
    .A1(_1161_),
    .S(_1194_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(\rf_reg[719] ),
    .A1(_1162_),
    .S(_1194_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(\rf_reg[720] ),
    .A1(_1163_),
    .S(_1194_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(\rf_reg[721] ),
    .A1(_1164_),
    .S(_1194_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(_1055_),
    .A1(\rf_reg[100] ),
    .S(_1189_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(\rf_reg[722] ),
    .A1(_1165_),
    .S(_1194_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(\rf_reg[723] ),
    .A1(_1166_),
    .S(_1194_),
    .X(_0656_));
 sky130_fd_sc_hd__buf_16 _3186_ (.A(_1192_),
    .X(_1195_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(\rf_reg[724] ),
    .A1(_1167_),
    .S(_1195_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(\rf_reg[725] ),
    .A1(_1169_),
    .S(_1195_),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(\rf_reg[726] ),
    .A1(_1170_),
    .S(_1195_),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(\rf_reg[727] ),
    .A1(_1171_),
    .S(_1195_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(\rf_reg[728] ),
    .A1(_1172_),
    .S(_1195_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(\rf_reg[729] ),
    .A1(_1173_),
    .S(_1195_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(\rf_reg[730] ),
    .A1(_1174_),
    .S(_1195_),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(\rf_reg[731] ),
    .A1(_1175_),
    .S(_1195_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(_1056_),
    .A1(\rf_reg[101] ),
    .S(_1189_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(_1057_),
    .A1(\rf_reg[38] ),
    .S(_1097_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _3197_ (.A0(\rf_reg[732] ),
    .A1(_1176_),
    .S(_1195_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(\rf_reg[733] ),
    .A1(_1177_),
    .S(_1195_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _3199_ (.A0(\rf_reg[734] ),
    .A1(_1178_),
    .S(_1192_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(\rf_reg[735] ),
    .A1(_1179_),
    .S(_1192_),
    .X(_0670_));
 sky130_fd_sc_hd__nor2_8 _3201_ (.A(_1100_),
    .B(_1180_),
    .Y(_1196_));
 sky130_fd_sc_hd__buf_16 _3202_ (.A(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(\rf_reg[736] ),
    .A1(_1144_),
    .S(_1197_),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(\rf_reg[737] ),
    .A1(_1147_),
    .S(_1197_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(\rf_reg[738] ),
    .A1(_1148_),
    .S(_1197_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(\rf_reg[739] ),
    .A1(_1149_),
    .S(_1197_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(\rf_reg[740] ),
    .A1(_1150_),
    .S(_1197_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(\rf_reg[741] ),
    .A1(_1151_),
    .S(_1197_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(_1057_),
    .A1(\rf_reg[102] ),
    .S(_1189_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _3210_ (.A0(\rf_reg[742] ),
    .A1(_1152_),
    .S(_1197_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(\rf_reg[743] ),
    .A1(_1153_),
    .S(_1197_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(\rf_reg[744] ),
    .A1(_1154_),
    .S(_1197_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(\rf_reg[745] ),
    .A1(_1155_),
    .S(_1197_),
    .X(_0681_));
 sky130_fd_sc_hd__buf_8 _3214_ (.A(_1196_),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\rf_reg[746] ),
    .A1(_1156_),
    .S(_1198_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(\rf_reg[747] ),
    .A1(_1158_),
    .S(_1198_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(\rf_reg[748] ),
    .A1(_1159_),
    .S(_1198_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(\rf_reg[749] ),
    .A1(_1160_),
    .S(_1198_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(\rf_reg[750] ),
    .A1(_1161_),
    .S(_1198_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(\rf_reg[751] ),
    .A1(_1162_),
    .S(_1198_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(_1058_),
    .A1(\rf_reg[103] ),
    .S(_1189_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(\rf_reg[752] ),
    .A1(_1163_),
    .S(_1198_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(\rf_reg[753] ),
    .A1(_1164_),
    .S(_1198_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(\rf_reg[754] ),
    .A1(_1165_),
    .S(_1198_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(\rf_reg[755] ),
    .A1(_1166_),
    .S(_1198_),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_16 _3226_ (.A(_1196_),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(\rf_reg[756] ),
    .A1(_1167_),
    .S(_1199_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(\rf_reg[757] ),
    .A1(_1169_),
    .S(_1199_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(\rf_reg[758] ),
    .A1(_1170_),
    .S(_1199_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(\rf_reg[759] ),
    .A1(_1171_),
    .S(_1199_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(\rf_reg[760] ),
    .A1(_1172_),
    .S(_1199_),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(\rf_reg[761] ),
    .A1(_1173_),
    .S(_1199_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(_1060_),
    .A1(\rf_reg[104] ),
    .S(_1189_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(\rf_reg[762] ),
    .A1(_1174_),
    .S(_1199_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _3235_ (.A0(\rf_reg[763] ),
    .A1(_1175_),
    .S(_1199_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(\rf_reg[764] ),
    .A1(_1176_),
    .S(_1199_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(\rf_reg[765] ),
    .A1(_1177_),
    .S(_1199_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(\rf_reg[766] ),
    .A1(_1178_),
    .S(_1196_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(\rf_reg[767] ),
    .A1(_1179_),
    .S(_1196_),
    .X(_0705_));
 sky130_fd_sc_hd__nand4b_4 _3240_ (.A_N(_0997_),
    .B(net5),
    .C(net46),
    .D(_0996_),
    .Y(_1200_));
 sky130_fd_sc_hd__or3_1 _3241_ (.A(net4),
    .B(net3),
    .C(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__buf_6 _3242_ (.A(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__buf_16 _3243_ (.A(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(_1048_),
    .A1(\rf_reg[768] ),
    .S(_1203_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(_1052_),
    .A1(\rf_reg[769] ),
    .S(_1203_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(_1053_),
    .A1(\rf_reg[770] ),
    .S(_1203_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(_1054_),
    .A1(\rf_reg[771] ),
    .S(_1203_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(_1061_),
    .A1(\rf_reg[105] ),
    .S(_1189_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(_1055_),
    .A1(\rf_reg[772] ),
    .S(_1203_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(_1056_),
    .A1(\rf_reg[773] ),
    .S(_1203_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(_1057_),
    .A1(\rf_reg[774] ),
    .S(_1203_),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(_1058_),
    .A1(\rf_reg[775] ),
    .S(_1203_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(_1060_),
    .A1(\rf_reg[776] ),
    .S(_1203_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(_1061_),
    .A1(\rf_reg[777] ),
    .S(_1203_),
    .X(_0716_));
 sky130_fd_sc_hd__buf_8 _3255_ (.A(_1202_),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(_1062_),
    .A1(\rf_reg[778] ),
    .S(_1204_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(_1064_),
    .A1(\rf_reg[779] ),
    .S(_1204_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(_1065_),
    .A1(\rf_reg[780] ),
    .S(_1204_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _3259_ (.A0(_1066_),
    .A1(\rf_reg[781] ),
    .S(_1204_),
    .X(_0720_));
 sky130_fd_sc_hd__clkbuf_16 _3260_ (.A(_1188_),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(_1062_),
    .A1(\rf_reg[106] ),
    .S(_1205_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(_1067_),
    .A1(\rf_reg[782] ),
    .S(_1204_),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(_1068_),
    .A1(\rf_reg[783] ),
    .S(_1204_),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(_1069_),
    .A1(\rf_reg[784] ),
    .S(_1204_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(_1070_),
    .A1(\rf_reg[785] ),
    .S(_1204_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(_1071_),
    .A1(\rf_reg[786] ),
    .S(_1204_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(_1072_),
    .A1(\rf_reg[787] ),
    .S(_1204_),
    .X(_0727_));
 sky130_fd_sc_hd__buf_16 _3268_ (.A(_1202_),
    .X(_1206_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(_1073_),
    .A1(\rf_reg[788] ),
    .S(_1206_),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(_1075_),
    .A1(\rf_reg[789] ),
    .S(_1206_),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(_1076_),
    .A1(\rf_reg[790] ),
    .S(_1206_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _3272_ (.A0(_1077_),
    .A1(\rf_reg[791] ),
    .S(_1206_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(_1064_),
    .A1(\rf_reg[107] ),
    .S(_1205_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(_1078_),
    .A1(\rf_reg[792] ),
    .S(_1206_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(_1079_),
    .A1(\rf_reg[793] ),
    .S(_1206_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(_1080_),
    .A1(\rf_reg[794] ),
    .S(_1206_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _3277_ (.A0(_1081_),
    .A1(\rf_reg[795] ),
    .S(_1206_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(_1082_),
    .A1(\rf_reg[796] ),
    .S(_1206_),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(_1083_),
    .A1(\rf_reg[797] ),
    .S(_1206_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(_1084_),
    .A1(\rf_reg[798] ),
    .S(_1202_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(_1085_),
    .A1(\rf_reg[799] ),
    .S(_1202_),
    .X(_0740_));
 sky130_fd_sc_hd__nor2_8 _3282_ (.A(_1114_),
    .B(_1200_),
    .Y(_1207_));
 sky130_fd_sc_hd__buf_12 _3283_ (.A(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(\rf_reg[800] ),
    .A1(_1144_),
    .S(_1208_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _3285_ (.A0(\rf_reg[801] ),
    .A1(_1147_),
    .S(_1208_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(_1065_),
    .A1(\rf_reg[108] ),
    .S(_1205_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _3287_ (.A0(\rf_reg[802] ),
    .A1(_1148_),
    .S(_1208_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(\rf_reg[803] ),
    .A1(_1149_),
    .S(_1208_),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _3289_ (.A0(\rf_reg[804] ),
    .A1(_1150_),
    .S(_1208_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\rf_reg[805] ),
    .A1(_1151_),
    .S(_1208_),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _3291_ (.A0(\rf_reg[806] ),
    .A1(_1152_),
    .S(_1208_),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(\rf_reg[807] ),
    .A1(_1153_),
    .S(_1208_),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(\rf_reg[808] ),
    .A1(_1154_),
    .S(_1208_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(\rf_reg[809] ),
    .A1(_1155_),
    .S(_1208_),
    .X(_0751_));
 sky130_fd_sc_hd__buf_16 _3295_ (.A(_1207_),
    .X(_1209_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(\rf_reg[810] ),
    .A1(_1156_),
    .S(_1209_),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(\rf_reg[811] ),
    .A1(_1158_),
    .S(_1209_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(_1066_),
    .A1(\rf_reg[109] ),
    .S(_1205_),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(\rf_reg[812] ),
    .A1(_1159_),
    .S(_1209_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(\rf_reg[813] ),
    .A1(_1160_),
    .S(_1209_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(\rf_reg[814] ),
    .A1(_1161_),
    .S(_1209_),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _3302_ (.A0(\rf_reg[815] ),
    .A1(_1162_),
    .S(_1209_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(\rf_reg[816] ),
    .A1(_1163_),
    .S(_1209_),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _3304_ (.A0(\rf_reg[817] ),
    .A1(_1164_),
    .S(_1209_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(\rf_reg[818] ),
    .A1(_1165_),
    .S(_1209_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(\rf_reg[819] ),
    .A1(_1166_),
    .S(_1209_),
    .X(_0762_));
 sky130_fd_sc_hd__buf_16 _3307_ (.A(_1207_),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_1 _3308_ (.A0(\rf_reg[820] ),
    .A1(_1167_),
    .S(_1210_),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(\rf_reg[821] ),
    .A1(_1169_),
    .S(_1210_),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _3310_ (.A0(_1067_),
    .A1(\rf_reg[110] ),
    .S(_1205_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(\rf_reg[822] ),
    .A1(_1170_),
    .S(_1210_),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _3312_ (.A0(\rf_reg[823] ),
    .A1(_1171_),
    .S(_1210_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(\rf_reg[824] ),
    .A1(_1172_),
    .S(_1210_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(\rf_reg[825] ),
    .A1(_1173_),
    .S(_1210_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(\rf_reg[826] ),
    .A1(_1174_),
    .S(_1210_),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(\rf_reg[827] ),
    .A1(_1175_),
    .S(_1210_),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(\rf_reg[828] ),
    .A1(_1176_),
    .S(_1210_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(\rf_reg[829] ),
    .A1(_1177_),
    .S(_1210_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(\rf_reg[830] ),
    .A1(_1178_),
    .S(_1207_),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _3320_ (.A0(\rf_reg[831] ),
    .A1(_1179_),
    .S(_1207_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(_1068_),
    .A1(\rf_reg[111] ),
    .S(_1205_),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _3322_ (.A0(_1058_),
    .A1(\rf_reg[39] ),
    .S(_1097_),
    .X(_0777_));
 sky130_fd_sc_hd__nor2_8 _3323_ (.A(_1119_),
    .B(_1200_),
    .Y(_1211_));
 sky130_fd_sc_hd__buf_12 _3324_ (.A(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_1 _3325_ (.A0(\rf_reg[832] ),
    .A1(_1144_),
    .S(_1212_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _3326_ (.A0(\rf_reg[833] ),
    .A1(_1147_),
    .S(_1212_),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _3327_ (.A0(\rf_reg[834] ),
    .A1(_1148_),
    .S(_1212_),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(\rf_reg[835] ),
    .A1(_1149_),
    .S(_1212_),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _3329_ (.A0(\rf_reg[836] ),
    .A1(_1150_),
    .S(_1212_),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(\rf_reg[837] ),
    .A1(_1151_),
    .S(_1212_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _3331_ (.A0(\rf_reg[838] ),
    .A1(_1152_),
    .S(_1212_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _3332_ (.A0(\rf_reg[839] ),
    .A1(_1153_),
    .S(_1212_),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _3333_ (.A0(\rf_reg[840] ),
    .A1(_1154_),
    .S(_1212_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(\rf_reg[841] ),
    .A1(_1155_),
    .S(_1212_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _3335_ (.A0(_1069_),
    .A1(\rf_reg[112] ),
    .S(_1205_),
    .X(_0788_));
 sky130_fd_sc_hd__buf_16 _3336_ (.A(_1211_),
    .X(_1213_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(\rf_reg[842] ),
    .A1(_1156_),
    .S(_1213_),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _3338_ (.A0(\rf_reg[843] ),
    .A1(_1158_),
    .S(_1213_),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(\rf_reg[844] ),
    .A1(_1159_),
    .S(_1213_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(\rf_reg[845] ),
    .A1(_1160_),
    .S(_1213_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _3341_ (.A0(\rf_reg[846] ),
    .A1(_1161_),
    .S(_1213_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _3342_ (.A0(\rf_reg[847] ),
    .A1(_1162_),
    .S(_1213_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _3343_ (.A0(\rf_reg[848] ),
    .A1(_1163_),
    .S(_1213_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(\rf_reg[849] ),
    .A1(_1164_),
    .S(_1213_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _3345_ (.A0(\rf_reg[850] ),
    .A1(_1165_),
    .S(_1213_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _3346_ (.A0(\rf_reg[851] ),
    .A1(_1166_),
    .S(_1213_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _3347_ (.A0(_1070_),
    .A1(\rf_reg[113] ),
    .S(_1205_),
    .X(_0799_));
 sky130_fd_sc_hd__buf_16 _3348_ (.A(_1211_),
    .X(_1214_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(\rf_reg[852] ),
    .A1(_1167_),
    .S(_1214_),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _3350_ (.A0(\rf_reg[853] ),
    .A1(_1169_),
    .S(_1214_),
    .X(_0801_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(\rf_reg[854] ),
    .A1(_1170_),
    .S(_1214_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _3352_ (.A0(\rf_reg[855] ),
    .A1(_1171_),
    .S(_1214_),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _3353_ (.A0(\rf_reg[856] ),
    .A1(_1172_),
    .S(_1214_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _3354_ (.A0(\rf_reg[857] ),
    .A1(_1173_),
    .S(_1214_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(\rf_reg[858] ),
    .A1(_1174_),
    .S(_1214_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _3356_ (.A0(\rf_reg[859] ),
    .A1(_1175_),
    .S(_1214_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _3357_ (.A0(\rf_reg[860] ),
    .A1(_1176_),
    .S(_1214_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(\rf_reg[861] ),
    .A1(_1177_),
    .S(_1214_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(_1071_),
    .A1(\rf_reg[114] ),
    .S(_1205_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _3360_ (.A0(\rf_reg[862] ),
    .A1(_1178_),
    .S(_1211_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _3361_ (.A0(\rf_reg[863] ),
    .A1(_1179_),
    .S(_1211_),
    .X(_0812_));
 sky130_fd_sc_hd__nor2_8 _3362_ (.A(_1100_),
    .B(_1200_),
    .Y(_1215_));
 sky130_fd_sc_hd__buf_12 _3363_ (.A(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(\rf_reg[864] ),
    .A1(_1144_),
    .S(_1216_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(\rf_reg[865] ),
    .A1(_1147_),
    .S(_1216_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(\rf_reg[866] ),
    .A1(_1148_),
    .S(_1216_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _3367_ (.A0(\rf_reg[867] ),
    .A1(_1149_),
    .S(_1216_),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(\rf_reg[868] ),
    .A1(_1150_),
    .S(_1216_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(\rf_reg[869] ),
    .A1(_1151_),
    .S(_1216_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _3370_ (.A0(\rf_reg[870] ),
    .A1(_1152_),
    .S(_1216_),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(\rf_reg[871] ),
    .A1(_1153_),
    .S(_1216_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _3372_ (.A0(_1072_),
    .A1(\rf_reg[115] ),
    .S(_1205_),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(\rf_reg[872] ),
    .A1(_1154_),
    .S(_1216_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _3374_ (.A0(\rf_reg[873] ),
    .A1(_1155_),
    .S(_1216_),
    .X(_0823_));
 sky130_fd_sc_hd__clkbuf_16 _3375_ (.A(_1215_),
    .X(_1217_));
 sky130_fd_sc_hd__mux2_1 _3376_ (.A0(\rf_reg[874] ),
    .A1(_1156_),
    .S(_1217_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(\rf_reg[875] ),
    .A1(_1158_),
    .S(_1217_),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _3378_ (.A0(\rf_reg[876] ),
    .A1(_1159_),
    .S(_1217_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(\rf_reg[877] ),
    .A1(_1160_),
    .S(_1217_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(\rf_reg[878] ),
    .A1(_1161_),
    .S(_1217_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(\rf_reg[879] ),
    .A1(_1162_),
    .S(_1217_),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(\rf_reg[880] ),
    .A1(_1163_),
    .S(_1217_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(\rf_reg[881] ),
    .A1(_1164_),
    .S(_1217_),
    .X(_0831_));
 sky130_fd_sc_hd__buf_8 _3384_ (.A(_1188_),
    .X(_1218_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(_1073_),
    .A1(\rf_reg[116] ),
    .S(_1218_),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _3386_ (.A0(\rf_reg[882] ),
    .A1(_1165_),
    .S(_1217_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _3387_ (.A0(\rf_reg[883] ),
    .A1(_1166_),
    .S(_1217_),
    .X(_0834_));
 sky130_fd_sc_hd__buf_16 _3388_ (.A(_1215_),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _3389_ (.A0(\rf_reg[884] ),
    .A1(_1167_),
    .S(_1219_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(\rf_reg[885] ),
    .A1(_1169_),
    .S(_1219_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(\rf_reg[886] ),
    .A1(_1170_),
    .S(_1219_),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(\rf_reg[887] ),
    .A1(_1171_),
    .S(_1219_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(\rf_reg[888] ),
    .A1(_1172_),
    .S(_1219_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _3394_ (.A0(\rf_reg[889] ),
    .A1(_1173_),
    .S(_1219_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(\rf_reg[890] ),
    .A1(_1174_),
    .S(_1219_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(\rf_reg[891] ),
    .A1(_1175_),
    .S(_1219_),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _3397_ (.A0(_1075_),
    .A1(\rf_reg[117] ),
    .S(_1218_),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(\rf_reg[892] ),
    .A1(_1176_),
    .S(_1219_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _3399_ (.A0(\rf_reg[893] ),
    .A1(_1177_),
    .S(_1219_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(\rf_reg[894] ),
    .A1(_1178_),
    .S(_1215_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(\rf_reg[895] ),
    .A1(_1179_),
    .S(_1215_),
    .X(_0847_));
 sky130_fd_sc_hd__nand4_4 _3402_ (.A(_0996_),
    .B(_0997_),
    .C(net5),
    .D(net46),
    .Y(_1220_));
 sky130_fd_sc_hd__nor3_4 _3403_ (.A(_0993_),
    .B(_0994_),
    .C(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__buf_12 _3404_ (.A(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(\rf_reg[896] ),
    .A1(_1144_),
    .S(_1222_),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _3406_ (.A0(\rf_reg[897] ),
    .A1(_1147_),
    .S(_1222_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _3407_ (.A0(\rf_reg[898] ),
    .A1(_1148_),
    .S(_1222_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _3408_ (.A0(\rf_reg[899] ),
    .A1(_1149_),
    .S(_1222_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(\rf_reg[900] ),
    .A1(_1150_),
    .S(_1222_),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _3410_ (.A0(\rf_reg[901] ),
    .A1(_1151_),
    .S(_1222_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(_1076_),
    .A1(\rf_reg[118] ),
    .S(_1218_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(\rf_reg[902] ),
    .A1(_1152_),
    .S(_1222_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(\rf_reg[903] ),
    .A1(_1153_),
    .S(_1222_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(\rf_reg[904] ),
    .A1(_1154_),
    .S(_1222_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(\rf_reg[905] ),
    .A1(_1155_),
    .S(_1222_),
    .X(_0858_));
 sky130_fd_sc_hd__buf_8 _3416_ (.A(_1221_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(\rf_reg[906] ),
    .A1(_1156_),
    .S(_1223_),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _3418_ (.A0(\rf_reg[907] ),
    .A1(_1158_),
    .S(_1223_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(\rf_reg[908] ),
    .A1(_1159_),
    .S(_1223_),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _3420_ (.A0(\rf_reg[909] ),
    .A1(_1160_),
    .S(_1223_),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _3421_ (.A0(\rf_reg[910] ),
    .A1(_1161_),
    .S(_1223_),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(\rf_reg[911] ),
    .A1(_1162_),
    .S(_1223_),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(_1077_),
    .A1(\rf_reg[119] ),
    .S(_1218_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(\rf_reg[912] ),
    .A1(_1163_),
    .S(_1223_),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(\rf_reg[913] ),
    .A1(_1164_),
    .S(_1223_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(\rf_reg[914] ),
    .A1(_1165_),
    .S(_1223_),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _3427_ (.A0(\rf_reg[915] ),
    .A1(_1166_),
    .S(_1223_),
    .X(_0869_));
 sky130_fd_sc_hd__buf_16 _3428_ (.A(_1221_),
    .X(_1224_));
 sky130_fd_sc_hd__mux2_1 _3429_ (.A0(\rf_reg[916] ),
    .A1(_1167_),
    .S(_1224_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(\rf_reg[917] ),
    .A1(_1169_),
    .S(_1224_),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _3431_ (.A0(\rf_reg[918] ),
    .A1(_1170_),
    .S(_1224_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(\rf_reg[919] ),
    .A1(_1171_),
    .S(_1224_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(\rf_reg[920] ),
    .A1(_1172_),
    .S(_1224_),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(\rf_reg[921] ),
    .A1(_1173_),
    .S(_1224_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(_1078_),
    .A1(\rf_reg[120] ),
    .S(_1218_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(\rf_reg[922] ),
    .A1(_1174_),
    .S(_1224_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _3437_ (.A0(\rf_reg[923] ),
    .A1(_1175_),
    .S(_1224_),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(\rf_reg[924] ),
    .A1(_1176_),
    .S(_1224_),
    .X(_0879_));
 sky130_fd_sc_hd__mux2_1 _3439_ (.A0(\rf_reg[925] ),
    .A1(_1177_),
    .S(_1224_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(\rf_reg[926] ),
    .A1(_1178_),
    .S(_1221_),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(\rf_reg[927] ),
    .A1(_1179_),
    .S(_1221_),
    .X(_0882_));
 sky130_fd_sc_hd__nor2_8 _3442_ (.A(_1114_),
    .B(_1220_),
    .Y(_1225_));
 sky130_fd_sc_hd__buf_12 _3443_ (.A(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(\rf_reg[928] ),
    .A1(_1144_),
    .S(_1226_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(\rf_reg[929] ),
    .A1(_1147_),
    .S(_1226_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(\rf_reg[930] ),
    .A1(_1148_),
    .S(_1226_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(\rf_reg[931] ),
    .A1(_1149_),
    .S(_1226_),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(_1079_),
    .A1(\rf_reg[121] ),
    .S(_1218_),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(_1060_),
    .A1(\rf_reg[40] ),
    .S(_1000_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(\rf_reg[932] ),
    .A1(_1150_),
    .S(_1226_),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(\rf_reg[933] ),
    .A1(_1151_),
    .S(_1226_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(\rf_reg[934] ),
    .A1(_1152_),
    .S(_1226_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(\rf_reg[935] ),
    .A1(_1153_),
    .S(_1226_),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _3454_ (.A0(\rf_reg[936] ),
    .A1(_1154_),
    .S(_1226_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(\rf_reg[937] ),
    .A1(_1155_),
    .S(_1226_),
    .X(_0894_));
 sky130_fd_sc_hd__buf_16 _3456_ (.A(_1225_),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(\rf_reg[938] ),
    .A1(_1156_),
    .S(_1227_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(\rf_reg[939] ),
    .A1(_1158_),
    .S(_1227_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _3459_ (.A0(\rf_reg[940] ),
    .A1(_1159_),
    .S(_1227_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(\rf_reg[941] ),
    .A1(_1160_),
    .S(_1227_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(_1080_),
    .A1(\rf_reg[122] ),
    .S(_1218_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(\rf_reg[942] ),
    .A1(_1161_),
    .S(_1227_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _3463_ (.A0(\rf_reg[943] ),
    .A1(_1162_),
    .S(_1227_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(\rf_reg[944] ),
    .A1(_1163_),
    .S(_1227_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _3465_ (.A0(\rf_reg[945] ),
    .A1(_1164_),
    .S(_1227_),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _3466_ (.A0(\rf_reg[946] ),
    .A1(_1165_),
    .S(_1227_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _3467_ (.A0(\rf_reg[947] ),
    .A1(_1166_),
    .S(_1227_),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_16 _3468_ (.A(_1225_),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(\rf_reg[948] ),
    .A1(_1167_),
    .S(_1228_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(\rf_reg[949] ),
    .A1(_1169_),
    .S(_1228_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _3471_ (.A0(\rf_reg[950] ),
    .A1(_1170_),
    .S(_1228_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _3472_ (.A0(\rf_reg[951] ),
    .A1(_1171_),
    .S(_1228_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(_1081_),
    .A1(\rf_reg[123] ),
    .S(_1218_),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(\rf_reg[952] ),
    .A1(_1172_),
    .S(_1228_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _3475_ (.A0(\rf_reg[953] ),
    .A1(_1173_),
    .S(_1228_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(\rf_reg[954] ),
    .A1(_1174_),
    .S(_1228_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _3477_ (.A0(\rf_reg[955] ),
    .A1(_1175_),
    .S(_1228_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(\rf_reg[956] ),
    .A1(_1176_),
    .S(_1228_),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _3479_ (.A0(\rf_reg[957] ),
    .A1(_1177_),
    .S(_1228_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(\rf_reg[958] ),
    .A1(_1178_),
    .S(_1225_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _3481_ (.A0(\rf_reg[959] ),
    .A1(_1179_),
    .S(_1225_),
    .X(_0918_));
 sky130_fd_sc_hd__nor2_8 _3482_ (.A(_1119_),
    .B(_1220_),
    .Y(_1229_));
 sky130_fd_sc_hd__buf_16 _3483_ (.A(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _3484_ (.A0(\rf_reg[960] ),
    .A1(_1144_),
    .S(_1230_),
    .X(_0919_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(\rf_reg[961] ),
    .A1(_1147_),
    .S(_1230_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(_1082_),
    .A1(\rf_reg[124] ),
    .S(_1218_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _3487_ (.A0(\rf_reg[962] ),
    .A1(_1148_),
    .S(_1230_),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(\rf_reg[963] ),
    .A1(_1149_),
    .S(_1230_),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(\rf_reg[964] ),
    .A1(_1150_),
    .S(_1230_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(\rf_reg[965] ),
    .A1(_1151_),
    .S(_1230_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _3491_ (.A0(\rf_reg[966] ),
    .A1(_1152_),
    .S(_1230_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(\rf_reg[967] ),
    .A1(_1153_),
    .S(_1230_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(\rf_reg[968] ),
    .A1(_1154_),
    .S(_1230_),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(\rf_reg[969] ),
    .A1(_1155_),
    .S(_1230_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_16 _3495_ (.A(_1229_),
    .X(_1231_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(\rf_reg[970] ),
    .A1(_1156_),
    .S(_1231_),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_1 _3497_ (.A0(\rf_reg[971] ),
    .A1(_1158_),
    .S(_1231_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(_1083_),
    .A1(\rf_reg[125] ),
    .S(_1218_),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _3499_ (.A0(\rf_reg[972] ),
    .A1(_1159_),
    .S(_1231_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(\rf_reg[973] ),
    .A1(_1160_),
    .S(_1231_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _3501_ (.A0(\rf_reg[974] ),
    .A1(_1161_),
    .S(_1231_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _3502_ (.A0(\rf_reg[975] ),
    .A1(_1162_),
    .S(_1231_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _3503_ (.A0(\rf_reg[976] ),
    .A1(_1163_),
    .S(_1231_),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(\rf_reg[977] ),
    .A1(_1164_),
    .S(_1231_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(\rf_reg[978] ),
    .A1(_1165_),
    .S(_1231_),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(\rf_reg[979] ),
    .A1(_1166_),
    .S(_1231_),
    .X(_0940_));
 sky130_fd_sc_hd__clkbuf_16 _3507_ (.A(_1229_),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _3508_ (.A0(\rf_reg[980] ),
    .A1(_1167_),
    .S(_1232_),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_1 _3509_ (.A0(\rf_reg[981] ),
    .A1(_1169_),
    .S(_1232_),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _3510_ (.A0(_1084_),
    .A1(\rf_reg[126] ),
    .S(_1188_),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(\rf_reg[982] ),
    .A1(_1170_),
    .S(_1232_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(\rf_reg[983] ),
    .A1(_1171_),
    .S(_1232_),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _3513_ (.A0(\rf_reg[984] ),
    .A1(_1172_),
    .S(_1232_),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(\rf_reg[985] ),
    .A1(_1173_),
    .S(_1232_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(\rf_reg[986] ),
    .A1(_1174_),
    .S(_1232_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(\rf_reg[987] ),
    .A1(_1175_),
    .S(_1232_),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _3517_ (.A0(\rf_reg[988] ),
    .A1(_1176_),
    .S(_1232_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(\rf_reg[989] ),
    .A1(_1177_),
    .S(_1232_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(\rf_reg[990] ),
    .A1(_1178_),
    .S(_1229_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(\rf_reg[991] ),
    .A1(_1179_),
    .S(_1229_),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _3521_ (.A0(_1085_),
    .A1(\rf_reg[127] ),
    .S(_1188_),
    .X(_0954_));
 sky130_fd_sc_hd__nor2_8 _3522_ (.A(_1100_),
    .B(_1220_),
    .Y(_1233_));
 sky130_fd_sc_hd__buf_12 _3523_ (.A(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _3524_ (.A0(\rf_reg[992] ),
    .A1(net6),
    .S(_1234_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(\rf_reg[993] ),
    .A1(net25),
    .S(_1234_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _3526_ (.A0(\rf_reg[994] ),
    .A1(net36),
    .S(_1234_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3527_ (.A0(\rf_reg[995] ),
    .A1(net39),
    .S(_1234_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(\rf_reg[996] ),
    .A1(net40),
    .S(_1234_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _3529_ (.A0(\rf_reg[997] ),
    .A1(net41),
    .S(_1234_),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(\rf_reg[998] ),
    .A1(net42),
    .S(_1234_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _3531_ (.A0(\rf_reg[999] ),
    .A1(net43),
    .S(_1234_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(\rf_reg[1000] ),
    .A1(net44),
    .S(_1234_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _3533_ (.A0(\rf_reg[1001] ),
    .A1(net45),
    .S(_1234_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(_1048_),
    .A1(\rf_reg[128] ),
    .S(_1028_),
    .X(_0965_));
 sky130_fd_sc_hd__buf_16 _3535_ (.A(_1233_),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _3536_ (.A0(\rf_reg[1002] ),
    .A1(net7),
    .S(_1235_),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _3537_ (.A0(\rf_reg[1003] ),
    .A1(net16),
    .S(_1235_),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(\rf_reg[1004] ),
    .A1(net17),
    .S(_1235_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(\rf_reg[1005] ),
    .A1(net18),
    .S(_1235_),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _3540_ (.A0(\rf_reg[1006] ),
    .A1(net19),
    .S(_1235_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(\rf_reg[1007] ),
    .A1(net20),
    .S(_1235_),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(\rf_reg[1008] ),
    .A1(net21),
    .S(_1235_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(\rf_reg[1009] ),
    .A1(net22),
    .S(_1235_),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(\rf_reg[1010] ),
    .A1(net23),
    .S(_1235_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(\rf_reg[1011] ),
    .A1(net24),
    .S(_1235_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(_1052_),
    .A1(\rf_reg[129] ),
    .S(_1028_),
    .X(_0976_));
 sky130_fd_sc_hd__buf_16 _3547_ (.A(_1233_),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(\rf_reg[1012] ),
    .A1(net26),
    .S(_1236_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(\rf_reg[1013] ),
    .A1(net27),
    .S(_1236_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(\rf_reg[1014] ),
    .A1(net28),
    .S(_1236_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(\rf_reg[1015] ),
    .A1(net29),
    .S(_1236_),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(\rf_reg[1016] ),
    .A1(net30),
    .S(_1236_),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _3553_ (.A0(\rf_reg[1017] ),
    .A1(net31),
    .S(_1236_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _3554_ (.A0(\rf_reg[1018] ),
    .A1(net32),
    .S(_1236_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(\rf_reg[1019] ),
    .A1(net33),
    .S(_1236_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(\rf_reg[1020] ),
    .A1(net34),
    .S(_1236_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(\rf_reg[1021] ),
    .A1(net35),
    .S(_1236_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(_1053_),
    .A1(\rf_reg[130] ),
    .S(_1005_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(\rf_reg[1022] ),
    .A1(net37),
    .S(_1233_),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(\rf_reg[1023] ),
    .A1(net38),
    .S(_1233_),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(_1054_),
    .A1(\rf_reg[131] ),
    .S(_1005_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _3562_ (.A0(_1061_),
    .A1(\rf_reg[41] ),
    .S(_1000_),
    .X(_0991_));
 sky130_fd_sc_hd__buf_2 _3563_ (.A(raddr_a_i[0]),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_4 _3564_ (.A(raddr_a_i[1]),
    .X(_1238_));
 sky130_fd_sc_hd__nor2b_1 _3565_ (.A(_1237_),
    .B_N(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__buf_4 _3566_ (.A(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__buf_6 _3567_ (.A(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__buf_16 _3568_ (.A(_1238_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _3569_ (.A0(\rf_reg[32] ),
    .A1(\rf_reg[96] ),
    .S(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__buf_8 _3570_ (.A(_1237_),
    .X(_1244_));
 sky130_fd_sc_hd__buf_8 _3571_ (.A(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__buf_6 _3572_ (.A(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__a22o_1 _3573_ (.A1(\rf_reg[64] ),
    .A2(_1241_),
    .B1(_1243_),
    .B2(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__buf_16 _3574_ (.A(_1237_),
    .X(_1248_));
 sky130_fd_sc_hd__buf_16 _3575_ (.A(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__buf_8 _3576_ (.A(_1242_),
    .X(_1250_));
 sky130_fd_sc_hd__mux4_1 _3577_ (.A0(\rf_reg[128] ),
    .A1(\rf_reg[160] ),
    .A2(\rf_reg[192] ),
    .A3(\rf_reg[224] ),
    .S0(_1249_),
    .S1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__buf_16 _3578_ (.A(_1248_),
    .X(_1252_));
 sky130_fd_sc_hd__buf_6 _3579_ (.A(_1238_),
    .X(_1253_));
 sky130_fd_sc_hd__buf_16 _3580_ (.A(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__buf_16 _3581_ (.A(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__mux4_1 _3582_ (.A0(\rf_reg[512] ),
    .A1(\rf_reg[544] ),
    .A2(\rf_reg[576] ),
    .A3(\rf_reg[608] ),
    .S0(_1252_),
    .S1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__buf_12 _3583_ (.A(_1237_),
    .X(_1257_));
 sky130_fd_sc_hd__buf_16 _3584_ (.A(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__buf_8 _3585_ (.A(_1253_),
    .X(_1259_));
 sky130_fd_sc_hd__buf_8 _3586_ (.A(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__mux4_1 _3587_ (.A0(\rf_reg[640] ),
    .A1(\rf_reg[672] ),
    .A2(\rf_reg[704] ),
    .A3(\rf_reg[736] ),
    .S0(_1258_),
    .S1(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__buf_12 _3588_ (.A(raddr_a_i[2]),
    .X(_1262_));
 sky130_fd_sc_hd__buf_8 _3589_ (.A(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__buf_12 _3590_ (.A(raddr_a_i[4]),
    .X(_1264_));
 sky130_fd_sc_hd__buf_8 _3591_ (.A(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__mux4_1 _3592_ (.A0(_1247_),
    .A1(_1251_),
    .A2(_1256_),
    .A3(_1261_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__buf_12 _3593_ (.A(_1257_),
    .X(_1267_));
 sky130_fd_sc_hd__buf_12 _3594_ (.A(_1254_),
    .X(_1268_));
 sky130_fd_sc_hd__mux4_1 _3595_ (.A0(\rf_reg[256] ),
    .A1(\rf_reg[288] ),
    .A2(\rf_reg[320] ),
    .A3(\rf_reg[352] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__buf_12 _3596_ (.A(_1248_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_16 _3597_ (.A(_1242_),
    .X(_1271_));
 sky130_fd_sc_hd__mux4_1 _3598_ (.A0(\rf_reg[384] ),
    .A1(\rf_reg[416] ),
    .A2(\rf_reg[448] ),
    .A3(\rf_reg[480] ),
    .S0(_1270_),
    .S1(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_16 _3599_ (.A(_1257_),
    .X(_1273_));
 sky130_fd_sc_hd__buf_6 _3600_ (.A(_1254_),
    .X(_1274_));
 sky130_fd_sc_hd__mux4_1 _3601_ (.A0(\rf_reg[768] ),
    .A1(\rf_reg[800] ),
    .A2(\rf_reg[832] ),
    .A3(\rf_reg[864] ),
    .S0(_1273_),
    .S1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__buf_8 _3602_ (.A(_1259_),
    .X(_1276_));
 sky130_fd_sc_hd__mux4_1 _3603_ (.A0(\rf_reg[896] ),
    .A1(\rf_reg[928] ),
    .A2(\rf_reg[960] ),
    .A3(\rf_reg[992] ),
    .S0(_1245_),
    .S1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_16 _3604_ (.A(_1262_),
    .X(_1278_));
 sky130_fd_sc_hd__buf_16 _3605_ (.A(_1264_),
    .X(_1279_));
 sky130_fd_sc_hd__mux4_1 _3606_ (.A0(_1269_),
    .A1(_1272_),
    .A2(_1275_),
    .A3(_1277_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__buf_6 _3607_ (.A(raddr_a_i[3]),
    .X(_1281_));
 sky130_fd_sc_hd__buf_8 _3608_ (.A(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_2 _3609_ (.A0(_1266_),
    .A1(_1280_),
    .S(_1282_),
    .X(net47));
 sky130_fd_sc_hd__mux2_1 _3610_ (.A0(\rf_reg[42] ),
    .A1(\rf_reg[106] ),
    .S(_1242_),
    .X(_1283_));
 sky130_fd_sc_hd__a22o_1 _3611_ (.A1(\rf_reg[74] ),
    .A2(_1241_),
    .B1(_1283_),
    .B2(_1246_),
    .X(_1284_));
 sky130_fd_sc_hd__mux4_1 _3612_ (.A0(\rf_reg[138] ),
    .A1(\rf_reg[170] ),
    .A2(\rf_reg[202] ),
    .A3(\rf_reg[234] ),
    .S0(_1249_),
    .S1(_1250_),
    .X(_1285_));
 sky130_fd_sc_hd__mux4_1 _3613_ (.A0(\rf_reg[522] ),
    .A1(\rf_reg[554] ),
    .A2(\rf_reg[586] ),
    .A3(\rf_reg[618] ),
    .S0(_1252_),
    .S1(_1255_),
    .X(_1286_));
 sky130_fd_sc_hd__mux4_1 _3614_ (.A0(\rf_reg[650] ),
    .A1(\rf_reg[682] ),
    .A2(\rf_reg[714] ),
    .A3(\rf_reg[746] ),
    .S0(_1258_),
    .S1(_1260_),
    .X(_1287_));
 sky130_fd_sc_hd__mux4_1 _3615_ (.A0(_1284_),
    .A1(_1285_),
    .A2(_1286_),
    .A3(_1287_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1288_));
 sky130_fd_sc_hd__buf_16 _3616_ (.A(_1257_),
    .X(_1289_));
 sky130_fd_sc_hd__mux4_1 _3617_ (.A0(\rf_reg[266] ),
    .A1(\rf_reg[298] ),
    .A2(\rf_reg[330] ),
    .A3(\rf_reg[362] ),
    .S0(_1289_),
    .S1(_1268_),
    .X(_1290_));
 sky130_fd_sc_hd__mux4_1 _3618_ (.A0(\rf_reg[394] ),
    .A1(\rf_reg[426] ),
    .A2(\rf_reg[458] ),
    .A3(\rf_reg[490] ),
    .S0(_1270_),
    .S1(_1271_),
    .X(_1291_));
 sky130_fd_sc_hd__mux4_1 _3619_ (.A0(\rf_reg[778] ),
    .A1(\rf_reg[810] ),
    .A2(\rf_reg[842] ),
    .A3(\rf_reg[874] ),
    .S0(_1273_),
    .S1(_1274_),
    .X(_1292_));
 sky130_fd_sc_hd__mux4_1 _3620_ (.A0(\rf_reg[906] ),
    .A1(\rf_reg[938] ),
    .A2(\rf_reg[970] ),
    .A3(\rf_reg[1002] ),
    .S0(_1245_),
    .S1(_1276_),
    .X(_1293_));
 sky130_fd_sc_hd__mux4_1 _3621_ (.A0(_1290_),
    .A1(_1291_),
    .A2(_1292_),
    .A3(_1293_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_2 _3622_ (.A0(_1288_),
    .A1(_1294_),
    .S(_1282_),
    .X(net48));
 sky130_fd_sc_hd__mux2_1 _3623_ (.A0(\rf_reg[43] ),
    .A1(\rf_reg[107] ),
    .S(_1242_),
    .X(_1295_));
 sky130_fd_sc_hd__a22o_1 _3624_ (.A1(\rf_reg[75] ),
    .A2(_1241_),
    .B1(_1295_),
    .B2(_1246_),
    .X(_1296_));
 sky130_fd_sc_hd__mux4_1 _3625_ (.A0(\rf_reg[139] ),
    .A1(\rf_reg[171] ),
    .A2(\rf_reg[203] ),
    .A3(\rf_reg[235] ),
    .S0(_1249_),
    .S1(_1250_),
    .X(_1297_));
 sky130_fd_sc_hd__buf_8 _3626_ (.A(_1254_),
    .X(_1298_));
 sky130_fd_sc_hd__mux4_1 _3627_ (.A0(\rf_reg[523] ),
    .A1(\rf_reg[555] ),
    .A2(\rf_reg[587] ),
    .A3(\rf_reg[619] ),
    .S0(_1252_),
    .S1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__mux4_1 _3628_ (.A0(\rf_reg[651] ),
    .A1(\rf_reg[683] ),
    .A2(\rf_reg[715] ),
    .A3(\rf_reg[747] ),
    .S0(_1258_),
    .S1(_1260_),
    .X(_1300_));
 sky130_fd_sc_hd__mux4_1 _3629_ (.A0(_1296_),
    .A1(_1297_),
    .A2(_1299_),
    .A3(_1300_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1301_));
 sky130_fd_sc_hd__mux4_1 _3630_ (.A0(\rf_reg[267] ),
    .A1(\rf_reg[299] ),
    .A2(\rf_reg[331] ),
    .A3(\rf_reg[363] ),
    .S0(_1289_),
    .S1(_1268_),
    .X(_1302_));
 sky130_fd_sc_hd__mux4_1 _3631_ (.A0(\rf_reg[395] ),
    .A1(\rf_reg[427] ),
    .A2(\rf_reg[459] ),
    .A3(\rf_reg[491] ),
    .S0(_1270_),
    .S1(_1271_),
    .X(_1303_));
 sky130_fd_sc_hd__mux4_1 _3632_ (.A0(\rf_reg[779] ),
    .A1(\rf_reg[811] ),
    .A2(\rf_reg[843] ),
    .A3(\rf_reg[875] ),
    .S0(_1273_),
    .S1(_1274_),
    .X(_1304_));
 sky130_fd_sc_hd__mux4_1 _3633_ (.A0(\rf_reg[907] ),
    .A1(\rf_reg[939] ),
    .A2(\rf_reg[971] ),
    .A3(\rf_reg[1003] ),
    .S0(_1245_),
    .S1(_1276_),
    .X(_1305_));
 sky130_fd_sc_hd__mux4_1 _3634_ (.A0(_1302_),
    .A1(_1303_),
    .A2(_1304_),
    .A3(_1305_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1306_));
 sky130_fd_sc_hd__mux2_2 _3635_ (.A0(_1301_),
    .A1(_1306_),
    .S(_1282_),
    .X(net49));
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(\rf_reg[44] ),
    .A1(\rf_reg[108] ),
    .S(_1242_),
    .X(_1307_));
 sky130_fd_sc_hd__a22o_1 _3637_ (.A1(\rf_reg[76] ),
    .A2(_1241_),
    .B1(_1307_),
    .B2(_1246_),
    .X(_1308_));
 sky130_fd_sc_hd__buf_8 _3638_ (.A(_1248_),
    .X(_1309_));
 sky130_fd_sc_hd__mux4_1 _3639_ (.A0(\rf_reg[140] ),
    .A1(\rf_reg[172] ),
    .A2(\rf_reg[204] ),
    .A3(\rf_reg[236] ),
    .S0(_1309_),
    .S1(_1250_),
    .X(_1310_));
 sky130_fd_sc_hd__mux4_1 _3640_ (.A0(\rf_reg[524] ),
    .A1(\rf_reg[556] ),
    .A2(\rf_reg[588] ),
    .A3(\rf_reg[620] ),
    .S0(_1252_),
    .S1(_1298_),
    .X(_1311_));
 sky130_fd_sc_hd__buf_8 _3641_ (.A(_1257_),
    .X(_1312_));
 sky130_fd_sc_hd__mux4_1 _3642_ (.A0(\rf_reg[652] ),
    .A1(\rf_reg[684] ),
    .A2(\rf_reg[716] ),
    .A3(\rf_reg[748] ),
    .S0(_1312_),
    .S1(_1260_),
    .X(_1313_));
 sky130_fd_sc_hd__mux4_1 _3643_ (.A0(_1308_),
    .A1(_1310_),
    .A2(_1311_),
    .A3(_1313_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1314_));
 sky130_fd_sc_hd__mux4_1 _3644_ (.A0(\rf_reg[268] ),
    .A1(\rf_reg[300] ),
    .A2(\rf_reg[332] ),
    .A3(\rf_reg[364] ),
    .S0(_1289_),
    .S1(_1268_),
    .X(_1315_));
 sky130_fd_sc_hd__mux4_1 _3645_ (.A0(\rf_reg[396] ),
    .A1(\rf_reg[428] ),
    .A2(\rf_reg[460] ),
    .A3(\rf_reg[492] ),
    .S0(_1270_),
    .S1(_1271_),
    .X(_1316_));
 sky130_fd_sc_hd__mux4_1 _3646_ (.A0(\rf_reg[780] ),
    .A1(\rf_reg[812] ),
    .A2(\rf_reg[844] ),
    .A3(\rf_reg[876] ),
    .S0(_1273_),
    .S1(_1274_),
    .X(_1317_));
 sky130_fd_sc_hd__mux4_1 _3647_ (.A0(\rf_reg[908] ),
    .A1(\rf_reg[940] ),
    .A2(\rf_reg[972] ),
    .A3(\rf_reg[1004] ),
    .S0(_1245_),
    .S1(_1276_),
    .X(_1318_));
 sky130_fd_sc_hd__mux4_1 _3648_ (.A0(_1315_),
    .A1(_1316_),
    .A2(_1317_),
    .A3(_1318_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(_1314_),
    .A1(_1319_),
    .S(_1282_),
    .X(net50));
 sky130_fd_sc_hd__buf_8 _3650_ (.A(_1238_),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_1 _3651_ (.A0(\rf_reg[45] ),
    .A1(\rf_reg[109] ),
    .S(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__a22o_1 _3652_ (.A1(\rf_reg[77] ),
    .A2(_1241_),
    .B1(_1321_),
    .B2(_1246_),
    .X(_1322_));
 sky130_fd_sc_hd__mux4_1 _3653_ (.A0(\rf_reg[141] ),
    .A1(\rf_reg[173] ),
    .A2(\rf_reg[205] ),
    .A3(\rf_reg[237] ),
    .S0(_1309_),
    .S1(_1250_),
    .X(_1323_));
 sky130_fd_sc_hd__mux4_1 _3654_ (.A0(\rf_reg[525] ),
    .A1(\rf_reg[557] ),
    .A2(\rf_reg[589] ),
    .A3(\rf_reg[621] ),
    .S0(_1252_),
    .S1(_1298_),
    .X(_1324_));
 sky130_fd_sc_hd__mux4_1 _3655_ (.A0(\rf_reg[653] ),
    .A1(\rf_reg[685] ),
    .A2(\rf_reg[717] ),
    .A3(\rf_reg[749] ),
    .S0(_1312_),
    .S1(_1260_),
    .X(_1325_));
 sky130_fd_sc_hd__mux4_1 _3656_ (.A0(_1322_),
    .A1(_1323_),
    .A2(_1324_),
    .A3(_1325_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1326_));
 sky130_fd_sc_hd__mux4_1 _3657_ (.A0(\rf_reg[269] ),
    .A1(\rf_reg[301] ),
    .A2(\rf_reg[333] ),
    .A3(\rf_reg[365] ),
    .S0(_1289_),
    .S1(_1268_),
    .X(_1327_));
 sky130_fd_sc_hd__mux4_1 _3658_ (.A0(\rf_reg[397] ),
    .A1(\rf_reg[429] ),
    .A2(\rf_reg[461] ),
    .A3(\rf_reg[493] ),
    .S0(_1270_),
    .S1(_1271_),
    .X(_1328_));
 sky130_fd_sc_hd__buf_8 _3659_ (.A(_1254_),
    .X(_1329_));
 sky130_fd_sc_hd__mux4_1 _3660_ (.A0(\rf_reg[781] ),
    .A1(\rf_reg[813] ),
    .A2(\rf_reg[845] ),
    .A3(\rf_reg[877] ),
    .S0(_1273_),
    .S1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__mux4_1 _3661_ (.A0(\rf_reg[909] ),
    .A1(\rf_reg[941] ),
    .A2(\rf_reg[973] ),
    .A3(\rf_reg[1005] ),
    .S0(_1245_),
    .S1(_1276_),
    .X(_1331_));
 sky130_fd_sc_hd__mux4_1 _3662_ (.A0(_1327_),
    .A1(_1328_),
    .A2(_1330_),
    .A3(_1331_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1332_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(_1326_),
    .A1(_1332_),
    .S(_1282_),
    .X(net51));
 sky130_fd_sc_hd__mux2_1 _3664_ (.A0(\rf_reg[46] ),
    .A1(\rf_reg[110] ),
    .S(_1320_),
    .X(_1333_));
 sky130_fd_sc_hd__a22o_1 _3665_ (.A1(\rf_reg[78] ),
    .A2(_1241_),
    .B1(_1333_),
    .B2(_1246_),
    .X(_1334_));
 sky130_fd_sc_hd__mux4_1 _3666_ (.A0(\rf_reg[142] ),
    .A1(\rf_reg[174] ),
    .A2(\rf_reg[206] ),
    .A3(\rf_reg[238] ),
    .S0(_1309_),
    .S1(_1250_),
    .X(_1335_));
 sky130_fd_sc_hd__mux4_1 _3667_ (.A0(\rf_reg[526] ),
    .A1(\rf_reg[558] ),
    .A2(\rf_reg[590] ),
    .A3(\rf_reg[622] ),
    .S0(_1252_),
    .S1(_1298_),
    .X(_1336_));
 sky130_fd_sc_hd__mux4_1 _3668_ (.A0(\rf_reg[654] ),
    .A1(\rf_reg[686] ),
    .A2(\rf_reg[718] ),
    .A3(\rf_reg[750] ),
    .S0(_1312_),
    .S1(_1260_),
    .X(_1337_));
 sky130_fd_sc_hd__mux4_1 _3669_ (.A0(_1334_),
    .A1(_1335_),
    .A2(_1336_),
    .A3(_1337_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1338_));
 sky130_fd_sc_hd__mux4_1 _3670_ (.A0(\rf_reg[270] ),
    .A1(\rf_reg[302] ),
    .A2(\rf_reg[334] ),
    .A3(\rf_reg[366] ),
    .S0(_1289_),
    .S1(_1268_),
    .X(_1339_));
 sky130_fd_sc_hd__buf_16 _3671_ (.A(_1248_),
    .X(_1340_));
 sky130_fd_sc_hd__mux4_1 _3672_ (.A0(\rf_reg[398] ),
    .A1(\rf_reg[430] ),
    .A2(\rf_reg[462] ),
    .A3(\rf_reg[494] ),
    .S0(_1340_),
    .S1(_1271_),
    .X(_1341_));
 sky130_fd_sc_hd__mux4_1 _3673_ (.A0(\rf_reg[782] ),
    .A1(\rf_reg[814] ),
    .A2(\rf_reg[846] ),
    .A3(\rf_reg[878] ),
    .S0(_1273_),
    .S1(_1329_),
    .X(_1342_));
 sky130_fd_sc_hd__buf_16 _3674_ (.A(_1257_),
    .X(_1343_));
 sky130_fd_sc_hd__mux4_1 _3675_ (.A0(\rf_reg[910] ),
    .A1(\rf_reg[942] ),
    .A2(\rf_reg[974] ),
    .A3(\rf_reg[1006] ),
    .S0(_1343_),
    .S1(_1276_),
    .X(_1344_));
 sky130_fd_sc_hd__mux4_1 _3676_ (.A0(_1339_),
    .A1(_1341_),
    .A2(_1342_),
    .A3(_1344_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1345_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(_1338_),
    .A1(_1345_),
    .S(_1282_),
    .X(net52));
 sky130_fd_sc_hd__mux2_1 _3678_ (.A0(\rf_reg[47] ),
    .A1(\rf_reg[111] ),
    .S(_1320_),
    .X(_1346_));
 sky130_fd_sc_hd__a22o_1 _3679_ (.A1(\rf_reg[79] ),
    .A2(_1241_),
    .B1(_1346_),
    .B2(_1246_),
    .X(_1347_));
 sky130_fd_sc_hd__mux4_1 _3680_ (.A0(\rf_reg[143] ),
    .A1(\rf_reg[175] ),
    .A2(\rf_reg[207] ),
    .A3(\rf_reg[239] ),
    .S0(_1309_),
    .S1(_1250_),
    .X(_1348_));
 sky130_fd_sc_hd__mux4_1 _3681_ (.A0(\rf_reg[527] ),
    .A1(\rf_reg[559] ),
    .A2(\rf_reg[591] ),
    .A3(\rf_reg[623] ),
    .S0(_1252_),
    .S1(_1298_),
    .X(_1349_));
 sky130_fd_sc_hd__mux4_1 _3682_ (.A0(\rf_reg[655] ),
    .A1(\rf_reg[687] ),
    .A2(\rf_reg[719] ),
    .A3(\rf_reg[751] ),
    .S0(_1312_),
    .S1(_1260_),
    .X(_1350_));
 sky130_fd_sc_hd__mux4_1 _3683_ (.A0(_1347_),
    .A1(_1348_),
    .A2(_1349_),
    .A3(_1350_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1351_));
 sky130_fd_sc_hd__buf_8 _3684_ (.A(_1254_),
    .X(_1352_));
 sky130_fd_sc_hd__mux4_1 _3685_ (.A0(\rf_reg[271] ),
    .A1(\rf_reg[303] ),
    .A2(\rf_reg[335] ),
    .A3(\rf_reg[367] ),
    .S0(_1289_),
    .S1(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__mux4_1 _3686_ (.A0(\rf_reg[399] ),
    .A1(\rf_reg[431] ),
    .A2(\rf_reg[463] ),
    .A3(\rf_reg[495] ),
    .S0(_1340_),
    .S1(_1271_),
    .X(_1354_));
 sky130_fd_sc_hd__mux4_1 _3687_ (.A0(\rf_reg[783] ),
    .A1(\rf_reg[815] ),
    .A2(\rf_reg[847] ),
    .A3(\rf_reg[879] ),
    .S0(_1273_),
    .S1(_1329_),
    .X(_1355_));
 sky130_fd_sc_hd__mux4_1 _3688_ (.A0(\rf_reg[911] ),
    .A1(\rf_reg[943] ),
    .A2(\rf_reg[975] ),
    .A3(\rf_reg[1007] ),
    .S0(_1343_),
    .S1(_1276_),
    .X(_1356_));
 sky130_fd_sc_hd__mux4_1 _3689_ (.A0(_1353_),
    .A1(_1354_),
    .A2(_1355_),
    .A3(_1356_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1357_));
 sky130_fd_sc_hd__mux2_1 _3690_ (.A0(_1351_),
    .A1(_1357_),
    .S(_1282_),
    .X(net53));
 sky130_fd_sc_hd__mux2_1 _3691_ (.A0(\rf_reg[48] ),
    .A1(\rf_reg[112] ),
    .S(_1320_),
    .X(_1358_));
 sky130_fd_sc_hd__a22o_1 _3692_ (.A1(\rf_reg[80] ),
    .A2(_1241_),
    .B1(_1358_),
    .B2(_1246_),
    .X(_1359_));
 sky130_fd_sc_hd__mux4_1 _3693_ (.A0(\rf_reg[144] ),
    .A1(\rf_reg[176] ),
    .A2(\rf_reg[208] ),
    .A3(\rf_reg[240] ),
    .S0(_1309_),
    .S1(_1250_),
    .X(_1360_));
 sky130_fd_sc_hd__buf_8 _3694_ (.A(_1248_),
    .X(_1361_));
 sky130_fd_sc_hd__mux4_1 _3695_ (.A0(\rf_reg[528] ),
    .A1(\rf_reg[560] ),
    .A2(\rf_reg[592] ),
    .A3(\rf_reg[624] ),
    .S0(_1361_),
    .S1(_1298_),
    .X(_1362_));
 sky130_fd_sc_hd__mux4_1 _3696_ (.A0(\rf_reg[656] ),
    .A1(\rf_reg[688] ),
    .A2(\rf_reg[720] ),
    .A3(\rf_reg[752] ),
    .S0(_1312_),
    .S1(_1260_),
    .X(_1363_));
 sky130_fd_sc_hd__mux4_1 _3697_ (.A0(_1359_),
    .A1(_1360_),
    .A2(_1362_),
    .A3(_1363_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1364_));
 sky130_fd_sc_hd__mux4_1 _3698_ (.A0(\rf_reg[272] ),
    .A1(\rf_reg[304] ),
    .A2(\rf_reg[336] ),
    .A3(\rf_reg[368] ),
    .S0(_1289_),
    .S1(_1352_),
    .X(_1365_));
 sky130_fd_sc_hd__mux4_1 _3699_ (.A0(\rf_reg[400] ),
    .A1(\rf_reg[432] ),
    .A2(\rf_reg[464] ),
    .A3(\rf_reg[496] ),
    .S0(_1340_),
    .S1(_1271_),
    .X(_1366_));
 sky130_fd_sc_hd__mux4_1 _3700_ (.A0(\rf_reg[784] ),
    .A1(\rf_reg[816] ),
    .A2(\rf_reg[848] ),
    .A3(\rf_reg[880] ),
    .S0(_1273_),
    .S1(_1329_),
    .X(_1367_));
 sky130_fd_sc_hd__mux4_1 _3701_ (.A0(\rf_reg[912] ),
    .A1(\rf_reg[944] ),
    .A2(\rf_reg[976] ),
    .A3(\rf_reg[1008] ),
    .S0(_1343_),
    .S1(_1276_),
    .X(_1368_));
 sky130_fd_sc_hd__mux4_1 _3702_ (.A0(_1365_),
    .A1(_1366_),
    .A2(_1367_),
    .A3(_1368_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_1 _3703_ (.A0(_1364_),
    .A1(_1369_),
    .S(_1282_),
    .X(net54));
 sky130_fd_sc_hd__mux2_1 _3704_ (.A0(\rf_reg[49] ),
    .A1(\rf_reg[113] ),
    .S(_1320_),
    .X(_1370_));
 sky130_fd_sc_hd__a22o_1 _3705_ (.A1(\rf_reg[81] ),
    .A2(_1241_),
    .B1(_1370_),
    .B2(_1246_),
    .X(_1371_));
 sky130_fd_sc_hd__buf_6 _3706_ (.A(_1242_),
    .X(_1372_));
 sky130_fd_sc_hd__mux4_1 _3707_ (.A0(\rf_reg[145] ),
    .A1(\rf_reg[177] ),
    .A2(\rf_reg[209] ),
    .A3(\rf_reg[241] ),
    .S0(_1309_),
    .S1(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__mux4_1 _3708_ (.A0(\rf_reg[529] ),
    .A1(\rf_reg[561] ),
    .A2(\rf_reg[593] ),
    .A3(\rf_reg[625] ),
    .S0(_1361_),
    .S1(_1298_),
    .X(_1374_));
 sky130_fd_sc_hd__buf_6 _3709_ (.A(_1259_),
    .X(_1375_));
 sky130_fd_sc_hd__mux4_1 _3710_ (.A0(\rf_reg[657] ),
    .A1(\rf_reg[689] ),
    .A2(\rf_reg[721] ),
    .A3(\rf_reg[753] ),
    .S0(_1312_),
    .S1(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__buf_8 _3711_ (.A(_1262_),
    .X(_1377_));
 sky130_fd_sc_hd__buf_6 _3712_ (.A(_1264_),
    .X(_1378_));
 sky130_fd_sc_hd__mux4_1 _3713_ (.A0(_1371_),
    .A1(_1373_),
    .A2(_1374_),
    .A3(_1376_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__mux4_1 _3714_ (.A0(\rf_reg[273] ),
    .A1(\rf_reg[305] ),
    .A2(\rf_reg[337] ),
    .A3(\rf_reg[369] ),
    .S0(_1289_),
    .S1(_1352_),
    .X(_1380_));
 sky130_fd_sc_hd__mux4_1 _3715_ (.A0(\rf_reg[401] ),
    .A1(\rf_reg[433] ),
    .A2(\rf_reg[465] ),
    .A3(\rf_reg[497] ),
    .S0(_1340_),
    .S1(_1271_),
    .X(_1381_));
 sky130_fd_sc_hd__mux4_1 _3716_ (.A0(\rf_reg[785] ),
    .A1(\rf_reg[817] ),
    .A2(\rf_reg[849] ),
    .A3(\rf_reg[881] ),
    .S0(_1273_),
    .S1(_1329_),
    .X(_1382_));
 sky130_fd_sc_hd__mux4_1 _3717_ (.A0(\rf_reg[913] ),
    .A1(\rf_reg[945] ),
    .A2(\rf_reg[977] ),
    .A3(\rf_reg[1009] ),
    .S0(_1343_),
    .S1(_1276_),
    .X(_1383_));
 sky130_fd_sc_hd__mux4_1 _3718_ (.A0(_1380_),
    .A1(_1381_),
    .A2(_1382_),
    .A3(_1383_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_2 _3719_ (.A0(_1379_),
    .A1(_1384_),
    .S(_1282_),
    .X(net55));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(\rf_reg[50] ),
    .A1(\rf_reg[114] ),
    .S(_1320_),
    .X(_1385_));
 sky130_fd_sc_hd__a22o_1 _3721_ (.A1(\rf_reg[82] ),
    .A2(_1241_),
    .B1(_1385_),
    .B2(_1246_),
    .X(_1386_));
 sky130_fd_sc_hd__mux4_1 _3722_ (.A0(\rf_reg[146] ),
    .A1(\rf_reg[178] ),
    .A2(\rf_reg[210] ),
    .A3(\rf_reg[242] ),
    .S0(_1309_),
    .S1(_1372_),
    .X(_1387_));
 sky130_fd_sc_hd__mux4_1 _3723_ (.A0(\rf_reg[530] ),
    .A1(\rf_reg[562] ),
    .A2(\rf_reg[594] ),
    .A3(\rf_reg[626] ),
    .S0(_1361_),
    .S1(_1298_),
    .X(_1388_));
 sky130_fd_sc_hd__mux4_1 _3724_ (.A0(\rf_reg[658] ),
    .A1(\rf_reg[690] ),
    .A2(\rf_reg[722] ),
    .A3(\rf_reg[754] ),
    .S0(_1312_),
    .S1(_1375_),
    .X(_1389_));
 sky130_fd_sc_hd__mux4_1 _3725_ (.A0(_1386_),
    .A1(_1387_),
    .A2(_1388_),
    .A3(_1389_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1390_));
 sky130_fd_sc_hd__mux4_1 _3726_ (.A0(\rf_reg[274] ),
    .A1(\rf_reg[306] ),
    .A2(\rf_reg[338] ),
    .A3(\rf_reg[370] ),
    .S0(_1289_),
    .S1(_1352_),
    .X(_1391_));
 sky130_fd_sc_hd__mux4_1 _3727_ (.A0(\rf_reg[402] ),
    .A1(\rf_reg[434] ),
    .A2(\rf_reg[466] ),
    .A3(\rf_reg[498] ),
    .S0(_1340_),
    .S1(_1271_),
    .X(_1392_));
 sky130_fd_sc_hd__buf_16 _3728_ (.A(_1248_),
    .X(_1393_));
 sky130_fd_sc_hd__mux4_1 _3729_ (.A0(\rf_reg[786] ),
    .A1(\rf_reg[818] ),
    .A2(\rf_reg[850] ),
    .A3(\rf_reg[882] ),
    .S0(_1393_),
    .S1(_1329_),
    .X(_1394_));
 sky130_fd_sc_hd__mux4_1 _3730_ (.A0(\rf_reg[914] ),
    .A1(\rf_reg[946] ),
    .A2(\rf_reg[978] ),
    .A3(\rf_reg[1010] ),
    .S0(_1343_),
    .S1(_1276_),
    .X(_1395_));
 sky130_fd_sc_hd__mux4_1 _3731_ (.A0(_1391_),
    .A1(_1392_),
    .A2(_1394_),
    .A3(_1395_),
    .S0(_1278_),
    .S1(_1279_),
    .X(_1396_));
 sky130_fd_sc_hd__mux2_2 _3732_ (.A0(_1390_),
    .A1(_1396_),
    .S(_1282_),
    .X(net56));
 sky130_fd_sc_hd__buf_6 _3733_ (.A(_1240_),
    .X(_1397_));
 sky130_fd_sc_hd__mux2_1 _3734_ (.A0(\rf_reg[51] ),
    .A1(\rf_reg[115] ),
    .S(_1320_),
    .X(_1398_));
 sky130_fd_sc_hd__buf_6 _3735_ (.A(_1245_),
    .X(_1399_));
 sky130_fd_sc_hd__a22o_1 _3736_ (.A1(\rf_reg[83] ),
    .A2(_1397_),
    .B1(_1398_),
    .B2(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__mux4_1 _3737_ (.A0(\rf_reg[147] ),
    .A1(\rf_reg[179] ),
    .A2(\rf_reg[211] ),
    .A3(\rf_reg[243] ),
    .S0(_1309_),
    .S1(_1372_),
    .X(_1401_));
 sky130_fd_sc_hd__mux4_1 _3738_ (.A0(\rf_reg[531] ),
    .A1(\rf_reg[563] ),
    .A2(\rf_reg[595] ),
    .A3(\rf_reg[627] ),
    .S0(_1361_),
    .S1(_1298_),
    .X(_1402_));
 sky130_fd_sc_hd__mux4_1 _3739_ (.A0(\rf_reg[659] ),
    .A1(\rf_reg[691] ),
    .A2(\rf_reg[723] ),
    .A3(\rf_reg[755] ),
    .S0(_1312_),
    .S1(_1375_),
    .X(_1403_));
 sky130_fd_sc_hd__mux4_1 _3740_ (.A0(_1400_),
    .A1(_1401_),
    .A2(_1402_),
    .A3(_1403_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1404_));
 sky130_fd_sc_hd__mux4_1 _3741_ (.A0(\rf_reg[275] ),
    .A1(\rf_reg[307] ),
    .A2(\rf_reg[339] ),
    .A3(\rf_reg[371] ),
    .S0(_1289_),
    .S1(_1352_),
    .X(_1405_));
 sky130_fd_sc_hd__buf_16 _3742_ (.A(_1242_),
    .X(_1406_));
 sky130_fd_sc_hd__mux4_1 _3743_ (.A0(\rf_reg[403] ),
    .A1(\rf_reg[435] ),
    .A2(\rf_reg[467] ),
    .A3(\rf_reg[499] ),
    .S0(_1340_),
    .S1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__mux4_1 _3744_ (.A0(\rf_reg[787] ),
    .A1(\rf_reg[819] ),
    .A2(\rf_reg[851] ),
    .A3(\rf_reg[883] ),
    .S0(_1393_),
    .S1(_1329_),
    .X(_1408_));
 sky130_fd_sc_hd__buf_8 _3745_ (.A(_1259_),
    .X(_1409_));
 sky130_fd_sc_hd__mux4_1 _3746_ (.A0(\rf_reg[915] ),
    .A1(\rf_reg[947] ),
    .A2(\rf_reg[979] ),
    .A3(\rf_reg[1011] ),
    .S0(_1343_),
    .S1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__buf_16 _3747_ (.A(_1262_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_16 _3748_ (.A(_1264_),
    .X(_1412_));
 sky130_fd_sc_hd__mux4_1 _3749_ (.A0(_1405_),
    .A1(_1407_),
    .A2(_1408_),
    .A3(_1410_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__buf_8 _3750_ (.A(_1281_),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_1 _3751_ (.A0(_1404_),
    .A1(_1413_),
    .S(_1414_),
    .X(net57));
 sky130_fd_sc_hd__mux2_1 _3752_ (.A0(\rf_reg[33] ),
    .A1(\rf_reg[97] ),
    .S(_1320_),
    .X(_1415_));
 sky130_fd_sc_hd__a22o_1 _3753_ (.A1(\rf_reg[65] ),
    .A2(_1397_),
    .B1(_1415_),
    .B2(_1399_),
    .X(_1416_));
 sky130_fd_sc_hd__mux4_1 _3754_ (.A0(\rf_reg[129] ),
    .A1(\rf_reg[161] ),
    .A2(\rf_reg[193] ),
    .A3(\rf_reg[225] ),
    .S0(_1309_),
    .S1(_1372_),
    .X(_1417_));
 sky130_fd_sc_hd__mux4_1 _3755_ (.A0(\rf_reg[513] ),
    .A1(\rf_reg[545] ),
    .A2(\rf_reg[577] ),
    .A3(\rf_reg[609] ),
    .S0(_1361_),
    .S1(_1298_),
    .X(_1418_));
 sky130_fd_sc_hd__mux4_1 _3756_ (.A0(\rf_reg[641] ),
    .A1(\rf_reg[673] ),
    .A2(\rf_reg[705] ),
    .A3(\rf_reg[737] ),
    .S0(_1312_),
    .S1(_1375_),
    .X(_1419_));
 sky130_fd_sc_hd__mux4_1 _3757_ (.A0(_1416_),
    .A1(_1417_),
    .A2(_1418_),
    .A3(_1419_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_16 _3758_ (.A(_1257_),
    .X(_1421_));
 sky130_fd_sc_hd__mux4_1 _3759_ (.A0(\rf_reg[257] ),
    .A1(\rf_reg[289] ),
    .A2(\rf_reg[321] ),
    .A3(\rf_reg[353] ),
    .S0(_1421_),
    .S1(_1352_),
    .X(_1422_));
 sky130_fd_sc_hd__mux4_1 _3760_ (.A0(\rf_reg[385] ),
    .A1(\rf_reg[417] ),
    .A2(\rf_reg[449] ),
    .A3(\rf_reg[481] ),
    .S0(_1340_),
    .S1(_1406_),
    .X(_1423_));
 sky130_fd_sc_hd__mux4_1 _3761_ (.A0(\rf_reg[769] ),
    .A1(\rf_reg[801] ),
    .A2(\rf_reg[833] ),
    .A3(\rf_reg[865] ),
    .S0(_1393_),
    .S1(_1329_),
    .X(_1424_));
 sky130_fd_sc_hd__mux4_1 _3762_ (.A0(\rf_reg[897] ),
    .A1(\rf_reg[929] ),
    .A2(\rf_reg[961] ),
    .A3(\rf_reg[993] ),
    .S0(_1343_),
    .S1(_1409_),
    .X(_1425_));
 sky130_fd_sc_hd__mux4_1 _3763_ (.A0(_1422_),
    .A1(_1423_),
    .A2(_1424_),
    .A3(_1425_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1426_));
 sky130_fd_sc_hd__mux2_2 _3764_ (.A0(_1420_),
    .A1(_1426_),
    .S(_1414_),
    .X(net58));
 sky130_fd_sc_hd__mux2_1 _3765_ (.A0(\rf_reg[52] ),
    .A1(\rf_reg[116] ),
    .S(_1320_),
    .X(_1427_));
 sky130_fd_sc_hd__a22o_1 _3766_ (.A1(\rf_reg[84] ),
    .A2(_1397_),
    .B1(_1427_),
    .B2(_1399_),
    .X(_1428_));
 sky130_fd_sc_hd__mux4_1 _3767_ (.A0(\rf_reg[148] ),
    .A1(\rf_reg[180] ),
    .A2(\rf_reg[212] ),
    .A3(\rf_reg[244] ),
    .S0(_1309_),
    .S1(_1372_),
    .X(_1429_));
 sky130_fd_sc_hd__buf_6 _3768_ (.A(_1254_),
    .X(_1430_));
 sky130_fd_sc_hd__mux4_1 _3769_ (.A0(\rf_reg[532] ),
    .A1(\rf_reg[564] ),
    .A2(\rf_reg[596] ),
    .A3(\rf_reg[628] ),
    .S0(_1361_),
    .S1(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__mux4_1 _3770_ (.A0(\rf_reg[660] ),
    .A1(\rf_reg[692] ),
    .A2(\rf_reg[724] ),
    .A3(\rf_reg[756] ),
    .S0(_1312_),
    .S1(_1375_),
    .X(_1432_));
 sky130_fd_sc_hd__mux4_1 _3771_ (.A0(_1428_),
    .A1(_1429_),
    .A2(_1431_),
    .A3(_1432_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1433_));
 sky130_fd_sc_hd__mux4_1 _3772_ (.A0(\rf_reg[276] ),
    .A1(\rf_reg[308] ),
    .A2(\rf_reg[340] ),
    .A3(\rf_reg[372] ),
    .S0(_1421_),
    .S1(_1352_),
    .X(_1434_));
 sky130_fd_sc_hd__mux4_1 _3773_ (.A0(\rf_reg[404] ),
    .A1(\rf_reg[436] ),
    .A2(\rf_reg[468] ),
    .A3(\rf_reg[500] ),
    .S0(_1340_),
    .S1(_1406_),
    .X(_1435_));
 sky130_fd_sc_hd__mux4_1 _3774_ (.A0(\rf_reg[788] ),
    .A1(\rf_reg[820] ),
    .A2(\rf_reg[852] ),
    .A3(\rf_reg[884] ),
    .S0(_1393_),
    .S1(_1329_),
    .X(_1436_));
 sky130_fd_sc_hd__mux4_1 _3775_ (.A0(\rf_reg[916] ),
    .A1(\rf_reg[948] ),
    .A2(\rf_reg[980] ),
    .A3(\rf_reg[1012] ),
    .S0(_1343_),
    .S1(_1409_),
    .X(_1437_));
 sky130_fd_sc_hd__mux4_1 _3776_ (.A0(_1434_),
    .A1(_1435_),
    .A2(_1436_),
    .A3(_1437_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1438_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(_1433_),
    .A1(_1438_),
    .S(_1414_),
    .X(net59));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(\rf_reg[53] ),
    .A1(\rf_reg[117] ),
    .S(_1320_),
    .X(_1439_));
 sky130_fd_sc_hd__a22o_1 _3779_ (.A1(\rf_reg[85] ),
    .A2(_1397_),
    .B1(_1439_),
    .B2(_1399_),
    .X(_1440_));
 sky130_fd_sc_hd__buf_8 _3780_ (.A(_1237_),
    .X(_1441_));
 sky130_fd_sc_hd__mux4_1 _3781_ (.A0(\rf_reg[149] ),
    .A1(\rf_reg[181] ),
    .A2(\rf_reg[213] ),
    .A3(\rf_reg[245] ),
    .S0(_1441_),
    .S1(_1372_),
    .X(_1442_));
 sky130_fd_sc_hd__mux4_1 _3782_ (.A0(\rf_reg[533] ),
    .A1(\rf_reg[565] ),
    .A2(\rf_reg[597] ),
    .A3(\rf_reg[629] ),
    .S0(_1361_),
    .S1(_1430_),
    .X(_1443_));
 sky130_fd_sc_hd__buf_16 _3783_ (.A(_1257_),
    .X(_1444_));
 sky130_fd_sc_hd__mux4_1 _3784_ (.A0(\rf_reg[661] ),
    .A1(\rf_reg[693] ),
    .A2(\rf_reg[725] ),
    .A3(\rf_reg[757] ),
    .S0(_1444_),
    .S1(_1375_),
    .X(_1445_));
 sky130_fd_sc_hd__mux4_1 _3785_ (.A0(_1440_),
    .A1(_1442_),
    .A2(_1443_),
    .A3(_1445_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1446_));
 sky130_fd_sc_hd__mux4_1 _3786_ (.A0(\rf_reg[277] ),
    .A1(\rf_reg[309] ),
    .A2(\rf_reg[341] ),
    .A3(\rf_reg[373] ),
    .S0(_1421_),
    .S1(_1352_),
    .X(_1447_));
 sky130_fd_sc_hd__mux4_1 _3787_ (.A0(\rf_reg[405] ),
    .A1(\rf_reg[437] ),
    .A2(\rf_reg[469] ),
    .A3(\rf_reg[501] ),
    .S0(_1340_),
    .S1(_1406_),
    .X(_1448_));
 sky130_fd_sc_hd__mux4_1 _3788_ (.A0(\rf_reg[789] ),
    .A1(\rf_reg[821] ),
    .A2(\rf_reg[853] ),
    .A3(\rf_reg[885] ),
    .S0(_1393_),
    .S1(_1329_),
    .X(_1449_));
 sky130_fd_sc_hd__mux4_1 _3789_ (.A0(\rf_reg[917] ),
    .A1(\rf_reg[949] ),
    .A2(\rf_reg[981] ),
    .A3(\rf_reg[1013] ),
    .S0(_1343_),
    .S1(_1409_),
    .X(_1450_));
 sky130_fd_sc_hd__mux4_1 _3790_ (.A0(_1447_),
    .A1(_1448_),
    .A2(_1449_),
    .A3(_1450_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(_1446_),
    .A1(_1451_),
    .S(_1414_),
    .X(net60));
 sky130_fd_sc_hd__buf_6 _3792_ (.A(_1238_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(\rf_reg[54] ),
    .A1(\rf_reg[118] ),
    .S(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__a22o_1 _3794_ (.A1(\rf_reg[86] ),
    .A2(_1397_),
    .B1(_1453_),
    .B2(_1399_),
    .X(_1454_));
 sky130_fd_sc_hd__mux4_1 _3795_ (.A0(\rf_reg[150] ),
    .A1(\rf_reg[182] ),
    .A2(\rf_reg[214] ),
    .A3(\rf_reg[246] ),
    .S0(_1441_),
    .S1(_1372_),
    .X(_1455_));
 sky130_fd_sc_hd__mux4_1 _3796_ (.A0(\rf_reg[534] ),
    .A1(\rf_reg[566] ),
    .A2(\rf_reg[598] ),
    .A3(\rf_reg[630] ),
    .S0(_1361_),
    .S1(_1430_),
    .X(_1456_));
 sky130_fd_sc_hd__mux4_1 _3797_ (.A0(\rf_reg[662] ),
    .A1(\rf_reg[694] ),
    .A2(\rf_reg[726] ),
    .A3(\rf_reg[758] ),
    .S0(_1444_),
    .S1(_1375_),
    .X(_1457_));
 sky130_fd_sc_hd__mux4_1 _3798_ (.A0(_1454_),
    .A1(_1455_),
    .A2(_1456_),
    .A3(_1457_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1458_));
 sky130_fd_sc_hd__mux4_1 _3799_ (.A0(\rf_reg[278] ),
    .A1(\rf_reg[310] ),
    .A2(\rf_reg[342] ),
    .A3(\rf_reg[374] ),
    .S0(_1421_),
    .S1(_1352_),
    .X(_1459_));
 sky130_fd_sc_hd__mux4_1 _3800_ (.A0(\rf_reg[406] ),
    .A1(\rf_reg[438] ),
    .A2(\rf_reg[470] ),
    .A3(\rf_reg[502] ),
    .S0(_1340_),
    .S1(_1406_),
    .X(_1460_));
 sky130_fd_sc_hd__buf_8 _3801_ (.A(_1254_),
    .X(_1461_));
 sky130_fd_sc_hd__mux4_1 _3802_ (.A0(\rf_reg[790] ),
    .A1(\rf_reg[822] ),
    .A2(\rf_reg[854] ),
    .A3(\rf_reg[886] ),
    .S0(_1393_),
    .S1(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__mux4_1 _3803_ (.A0(\rf_reg[918] ),
    .A1(\rf_reg[950] ),
    .A2(\rf_reg[982] ),
    .A3(\rf_reg[1014] ),
    .S0(_1343_),
    .S1(_1409_),
    .X(_1463_));
 sky130_fd_sc_hd__mux4_1 _3804_ (.A0(_1459_),
    .A1(_1460_),
    .A2(_1462_),
    .A3(_1463_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _3805_ (.A0(_1458_),
    .A1(_1464_),
    .S(_1414_),
    .X(net61));
 sky130_fd_sc_hd__mux2_1 _3806_ (.A0(\rf_reg[55] ),
    .A1(\rf_reg[119] ),
    .S(_1452_),
    .X(_1465_));
 sky130_fd_sc_hd__a22o_1 _3807_ (.A1(\rf_reg[87] ),
    .A2(_1397_),
    .B1(_1465_),
    .B2(_1399_),
    .X(_1466_));
 sky130_fd_sc_hd__mux4_2 _3808_ (.A0(\rf_reg[151] ),
    .A1(\rf_reg[183] ),
    .A2(\rf_reg[215] ),
    .A3(\rf_reg[247] ),
    .S0(_1441_),
    .S1(_1372_),
    .X(_1467_));
 sky130_fd_sc_hd__mux4_1 _3809_ (.A0(\rf_reg[535] ),
    .A1(\rf_reg[567] ),
    .A2(\rf_reg[599] ),
    .A3(\rf_reg[631] ),
    .S0(_1361_),
    .S1(_1430_),
    .X(_1468_));
 sky130_fd_sc_hd__mux4_1 _3810_ (.A0(\rf_reg[663] ),
    .A1(\rf_reg[695] ),
    .A2(\rf_reg[727] ),
    .A3(\rf_reg[759] ),
    .S0(_1444_),
    .S1(_1375_),
    .X(_1469_));
 sky130_fd_sc_hd__mux4_1 _3811_ (.A0(_1466_),
    .A1(_1467_),
    .A2(_1468_),
    .A3(_1469_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1470_));
 sky130_fd_sc_hd__mux4_1 _3812_ (.A0(\rf_reg[279] ),
    .A1(\rf_reg[311] ),
    .A2(\rf_reg[343] ),
    .A3(\rf_reg[375] ),
    .S0(_1421_),
    .S1(_1352_),
    .X(_1471_));
 sky130_fd_sc_hd__buf_8 _3813_ (.A(_1248_),
    .X(_1472_));
 sky130_fd_sc_hd__mux4_1 _3814_ (.A0(\rf_reg[407] ),
    .A1(\rf_reg[439] ),
    .A2(\rf_reg[471] ),
    .A3(\rf_reg[503] ),
    .S0(_1472_),
    .S1(_1406_),
    .X(_1473_));
 sky130_fd_sc_hd__mux4_1 _3815_ (.A0(\rf_reg[791] ),
    .A1(\rf_reg[823] ),
    .A2(\rf_reg[855] ),
    .A3(\rf_reg[887] ),
    .S0(_1393_),
    .S1(_1461_),
    .X(_1474_));
 sky130_fd_sc_hd__buf_16 _3816_ (.A(_1257_),
    .X(_1475_));
 sky130_fd_sc_hd__mux4_1 _3817_ (.A0(\rf_reg[919] ),
    .A1(\rf_reg[951] ),
    .A2(\rf_reg[983] ),
    .A3(\rf_reg[1015] ),
    .S0(_1475_),
    .S1(_1409_),
    .X(_1476_));
 sky130_fd_sc_hd__mux4_1 _3818_ (.A0(_1471_),
    .A1(_1473_),
    .A2(_1474_),
    .A3(_1476_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _3819_ (.A0(_1470_),
    .A1(_1477_),
    .S(_1414_),
    .X(net62));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(\rf_reg[56] ),
    .A1(\rf_reg[120] ),
    .S(_1452_),
    .X(_1478_));
 sky130_fd_sc_hd__a22o_1 _3821_ (.A1(\rf_reg[88] ),
    .A2(_1397_),
    .B1(_1478_),
    .B2(_1399_),
    .X(_1479_));
 sky130_fd_sc_hd__mux4_2 _3822_ (.A0(\rf_reg[152] ),
    .A1(\rf_reg[184] ),
    .A2(\rf_reg[216] ),
    .A3(\rf_reg[248] ),
    .S0(_1441_),
    .S1(_1372_),
    .X(_1480_));
 sky130_fd_sc_hd__mux4_1 _3823_ (.A0(\rf_reg[536] ),
    .A1(\rf_reg[568] ),
    .A2(\rf_reg[600] ),
    .A3(\rf_reg[632] ),
    .S0(_1361_),
    .S1(_1430_),
    .X(_1481_));
 sky130_fd_sc_hd__mux4_1 _3824_ (.A0(\rf_reg[664] ),
    .A1(\rf_reg[696] ),
    .A2(\rf_reg[728] ),
    .A3(\rf_reg[760] ),
    .S0(_1444_),
    .S1(_1375_),
    .X(_1482_));
 sky130_fd_sc_hd__mux4_1 _3825_ (.A0(_1479_),
    .A1(_1480_),
    .A2(_1481_),
    .A3(_1482_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1483_));
 sky130_fd_sc_hd__buf_8 _3826_ (.A(_1254_),
    .X(_1484_));
 sky130_fd_sc_hd__mux4_1 _3827_ (.A0(\rf_reg[280] ),
    .A1(\rf_reg[312] ),
    .A2(\rf_reg[344] ),
    .A3(\rf_reg[376] ),
    .S0(_1421_),
    .S1(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__mux4_1 _3828_ (.A0(\rf_reg[408] ),
    .A1(\rf_reg[440] ),
    .A2(\rf_reg[472] ),
    .A3(\rf_reg[504] ),
    .S0(_1472_),
    .S1(_1406_),
    .X(_1486_));
 sky130_fd_sc_hd__mux4_1 _3829_ (.A0(\rf_reg[792] ),
    .A1(\rf_reg[824] ),
    .A2(\rf_reg[856] ),
    .A3(\rf_reg[888] ),
    .S0(_1393_),
    .S1(_1461_),
    .X(_1487_));
 sky130_fd_sc_hd__mux4_1 _3830_ (.A0(\rf_reg[920] ),
    .A1(\rf_reg[952] ),
    .A2(\rf_reg[984] ),
    .A3(\rf_reg[1016] ),
    .S0(_1475_),
    .S1(_1409_),
    .X(_1488_));
 sky130_fd_sc_hd__mux4_1 _3831_ (.A0(_1485_),
    .A1(_1486_),
    .A2(_1487_),
    .A3(_1488_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_2 _3832_ (.A0(_1483_),
    .A1(_1489_),
    .S(_1414_),
    .X(net63));
 sky130_fd_sc_hd__mux2_1 _3833_ (.A0(\rf_reg[57] ),
    .A1(\rf_reg[121] ),
    .S(_1452_),
    .X(_1490_));
 sky130_fd_sc_hd__a22o_1 _3834_ (.A1(\rf_reg[89] ),
    .A2(_1397_),
    .B1(_1490_),
    .B2(_1399_),
    .X(_1491_));
 sky130_fd_sc_hd__mux4_2 _3835_ (.A0(\rf_reg[153] ),
    .A1(\rf_reg[185] ),
    .A2(\rf_reg[217] ),
    .A3(\rf_reg[249] ),
    .S0(_1441_),
    .S1(_1372_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_16 _3836_ (.A(_1248_),
    .X(_1493_));
 sky130_fd_sc_hd__mux4_1 _3837_ (.A0(\rf_reg[537] ),
    .A1(\rf_reg[569] ),
    .A2(\rf_reg[601] ),
    .A3(\rf_reg[633] ),
    .S0(_1493_),
    .S1(_1430_),
    .X(_1494_));
 sky130_fd_sc_hd__mux4_1 _3838_ (.A0(\rf_reg[665] ),
    .A1(\rf_reg[697] ),
    .A2(\rf_reg[729] ),
    .A3(\rf_reg[761] ),
    .S0(_1444_),
    .S1(_1375_),
    .X(_1495_));
 sky130_fd_sc_hd__mux4_1 _3839_ (.A0(_1491_),
    .A1(_1492_),
    .A2(_1494_),
    .A3(_1495_),
    .S0(_1377_),
    .S1(_1378_),
    .X(_1496_));
 sky130_fd_sc_hd__mux4_1 _3840_ (.A0(\rf_reg[281] ),
    .A1(\rf_reg[313] ),
    .A2(\rf_reg[345] ),
    .A3(\rf_reg[377] ),
    .S0(_1421_),
    .S1(_1484_),
    .X(_1497_));
 sky130_fd_sc_hd__mux4_1 _3841_ (.A0(\rf_reg[409] ),
    .A1(\rf_reg[441] ),
    .A2(\rf_reg[473] ),
    .A3(\rf_reg[505] ),
    .S0(_1472_),
    .S1(_1406_),
    .X(_1498_));
 sky130_fd_sc_hd__mux4_1 _3842_ (.A0(\rf_reg[793] ),
    .A1(\rf_reg[825] ),
    .A2(\rf_reg[857] ),
    .A3(\rf_reg[889] ),
    .S0(_1393_),
    .S1(_1461_),
    .X(_1499_));
 sky130_fd_sc_hd__mux4_1 _3843_ (.A0(\rf_reg[921] ),
    .A1(\rf_reg[953] ),
    .A2(\rf_reg[985] ),
    .A3(\rf_reg[1017] ),
    .S0(_1475_),
    .S1(_1409_),
    .X(_1500_));
 sky130_fd_sc_hd__mux4_1 _3844_ (.A0(_1497_),
    .A1(_1498_),
    .A2(_1499_),
    .A3(_1500_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(_1496_),
    .A1(_1501_),
    .S(_1414_),
    .X(net64));
 sky130_fd_sc_hd__mux2_1 _3846_ (.A0(\rf_reg[58] ),
    .A1(\rf_reg[122] ),
    .S(_1452_),
    .X(_1502_));
 sky130_fd_sc_hd__a22o_1 _3847_ (.A1(\rf_reg[90] ),
    .A2(_1397_),
    .B1(_1502_),
    .B2(_1399_),
    .X(_1503_));
 sky130_fd_sc_hd__buf_6 _3848_ (.A(_1242_),
    .X(_1504_));
 sky130_fd_sc_hd__mux4_2 _3849_ (.A0(\rf_reg[154] ),
    .A1(\rf_reg[186] ),
    .A2(\rf_reg[218] ),
    .A3(\rf_reg[250] ),
    .S0(_1441_),
    .S1(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__mux4_1 _3850_ (.A0(\rf_reg[538] ),
    .A1(\rf_reg[570] ),
    .A2(\rf_reg[602] ),
    .A3(\rf_reg[634] ),
    .S0(_1493_),
    .S1(_1430_),
    .X(_1506_));
 sky130_fd_sc_hd__buf_8 _3851_ (.A(_1259_),
    .X(_1507_));
 sky130_fd_sc_hd__mux4_1 _3852_ (.A0(\rf_reg[666] ),
    .A1(\rf_reg[698] ),
    .A2(\rf_reg[730] ),
    .A3(\rf_reg[762] ),
    .S0(_1444_),
    .S1(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_16 _3853_ (.A(_1262_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_16 _3854_ (.A(_1264_),
    .X(_1510_));
 sky130_fd_sc_hd__mux4_1 _3855_ (.A0(_1503_),
    .A1(_1505_),
    .A2(_1506_),
    .A3(_1508_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__mux4_1 _3856_ (.A0(\rf_reg[282] ),
    .A1(\rf_reg[314] ),
    .A2(\rf_reg[346] ),
    .A3(\rf_reg[378] ),
    .S0(_1421_),
    .S1(_1484_),
    .X(_1512_));
 sky130_fd_sc_hd__mux4_1 _3857_ (.A0(\rf_reg[410] ),
    .A1(\rf_reg[442] ),
    .A2(\rf_reg[474] ),
    .A3(\rf_reg[506] ),
    .S0(_1472_),
    .S1(_1406_),
    .X(_1513_));
 sky130_fd_sc_hd__mux4_1 _3858_ (.A0(\rf_reg[794] ),
    .A1(\rf_reg[826] ),
    .A2(\rf_reg[858] ),
    .A3(\rf_reg[890] ),
    .S0(_1393_),
    .S1(_1461_),
    .X(_1514_));
 sky130_fd_sc_hd__mux4_1 _3859_ (.A0(\rf_reg[922] ),
    .A1(\rf_reg[954] ),
    .A2(\rf_reg[986] ),
    .A3(\rf_reg[1018] ),
    .S0(_1475_),
    .S1(_1409_),
    .X(_1515_));
 sky130_fd_sc_hd__mux4_1 _3860_ (.A0(_1512_),
    .A1(_1513_),
    .A2(_1514_),
    .A3(_1515_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _3861_ (.A0(_1511_),
    .A1(_1516_),
    .S(_1414_),
    .X(net65));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(\rf_reg[59] ),
    .A1(\rf_reg[123] ),
    .S(_1452_),
    .X(_1517_));
 sky130_fd_sc_hd__a22o_1 _3863_ (.A1(\rf_reg[91] ),
    .A2(_1397_),
    .B1(_1517_),
    .B2(_1399_),
    .X(_1518_));
 sky130_fd_sc_hd__mux4_2 _3864_ (.A0(\rf_reg[155] ),
    .A1(\rf_reg[187] ),
    .A2(\rf_reg[219] ),
    .A3(\rf_reg[251] ),
    .S0(_1441_),
    .S1(_1504_),
    .X(_1519_));
 sky130_fd_sc_hd__mux4_1 _3865_ (.A0(\rf_reg[539] ),
    .A1(\rf_reg[571] ),
    .A2(\rf_reg[603] ),
    .A3(\rf_reg[635] ),
    .S0(_1493_),
    .S1(_1430_),
    .X(_1520_));
 sky130_fd_sc_hd__mux4_1 _3866_ (.A0(\rf_reg[667] ),
    .A1(\rf_reg[699] ),
    .A2(\rf_reg[731] ),
    .A3(\rf_reg[763] ),
    .S0(_1444_),
    .S1(_1507_),
    .X(_1521_));
 sky130_fd_sc_hd__mux4_1 _3867_ (.A0(_1518_),
    .A1(_1519_),
    .A2(_1520_),
    .A3(_1521_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1522_));
 sky130_fd_sc_hd__mux4_1 _3868_ (.A0(\rf_reg[283] ),
    .A1(\rf_reg[315] ),
    .A2(\rf_reg[347] ),
    .A3(\rf_reg[379] ),
    .S0(_1421_),
    .S1(_1484_),
    .X(_1523_));
 sky130_fd_sc_hd__mux4_1 _3869_ (.A0(\rf_reg[411] ),
    .A1(\rf_reg[443] ),
    .A2(\rf_reg[475] ),
    .A3(\rf_reg[507] ),
    .S0(_1472_),
    .S1(_1406_),
    .X(_1524_));
 sky130_fd_sc_hd__buf_16 _3870_ (.A(_1248_),
    .X(_1525_));
 sky130_fd_sc_hd__mux4_1 _3871_ (.A0(\rf_reg[795] ),
    .A1(\rf_reg[827] ),
    .A2(\rf_reg[859] ),
    .A3(\rf_reg[891] ),
    .S0(_1525_),
    .S1(_1461_),
    .X(_1526_));
 sky130_fd_sc_hd__mux4_1 _3872_ (.A0(\rf_reg[923] ),
    .A1(\rf_reg[955] ),
    .A2(\rf_reg[987] ),
    .A3(\rf_reg[1019] ),
    .S0(_1475_),
    .S1(_1409_),
    .X(_1527_));
 sky130_fd_sc_hd__mux4_1 _3873_ (.A0(_1523_),
    .A1(_1524_),
    .A2(_1526_),
    .A3(_1527_),
    .S0(_1411_),
    .S1(_1412_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(_1522_),
    .A1(_1528_),
    .S(_1414_),
    .X(net66));
 sky130_fd_sc_hd__buf_6 _3875_ (.A(_1240_),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(\rf_reg[60] ),
    .A1(\rf_reg[124] ),
    .S(_1452_),
    .X(_1530_));
 sky130_fd_sc_hd__buf_6 _3877_ (.A(_1245_),
    .X(_1531_));
 sky130_fd_sc_hd__a22o_1 _3878_ (.A1(\rf_reg[92] ),
    .A2(_1529_),
    .B1(_1530_),
    .B2(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__mux4_1 _3879_ (.A0(\rf_reg[156] ),
    .A1(\rf_reg[188] ),
    .A2(\rf_reg[220] ),
    .A3(\rf_reg[252] ),
    .S0(_1441_),
    .S1(_1504_),
    .X(_1533_));
 sky130_fd_sc_hd__mux4_1 _3880_ (.A0(\rf_reg[540] ),
    .A1(\rf_reg[572] ),
    .A2(\rf_reg[604] ),
    .A3(\rf_reg[636] ),
    .S0(_1493_),
    .S1(_1430_),
    .X(_1534_));
 sky130_fd_sc_hd__mux4_1 _3881_ (.A0(\rf_reg[668] ),
    .A1(\rf_reg[700] ),
    .A2(\rf_reg[732] ),
    .A3(\rf_reg[764] ),
    .S0(_1444_),
    .S1(_1507_),
    .X(_1535_));
 sky130_fd_sc_hd__mux4_1 _3882_ (.A0(_1532_),
    .A1(_1533_),
    .A2(_1534_),
    .A3(_1535_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1536_));
 sky130_fd_sc_hd__mux4_1 _3883_ (.A0(\rf_reg[284] ),
    .A1(\rf_reg[316] ),
    .A2(\rf_reg[348] ),
    .A3(\rf_reg[380] ),
    .S0(_1421_),
    .S1(_1484_),
    .X(_1537_));
 sky130_fd_sc_hd__buf_8 _3884_ (.A(_1242_),
    .X(_1538_));
 sky130_fd_sc_hd__mux4_1 _3885_ (.A0(\rf_reg[412] ),
    .A1(\rf_reg[444] ),
    .A2(\rf_reg[476] ),
    .A3(\rf_reg[508] ),
    .S0(_1472_),
    .S1(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__mux4_1 _3886_ (.A0(\rf_reg[796] ),
    .A1(\rf_reg[828] ),
    .A2(\rf_reg[860] ),
    .A3(\rf_reg[892] ),
    .S0(_1525_),
    .S1(_1461_),
    .X(_1540_));
 sky130_fd_sc_hd__buf_16 _3887_ (.A(_1259_),
    .X(_1541_));
 sky130_fd_sc_hd__mux4_1 _3888_ (.A0(\rf_reg[924] ),
    .A1(\rf_reg[956] ),
    .A2(\rf_reg[988] ),
    .A3(\rf_reg[1020] ),
    .S0(_1475_),
    .S1(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__buf_8 _3889_ (.A(_1262_),
    .X(_1543_));
 sky130_fd_sc_hd__buf_8 _3890_ (.A(_1264_),
    .X(_1544_));
 sky130_fd_sc_hd__mux4_1 _3891_ (.A0(_1537_),
    .A1(_1539_),
    .A2(_1540_),
    .A3(_1542_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_16 _3892_ (.A(_1281_),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_1 _3893_ (.A0(_1536_),
    .A1(_1545_),
    .S(_1546_),
    .X(net67));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(\rf_reg[61] ),
    .A1(\rf_reg[125] ),
    .S(_1452_),
    .X(_1547_));
 sky130_fd_sc_hd__a22o_1 _3895_ (.A1(\rf_reg[93] ),
    .A2(_1529_),
    .B1(_1547_),
    .B2(_1531_),
    .X(_1548_));
 sky130_fd_sc_hd__mux4_1 _3896_ (.A0(\rf_reg[157] ),
    .A1(\rf_reg[189] ),
    .A2(\rf_reg[221] ),
    .A3(\rf_reg[253] ),
    .S0(_1441_),
    .S1(_1504_),
    .X(_1549_));
 sky130_fd_sc_hd__mux4_1 _3897_ (.A0(\rf_reg[541] ),
    .A1(\rf_reg[573] ),
    .A2(\rf_reg[605] ),
    .A3(\rf_reg[637] ),
    .S0(_1493_),
    .S1(_1430_),
    .X(_1550_));
 sky130_fd_sc_hd__mux4_1 _3898_ (.A0(\rf_reg[669] ),
    .A1(\rf_reg[701] ),
    .A2(\rf_reg[733] ),
    .A3(\rf_reg[765] ),
    .S0(_1444_),
    .S1(_1507_),
    .X(_1551_));
 sky130_fd_sc_hd__mux4_1 _3899_ (.A0(_1548_),
    .A1(_1549_),
    .A2(_1550_),
    .A3(_1551_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1552_));
 sky130_fd_sc_hd__buf_16 _3900_ (.A(_1257_),
    .X(_1553_));
 sky130_fd_sc_hd__mux4_1 _3901_ (.A0(\rf_reg[285] ),
    .A1(\rf_reg[317] ),
    .A2(\rf_reg[349] ),
    .A3(\rf_reg[381] ),
    .S0(_1553_),
    .S1(_1484_),
    .X(_1554_));
 sky130_fd_sc_hd__mux4_1 _3902_ (.A0(\rf_reg[413] ),
    .A1(\rf_reg[445] ),
    .A2(\rf_reg[477] ),
    .A3(\rf_reg[509] ),
    .S0(_1472_),
    .S1(_1538_),
    .X(_1555_));
 sky130_fd_sc_hd__mux4_1 _3903_ (.A0(\rf_reg[797] ),
    .A1(\rf_reg[829] ),
    .A2(\rf_reg[861] ),
    .A3(\rf_reg[893] ),
    .S0(_1525_),
    .S1(_1461_),
    .X(_1556_));
 sky130_fd_sc_hd__mux4_1 _3904_ (.A0(\rf_reg[925] ),
    .A1(\rf_reg[957] ),
    .A2(\rf_reg[989] ),
    .A3(\rf_reg[1021] ),
    .S0(_1475_),
    .S1(_1541_),
    .X(_1557_));
 sky130_fd_sc_hd__mux4_1 _3905_ (.A0(_1554_),
    .A1(_1555_),
    .A2(_1556_),
    .A3(_1557_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(_1552_),
    .A1(_1558_),
    .S(_1546_),
    .X(net68));
 sky130_fd_sc_hd__mux2_1 _3907_ (.A0(\rf_reg[34] ),
    .A1(\rf_reg[98] ),
    .S(_1452_),
    .X(_1559_));
 sky130_fd_sc_hd__a22o_1 _3908_ (.A1(\rf_reg[66] ),
    .A2(_1529_),
    .B1(_1559_),
    .B2(_1531_),
    .X(_1560_));
 sky130_fd_sc_hd__mux4_1 _3909_ (.A0(\rf_reg[130] ),
    .A1(\rf_reg[162] ),
    .A2(\rf_reg[194] ),
    .A3(\rf_reg[226] ),
    .S0(_1441_),
    .S1(_1504_),
    .X(_1561_));
 sky130_fd_sc_hd__buf_8 _3910_ (.A(_1254_),
    .X(_1562_));
 sky130_fd_sc_hd__mux4_1 _3911_ (.A0(\rf_reg[514] ),
    .A1(\rf_reg[546] ),
    .A2(\rf_reg[578] ),
    .A3(\rf_reg[610] ),
    .S0(_1493_),
    .S1(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__mux4_1 _3912_ (.A0(\rf_reg[642] ),
    .A1(\rf_reg[674] ),
    .A2(\rf_reg[706] ),
    .A3(\rf_reg[738] ),
    .S0(_1444_),
    .S1(_1507_),
    .X(_1564_));
 sky130_fd_sc_hd__mux4_1 _3913_ (.A0(_1560_),
    .A1(_1561_),
    .A2(_1563_),
    .A3(_1564_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1565_));
 sky130_fd_sc_hd__mux4_1 _3914_ (.A0(\rf_reg[258] ),
    .A1(\rf_reg[290] ),
    .A2(\rf_reg[322] ),
    .A3(\rf_reg[354] ),
    .S0(_1553_),
    .S1(_1484_),
    .X(_1566_));
 sky130_fd_sc_hd__mux4_1 _3915_ (.A0(\rf_reg[386] ),
    .A1(\rf_reg[418] ),
    .A2(\rf_reg[450] ),
    .A3(\rf_reg[482] ),
    .S0(_1472_),
    .S1(_1538_),
    .X(_1567_));
 sky130_fd_sc_hd__mux4_1 _3916_ (.A0(\rf_reg[770] ),
    .A1(\rf_reg[802] ),
    .A2(\rf_reg[834] ),
    .A3(\rf_reg[866] ),
    .S0(_1525_),
    .S1(_1461_),
    .X(_1568_));
 sky130_fd_sc_hd__mux4_1 _3917_ (.A0(\rf_reg[898] ),
    .A1(\rf_reg[930] ),
    .A2(\rf_reg[962] ),
    .A3(\rf_reg[994] ),
    .S0(_1475_),
    .S1(_1541_),
    .X(_1569_));
 sky130_fd_sc_hd__mux4_1 _3918_ (.A0(_1566_),
    .A1(_1567_),
    .A2(_1568_),
    .A3(_1569_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1570_));
 sky130_fd_sc_hd__mux2_1 _3919_ (.A0(_1565_),
    .A1(_1570_),
    .S(_1546_),
    .X(net69));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(\rf_reg[62] ),
    .A1(\rf_reg[126] ),
    .S(_1452_),
    .X(_1571_));
 sky130_fd_sc_hd__a22o_1 _3921_ (.A1(\rf_reg[94] ),
    .A2(_1529_),
    .B1(_1571_),
    .B2(_1531_),
    .X(_1572_));
 sky130_fd_sc_hd__mux4_1 _3922_ (.A0(\rf_reg[158] ),
    .A1(\rf_reg[190] ),
    .A2(\rf_reg[222] ),
    .A3(\rf_reg[254] ),
    .S0(_1244_),
    .S1(_1504_),
    .X(_1573_));
 sky130_fd_sc_hd__mux4_1 _3923_ (.A0(\rf_reg[542] ),
    .A1(\rf_reg[574] ),
    .A2(\rf_reg[606] ),
    .A3(\rf_reg[638] ),
    .S0(_1493_),
    .S1(_1562_),
    .X(_1574_));
 sky130_fd_sc_hd__mux4_1 _3924_ (.A0(\rf_reg[670] ),
    .A1(\rf_reg[702] ),
    .A2(\rf_reg[734] ),
    .A3(\rf_reg[766] ),
    .S0(_1267_),
    .S1(_1507_),
    .X(_1575_));
 sky130_fd_sc_hd__mux4_1 _3925_ (.A0(_1572_),
    .A1(_1573_),
    .A2(_1574_),
    .A3(_1575_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1576_));
 sky130_fd_sc_hd__mux4_1 _3926_ (.A0(\rf_reg[286] ),
    .A1(\rf_reg[318] ),
    .A2(\rf_reg[350] ),
    .A3(\rf_reg[382] ),
    .S0(_1553_),
    .S1(_1484_),
    .X(_1577_));
 sky130_fd_sc_hd__mux4_1 _3927_ (.A0(\rf_reg[414] ),
    .A1(\rf_reg[446] ),
    .A2(\rf_reg[478] ),
    .A3(\rf_reg[510] ),
    .S0(_1472_),
    .S1(_1538_),
    .X(_1578_));
 sky130_fd_sc_hd__mux4_1 _3928_ (.A0(\rf_reg[798] ),
    .A1(\rf_reg[830] ),
    .A2(\rf_reg[862] ),
    .A3(\rf_reg[894] ),
    .S0(_1525_),
    .S1(_1461_),
    .X(_1579_));
 sky130_fd_sc_hd__mux4_1 _3929_ (.A0(\rf_reg[926] ),
    .A1(\rf_reg[958] ),
    .A2(\rf_reg[990] ),
    .A3(\rf_reg[1022] ),
    .S0(_1475_),
    .S1(_1541_),
    .X(_1580_));
 sky130_fd_sc_hd__mux4_1 _3930_ (.A0(_1577_),
    .A1(_1578_),
    .A2(_1579_),
    .A3(_1580_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1581_));
 sky130_fd_sc_hd__mux2_4 _3931_ (.A0(_1576_),
    .A1(_1581_),
    .S(_1546_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _3932_ (.A0(\rf_reg[63] ),
    .A1(\rf_reg[127] ),
    .S(_1253_),
    .X(_1582_));
 sky130_fd_sc_hd__a22o_1 _3933_ (.A1(\rf_reg[95] ),
    .A2(_1529_),
    .B1(_1582_),
    .B2(_1531_),
    .X(_1583_));
 sky130_fd_sc_hd__mux4_1 _3934_ (.A0(\rf_reg[159] ),
    .A1(\rf_reg[191] ),
    .A2(\rf_reg[223] ),
    .A3(\rf_reg[255] ),
    .S0(_1244_),
    .S1(_1504_),
    .X(_1584_));
 sky130_fd_sc_hd__mux4_1 _3935_ (.A0(\rf_reg[543] ),
    .A1(\rf_reg[575] ),
    .A2(\rf_reg[607] ),
    .A3(\rf_reg[639] ),
    .S0(_1493_),
    .S1(_1562_),
    .X(_1585_));
 sky130_fd_sc_hd__mux4_1 _3936_ (.A0(\rf_reg[671] ),
    .A1(\rf_reg[703] ),
    .A2(\rf_reg[735] ),
    .A3(\rf_reg[767] ),
    .S0(_1267_),
    .S1(_1507_),
    .X(_1586_));
 sky130_fd_sc_hd__mux4_1 _3937_ (.A0(_1583_),
    .A1(_1584_),
    .A2(_1585_),
    .A3(_1586_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1587_));
 sky130_fd_sc_hd__mux4_1 _3938_ (.A0(\rf_reg[287] ),
    .A1(\rf_reg[319] ),
    .A2(\rf_reg[351] ),
    .A3(\rf_reg[383] ),
    .S0(_1553_),
    .S1(_1484_),
    .X(_1588_));
 sky130_fd_sc_hd__mux4_1 _3939_ (.A0(\rf_reg[415] ),
    .A1(\rf_reg[447] ),
    .A2(\rf_reg[479] ),
    .A3(\rf_reg[511] ),
    .S0(_1472_),
    .S1(_1538_),
    .X(_1589_));
 sky130_fd_sc_hd__mux4_1 _3940_ (.A0(\rf_reg[799] ),
    .A1(\rf_reg[831] ),
    .A2(\rf_reg[863] ),
    .A3(\rf_reg[895] ),
    .S0(_1525_),
    .S1(_1255_),
    .X(_1590_));
 sky130_fd_sc_hd__mux4_1 _3941_ (.A0(\rf_reg[927] ),
    .A1(\rf_reg[959] ),
    .A2(\rf_reg[991] ),
    .A3(\rf_reg[1023] ),
    .S0(_1475_),
    .S1(_1541_),
    .X(_1591_));
 sky130_fd_sc_hd__mux4_1 _3942_ (.A0(_1588_),
    .A1(_1589_),
    .A2(_1590_),
    .A3(_1591_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1592_));
 sky130_fd_sc_hd__mux2_4 _3943_ (.A0(_1587_),
    .A1(_1592_),
    .S(_1546_),
    .X(net71));
 sky130_fd_sc_hd__mux2_1 _3944_ (.A0(\rf_reg[35] ),
    .A1(\rf_reg[99] ),
    .S(_1253_),
    .X(_1593_));
 sky130_fd_sc_hd__a22o_1 _3945_ (.A1(\rf_reg[67] ),
    .A2(_1529_),
    .B1(_1593_),
    .B2(_1531_),
    .X(_1594_));
 sky130_fd_sc_hd__mux4_2 _3946_ (.A0(\rf_reg[131] ),
    .A1(\rf_reg[163] ),
    .A2(\rf_reg[195] ),
    .A3(\rf_reg[227] ),
    .S0(_1244_),
    .S1(_1504_),
    .X(_1595_));
 sky130_fd_sc_hd__mux4_1 _3947_ (.A0(\rf_reg[515] ),
    .A1(\rf_reg[547] ),
    .A2(\rf_reg[579] ),
    .A3(\rf_reg[611] ),
    .S0(_1493_),
    .S1(_1562_),
    .X(_1596_));
 sky130_fd_sc_hd__mux4_1 _3948_ (.A0(\rf_reg[643] ),
    .A1(\rf_reg[675] ),
    .A2(\rf_reg[707] ),
    .A3(\rf_reg[739] ),
    .S0(_1267_),
    .S1(_1507_),
    .X(_1597_));
 sky130_fd_sc_hd__mux4_1 _3949_ (.A0(_1594_),
    .A1(_1595_),
    .A2(_1596_),
    .A3(_1597_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1598_));
 sky130_fd_sc_hd__mux4_1 _3950_ (.A0(\rf_reg[259] ),
    .A1(\rf_reg[291] ),
    .A2(\rf_reg[323] ),
    .A3(\rf_reg[355] ),
    .S0(_1553_),
    .S1(_1484_),
    .X(_1599_));
 sky130_fd_sc_hd__mux4_1 _3951_ (.A0(\rf_reg[387] ),
    .A1(\rf_reg[419] ),
    .A2(\rf_reg[451] ),
    .A3(\rf_reg[483] ),
    .S0(_1249_),
    .S1(_1538_),
    .X(_1600_));
 sky130_fd_sc_hd__mux4_1 _3952_ (.A0(\rf_reg[771] ),
    .A1(\rf_reg[803] ),
    .A2(\rf_reg[835] ),
    .A3(\rf_reg[867] ),
    .S0(_1525_),
    .S1(_1255_),
    .X(_1601_));
 sky130_fd_sc_hd__mux4_1 _3953_ (.A0(\rf_reg[899] ),
    .A1(\rf_reg[931] ),
    .A2(\rf_reg[963] ),
    .A3(\rf_reg[995] ),
    .S0(_1258_),
    .S1(_1541_),
    .X(_1602_));
 sky130_fd_sc_hd__mux4_1 _3954_ (.A0(_1599_),
    .A1(_1600_),
    .A2(_1601_),
    .A3(_1602_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(_1598_),
    .A1(_1603_),
    .S(_1546_),
    .X(net72));
 sky130_fd_sc_hd__mux2_1 _3956_ (.A0(\rf_reg[36] ),
    .A1(\rf_reg[100] ),
    .S(_1253_),
    .X(_1604_));
 sky130_fd_sc_hd__a22o_1 _3957_ (.A1(\rf_reg[68] ),
    .A2(_1529_),
    .B1(_1604_),
    .B2(_1531_),
    .X(_1605_));
 sky130_fd_sc_hd__mux4_4 _3958_ (.A0(\rf_reg[132] ),
    .A1(\rf_reg[164] ),
    .A2(\rf_reg[196] ),
    .A3(\rf_reg[228] ),
    .S0(_1244_),
    .S1(_1504_),
    .X(_1606_));
 sky130_fd_sc_hd__mux4_1 _3959_ (.A0(\rf_reg[516] ),
    .A1(\rf_reg[548] ),
    .A2(\rf_reg[580] ),
    .A3(\rf_reg[612] ),
    .S0(_1493_),
    .S1(_1562_),
    .X(_1607_));
 sky130_fd_sc_hd__mux4_1 _3960_ (.A0(\rf_reg[644] ),
    .A1(\rf_reg[676] ),
    .A2(\rf_reg[708] ),
    .A3(\rf_reg[740] ),
    .S0(_1267_),
    .S1(_1507_),
    .X(_1608_));
 sky130_fd_sc_hd__mux4_1 _3961_ (.A0(_1605_),
    .A1(_1606_),
    .A2(_1607_),
    .A3(_1608_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1609_));
 sky130_fd_sc_hd__mux4_1 _3962_ (.A0(\rf_reg[260] ),
    .A1(\rf_reg[292] ),
    .A2(\rf_reg[324] ),
    .A3(\rf_reg[356] ),
    .S0(_1553_),
    .S1(_1274_),
    .X(_1610_));
 sky130_fd_sc_hd__mux4_1 _3963_ (.A0(\rf_reg[388] ),
    .A1(\rf_reg[420] ),
    .A2(\rf_reg[452] ),
    .A3(\rf_reg[484] ),
    .S0(_1249_),
    .S1(_1538_),
    .X(_1611_));
 sky130_fd_sc_hd__mux4_1 _3964_ (.A0(\rf_reg[772] ),
    .A1(\rf_reg[804] ),
    .A2(\rf_reg[836] ),
    .A3(\rf_reg[868] ),
    .S0(_1525_),
    .S1(_1255_),
    .X(_1612_));
 sky130_fd_sc_hd__mux4_1 _3965_ (.A0(\rf_reg[900] ),
    .A1(\rf_reg[932] ),
    .A2(\rf_reg[964] ),
    .A3(\rf_reg[996] ),
    .S0(_1258_),
    .S1(_1541_),
    .X(_1613_));
 sky130_fd_sc_hd__mux4_1 _3966_ (.A0(_1610_),
    .A1(_1611_),
    .A2(_1612_),
    .A3(_1613_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_2 _3967_ (.A0(_1609_),
    .A1(_1614_),
    .S(_1546_),
    .X(net73));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(\rf_reg[37] ),
    .A1(\rf_reg[101] ),
    .S(_1253_),
    .X(_1615_));
 sky130_fd_sc_hd__a22o_1 _3969_ (.A1(\rf_reg[69] ),
    .A2(_1529_),
    .B1(_1615_),
    .B2(_1531_),
    .X(_1616_));
 sky130_fd_sc_hd__mux4_1 _3970_ (.A0(\rf_reg[133] ),
    .A1(\rf_reg[165] ),
    .A2(\rf_reg[197] ),
    .A3(\rf_reg[229] ),
    .S0(_1244_),
    .S1(_1504_),
    .X(_1617_));
 sky130_fd_sc_hd__mux4_1 _3971_ (.A0(\rf_reg[517] ),
    .A1(\rf_reg[549] ),
    .A2(\rf_reg[581] ),
    .A3(\rf_reg[613] ),
    .S0(_1270_),
    .S1(_1562_),
    .X(_1618_));
 sky130_fd_sc_hd__mux4_1 _3972_ (.A0(\rf_reg[645] ),
    .A1(\rf_reg[677] ),
    .A2(\rf_reg[709] ),
    .A3(\rf_reg[741] ),
    .S0(_1267_),
    .S1(_1507_),
    .X(_1619_));
 sky130_fd_sc_hd__mux4_1 _3973_ (.A0(_1616_),
    .A1(_1617_),
    .A2(_1618_),
    .A3(_1619_),
    .S0(_1509_),
    .S1(_1510_),
    .X(_1620_));
 sky130_fd_sc_hd__mux4_1 _3974_ (.A0(\rf_reg[261] ),
    .A1(\rf_reg[293] ),
    .A2(\rf_reg[325] ),
    .A3(\rf_reg[357] ),
    .S0(_1553_),
    .S1(_1274_),
    .X(_1621_));
 sky130_fd_sc_hd__mux4_1 _3975_ (.A0(\rf_reg[389] ),
    .A1(\rf_reg[421] ),
    .A2(\rf_reg[453] ),
    .A3(\rf_reg[485] ),
    .S0(_1249_),
    .S1(_1538_),
    .X(_1622_));
 sky130_fd_sc_hd__mux4_1 _3976_ (.A0(\rf_reg[773] ),
    .A1(\rf_reg[805] ),
    .A2(\rf_reg[837] ),
    .A3(\rf_reg[869] ),
    .S0(_1525_),
    .S1(_1255_),
    .X(_1623_));
 sky130_fd_sc_hd__mux4_1 _3977_ (.A0(\rf_reg[901] ),
    .A1(\rf_reg[933] ),
    .A2(\rf_reg[965] ),
    .A3(\rf_reg[997] ),
    .S0(_1258_),
    .S1(_1541_),
    .X(_1624_));
 sky130_fd_sc_hd__mux4_1 _3978_ (.A0(_1621_),
    .A1(_1622_),
    .A2(_1623_),
    .A3(_1624_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1625_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(_1620_),
    .A1(_1625_),
    .S(_1546_),
    .X(net74));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(\rf_reg[38] ),
    .A1(\rf_reg[102] ),
    .S(_1253_),
    .X(_1626_));
 sky130_fd_sc_hd__a22o_1 _3981_ (.A1(\rf_reg[70] ),
    .A2(_1529_),
    .B1(_1626_),
    .B2(_1531_),
    .X(_1627_));
 sky130_fd_sc_hd__mux4_1 _3982_ (.A0(\rf_reg[134] ),
    .A1(\rf_reg[166] ),
    .A2(\rf_reg[198] ),
    .A3(\rf_reg[230] ),
    .S0(_1244_),
    .S1(_1259_),
    .X(_1628_));
 sky130_fd_sc_hd__mux4_1 _3983_ (.A0(\rf_reg[518] ),
    .A1(\rf_reg[550] ),
    .A2(\rf_reg[582] ),
    .A3(\rf_reg[614] ),
    .S0(_1270_),
    .S1(_1562_),
    .X(_1629_));
 sky130_fd_sc_hd__mux4_1 _3984_ (.A0(\rf_reg[646] ),
    .A1(\rf_reg[678] ),
    .A2(\rf_reg[710] ),
    .A3(\rf_reg[742] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1630_));
 sky130_fd_sc_hd__mux4_1 _3985_ (.A0(_1627_),
    .A1(_1628_),
    .A2(_1629_),
    .A3(_1630_),
    .S0(_1262_),
    .S1(_1264_),
    .X(_1631_));
 sky130_fd_sc_hd__mux4_1 _3986_ (.A0(\rf_reg[262] ),
    .A1(\rf_reg[294] ),
    .A2(\rf_reg[326] ),
    .A3(\rf_reg[358] ),
    .S0(_1553_),
    .S1(_1274_),
    .X(_1632_));
 sky130_fd_sc_hd__mux4_1 _3987_ (.A0(\rf_reg[390] ),
    .A1(\rf_reg[422] ),
    .A2(\rf_reg[454] ),
    .A3(\rf_reg[486] ),
    .S0(_1249_),
    .S1(_1538_),
    .X(_1633_));
 sky130_fd_sc_hd__mux4_1 _3988_ (.A0(\rf_reg[774] ),
    .A1(\rf_reg[806] ),
    .A2(\rf_reg[838] ),
    .A3(\rf_reg[870] ),
    .S0(_1525_),
    .S1(_1255_),
    .X(_1634_));
 sky130_fd_sc_hd__mux4_1 _3989_ (.A0(\rf_reg[902] ),
    .A1(\rf_reg[934] ),
    .A2(\rf_reg[966] ),
    .A3(\rf_reg[998] ),
    .S0(_1258_),
    .S1(_1541_),
    .X(_1635_));
 sky130_fd_sc_hd__mux4_1 _3990_ (.A0(_1632_),
    .A1(_1633_),
    .A2(_1634_),
    .A3(_1635_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1636_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(_1631_),
    .A1(_1636_),
    .S(_1546_),
    .X(net75));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(\rf_reg[39] ),
    .A1(\rf_reg[103] ),
    .S(_1253_),
    .X(_1637_));
 sky130_fd_sc_hd__a22o_1 _3993_ (.A1(\rf_reg[71] ),
    .A2(_1529_),
    .B1(_1637_),
    .B2(_1531_),
    .X(_1638_));
 sky130_fd_sc_hd__mux4_1 _3994_ (.A0(\rf_reg[135] ),
    .A1(\rf_reg[167] ),
    .A2(\rf_reg[199] ),
    .A3(\rf_reg[231] ),
    .S0(_1244_),
    .S1(_1259_),
    .X(_1639_));
 sky130_fd_sc_hd__mux4_1 _3995_ (.A0(\rf_reg[519] ),
    .A1(\rf_reg[551] ),
    .A2(\rf_reg[583] ),
    .A3(\rf_reg[615] ),
    .S0(_1270_),
    .S1(_1562_),
    .X(_1640_));
 sky130_fd_sc_hd__mux4_1 _3996_ (.A0(\rf_reg[647] ),
    .A1(\rf_reg[679] ),
    .A2(\rf_reg[711] ),
    .A3(\rf_reg[743] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1641_));
 sky130_fd_sc_hd__mux4_1 _3997_ (.A0(_1638_),
    .A1(_1639_),
    .A2(_1640_),
    .A3(_1641_),
    .S0(_1262_),
    .S1(_1264_),
    .X(_1642_));
 sky130_fd_sc_hd__mux4_1 _3998_ (.A0(\rf_reg[263] ),
    .A1(\rf_reg[295] ),
    .A2(\rf_reg[327] ),
    .A3(\rf_reg[359] ),
    .S0(_1553_),
    .S1(_1274_),
    .X(_1643_));
 sky130_fd_sc_hd__mux4_1 _3999_ (.A0(\rf_reg[391] ),
    .A1(\rf_reg[423] ),
    .A2(\rf_reg[455] ),
    .A3(\rf_reg[487] ),
    .S0(_1249_),
    .S1(_1538_),
    .X(_1644_));
 sky130_fd_sc_hd__mux4_1 _4000_ (.A0(\rf_reg[775] ),
    .A1(\rf_reg[807] ),
    .A2(\rf_reg[839] ),
    .A3(\rf_reg[871] ),
    .S0(_1252_),
    .S1(_1255_),
    .X(_1645_));
 sky130_fd_sc_hd__mux4_1 _4001_ (.A0(\rf_reg[903] ),
    .A1(\rf_reg[935] ),
    .A2(\rf_reg[967] ),
    .A3(\rf_reg[999] ),
    .S0(_1258_),
    .S1(_1541_),
    .X(_1646_));
 sky130_fd_sc_hd__mux4_1 _4002_ (.A0(_1643_),
    .A1(_1644_),
    .A2(_1645_),
    .A3(_1646_),
    .S0(_1543_),
    .S1(_1544_),
    .X(_1647_));
 sky130_fd_sc_hd__mux2_1 _4003_ (.A0(_1642_),
    .A1(_1647_),
    .S(_1546_),
    .X(net76));
 sky130_fd_sc_hd__mux2_1 _4004_ (.A0(\rf_reg[40] ),
    .A1(\rf_reg[104] ),
    .S(_1253_),
    .X(_1648_));
 sky130_fd_sc_hd__a22o_1 _4005_ (.A1(\rf_reg[72] ),
    .A2(_1240_),
    .B1(_1648_),
    .B2(_1245_),
    .X(_1649_));
 sky130_fd_sc_hd__mux4_1 _4006_ (.A0(\rf_reg[136] ),
    .A1(\rf_reg[168] ),
    .A2(\rf_reg[200] ),
    .A3(\rf_reg[232] ),
    .S0(_1244_),
    .S1(_1259_),
    .X(_1650_));
 sky130_fd_sc_hd__mux4_1 _4007_ (.A0(\rf_reg[520] ),
    .A1(\rf_reg[552] ),
    .A2(\rf_reg[584] ),
    .A3(\rf_reg[616] ),
    .S0(_1270_),
    .S1(_1562_),
    .X(_1651_));
 sky130_fd_sc_hd__mux4_1 _4008_ (.A0(\rf_reg[648] ),
    .A1(\rf_reg[680] ),
    .A2(\rf_reg[712] ),
    .A3(\rf_reg[744] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1652_));
 sky130_fd_sc_hd__mux4_1 _4009_ (.A0(_1649_),
    .A1(_1650_),
    .A2(_1651_),
    .A3(_1652_),
    .S0(_1262_),
    .S1(_1264_),
    .X(_1653_));
 sky130_fd_sc_hd__mux4_1 _4010_ (.A0(\rf_reg[264] ),
    .A1(\rf_reg[296] ),
    .A2(\rf_reg[328] ),
    .A3(\rf_reg[360] ),
    .S0(_1553_),
    .S1(_1274_),
    .X(_1654_));
 sky130_fd_sc_hd__mux4_1 _4011_ (.A0(\rf_reg[392] ),
    .A1(\rf_reg[424] ),
    .A2(\rf_reg[456] ),
    .A3(\rf_reg[488] ),
    .S0(_1249_),
    .S1(_1250_),
    .X(_1655_));
 sky130_fd_sc_hd__mux4_1 _4012_ (.A0(\rf_reg[776] ),
    .A1(\rf_reg[808] ),
    .A2(\rf_reg[840] ),
    .A3(\rf_reg[872] ),
    .S0(_1252_),
    .S1(_1255_),
    .X(_1656_));
 sky130_fd_sc_hd__mux4_1 _4013_ (.A0(\rf_reg[904] ),
    .A1(\rf_reg[936] ),
    .A2(\rf_reg[968] ),
    .A3(\rf_reg[1000] ),
    .S0(_1258_),
    .S1(_1260_),
    .X(_1657_));
 sky130_fd_sc_hd__mux4_1 _4014_ (.A0(_1654_),
    .A1(_1655_),
    .A2(_1656_),
    .A3(_1657_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1658_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(_1653_),
    .A1(_1658_),
    .S(_1281_),
    .X(net77));
 sky130_fd_sc_hd__mux2_1 _4016_ (.A0(\rf_reg[41] ),
    .A1(\rf_reg[105] ),
    .S(_1253_),
    .X(_1659_));
 sky130_fd_sc_hd__a22o_1 _4017_ (.A1(\rf_reg[73] ),
    .A2(_1240_),
    .B1(_1659_),
    .B2(_1245_),
    .X(_1660_));
 sky130_fd_sc_hd__mux4_1 _4018_ (.A0(\rf_reg[137] ),
    .A1(\rf_reg[169] ),
    .A2(\rf_reg[201] ),
    .A3(\rf_reg[233] ),
    .S0(_1244_),
    .S1(_1259_),
    .X(_1661_));
 sky130_fd_sc_hd__mux4_1 _4019_ (.A0(\rf_reg[521] ),
    .A1(\rf_reg[553] ),
    .A2(\rf_reg[585] ),
    .A3(\rf_reg[617] ),
    .S0(_1270_),
    .S1(_1562_),
    .X(_1662_));
 sky130_fd_sc_hd__mux4_1 _4020_ (.A0(\rf_reg[649] ),
    .A1(\rf_reg[681] ),
    .A2(\rf_reg[713] ),
    .A3(\rf_reg[745] ),
    .S0(_1267_),
    .S1(_1268_),
    .X(_1663_));
 sky130_fd_sc_hd__mux4_1 _4021_ (.A0(_1660_),
    .A1(_1661_),
    .A2(_1662_),
    .A3(_1663_),
    .S0(_1262_),
    .S1(_1264_),
    .X(_1664_));
 sky130_fd_sc_hd__mux4_1 _4022_ (.A0(\rf_reg[265] ),
    .A1(\rf_reg[297] ),
    .A2(\rf_reg[329] ),
    .A3(\rf_reg[361] ),
    .S0(_1273_),
    .S1(_1274_),
    .X(_1665_));
 sky130_fd_sc_hd__mux4_1 _4023_ (.A0(\rf_reg[393] ),
    .A1(\rf_reg[425] ),
    .A2(\rf_reg[457] ),
    .A3(\rf_reg[489] ),
    .S0(_1249_),
    .S1(_1250_),
    .X(_1666_));
 sky130_fd_sc_hd__mux4_1 _4024_ (.A0(\rf_reg[777] ),
    .A1(\rf_reg[809] ),
    .A2(\rf_reg[841] ),
    .A3(\rf_reg[873] ),
    .S0(_1252_),
    .S1(_1255_),
    .X(_1667_));
 sky130_fd_sc_hd__mux4_1 _4025_ (.A0(\rf_reg[905] ),
    .A1(\rf_reg[937] ),
    .A2(\rf_reg[969] ),
    .A3(\rf_reg[1001] ),
    .S0(_1258_),
    .S1(_1260_),
    .X(_1668_));
 sky130_fd_sc_hd__mux4_1 _4026_ (.A0(_1665_),
    .A1(_1666_),
    .A2(_1667_),
    .A3(_1668_),
    .S0(_1263_),
    .S1(_1265_),
    .X(_1669_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(_1664_),
    .A1(_1669_),
    .S(_1281_),
    .X(net78));
 sky130_fd_sc_hd__buf_12 _4028_ (.A(raddr_b_i[4]),
    .X(_1670_));
 sky130_fd_sc_hd__buf_16 _4029_ (.A(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__clkbuf_16 _4030_ (.A(net1),
    .X(_1672_));
 sky130_fd_sc_hd__buf_8 _4031_ (.A(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__buf_12 _4032_ (.A(raddr_b_i[0]),
    .X(_1674_));
 sky130_fd_sc_hd__buf_16 _4033_ (.A(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__buf_8 _4034_ (.A(raddr_b_i[2]),
    .X(_1676_));
 sky130_fd_sc_hd__buf_12 _4035_ (.A(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__buf_16 _4036_ (.A(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__mux4_1 _4037_ (.A0(\rf_reg[256] ),
    .A1(\rf_reg[288] ),
    .A2(\rf_reg[384] ),
    .A3(\rf_reg[416] ),
    .S0(_1675_),
    .S1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__buf_16 _4038_ (.A(_1674_),
    .X(_1680_));
 sky130_fd_sc_hd__buf_16 _4039_ (.A(_1676_),
    .X(_1681_));
 sky130_fd_sc_hd__mux4_1 _4040_ (.A0(\rf_reg[320] ),
    .A1(\rf_reg[352] ),
    .A2(\rf_reg[448] ),
    .A3(\rf_reg[480] ),
    .S0(_1680_),
    .S1(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__buf_6 _4041_ (.A(raddr_b_i[1]),
    .X(_1683_));
 sky130_fd_sc_hd__buf_12 _4042_ (.A(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__buf_12 _4043_ (.A(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__mux2i_1 _4044_ (.A0(_1679_),
    .A1(_1682_),
    .S(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__and2_0 _4045_ (.A(_1673_),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__buf_12 _4046_ (.A(_1676_),
    .X(_1688_));
 sky130_fd_sc_hd__buf_8 _4047_ (.A(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__inv_6 _4048_ (.A(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__buf_8 _4049_ (.A(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(\rf_reg[64] ),
    .B(_1685_),
    .Y(_1692_));
 sky130_fd_sc_hd__mux2i_1 _4051_ (.A0(\rf_reg[32] ),
    .A1(\rf_reg[96] ),
    .S(_1684_),
    .Y(_1693_));
 sky130_fd_sc_hd__buf_12 _4052_ (.A(_1674_),
    .X(_1694_));
 sky130_fd_sc_hd__buf_16 _4053_ (.A(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__buf_8 _4054_ (.A(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__buf_8 _4055_ (.A(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__mux2i_1 _4056_ (.A0(_1692_),
    .A1(_1693_),
    .S(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_8 _4057_ (.A(_1684_),
    .B(_1688_),
    .Y(_1699_));
 sky130_fd_sc_hd__buf_8 _4058_ (.A(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__buf_8 _4059_ (.A(_1694_),
    .X(_1701_));
 sky130_fd_sc_hd__buf_8 _4060_ (.A(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__mux2i_1 _4061_ (.A0(\rf_reg[192] ),
    .A1(\rf_reg[224] ),
    .S(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__nand2b_4 _4062_ (.A_N(_1684_),
    .B(_1677_),
    .Y(_1704_));
 sky130_fd_sc_hd__buf_8 _4063_ (.A(_1696_),
    .X(_1705_));
 sky130_fd_sc_hd__mux2i_1 _4064_ (.A0(\rf_reg[128] ),
    .A1(\rf_reg[160] ),
    .S(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__o22ai_2 _4065_ (.A1(_1700_),
    .A2(_1703_),
    .B1(_1704_),
    .B2(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__buf_8 _4066_ (.A(_1672_),
    .X(_1708_));
 sky130_fd_sc_hd__a211oi_2 _4067_ (.A1(_1691_),
    .A2(_1698_),
    .B1(_1707_),
    .C1(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__buf_8 _4068_ (.A(_1694_),
    .X(_1710_));
 sky130_fd_sc_hd__buf_6 _4069_ (.A(_1677_),
    .X(_1711_));
 sky130_fd_sc_hd__mux4_1 _4070_ (.A0(\rf_reg[768] ),
    .A1(\rf_reg[800] ),
    .A2(\rf_reg[896] ),
    .A3(\rf_reg[928] ),
    .S0(_1710_),
    .S1(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__nor2b_1 _4071_ (.A(_1683_),
    .B_N(net1),
    .Y(_1713_));
 sky130_fd_sc_hd__buf_4 _4072_ (.A(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__buf_16 _4073_ (.A(_1694_),
    .X(_1715_));
 sky130_fd_sc_hd__buf_8 _4074_ (.A(_1688_),
    .X(_1716_));
 sky130_fd_sc_hd__mux4_1 _4075_ (.A0(\rf_reg[512] ),
    .A1(\rf_reg[544] ),
    .A2(\rf_reg[640] ),
    .A3(\rf_reg[672] ),
    .S0(_1715_),
    .S1(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__nor2_8 _4076_ (.A(_1684_),
    .B(net1),
    .Y(_1718_));
 sky130_fd_sc_hd__buf_6 _4077_ (.A(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__a22o_1 _4078_ (.A1(_1712_),
    .A2(_1714_),
    .B1(_1717_),
    .B2(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__buf_16 _4079_ (.A(_1694_),
    .X(_1721_));
 sky130_fd_sc_hd__mux4_1 _4080_ (.A0(\rf_reg[832] ),
    .A1(\rf_reg[864] ),
    .A2(\rf_reg[960] ),
    .A3(\rf_reg[992] ),
    .S0(_1721_),
    .S1(_1711_),
    .X(_1722_));
 sky130_fd_sc_hd__and2_0 _4081_ (.A(_1683_),
    .B(net1),
    .X(_1723_));
 sky130_fd_sc_hd__buf_4 _4082_ (.A(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__mux4_1 _4083_ (.A0(\rf_reg[576] ),
    .A1(\rf_reg[608] ),
    .A2(\rf_reg[704] ),
    .A3(\rf_reg[736] ),
    .S0(_1701_),
    .S1(_1689_),
    .X(_1725_));
 sky130_fd_sc_hd__nor2b_1 _4084_ (.A(net1),
    .B_N(_1683_),
    .Y(_1726_));
 sky130_fd_sc_hd__buf_6 _4085_ (.A(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__buf_6 _4086_ (.A(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__a22o_1 _4087_ (.A1(_1722_),
    .A2(_1724_),
    .B1(_1725_),
    .B2(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__buf_6 _4088_ (.A(_1670_),
    .X(_1730_));
 sky130_fd_sc_hd__o21ai_1 _4089_ (.A1(_1720_),
    .A2(_1729_),
    .B1(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__o31ai_4 _4090_ (.A1(_1671_),
    .A2(_1687_),
    .A3(_1709_),
    .B1(_1731_),
    .Y(net79));
 sky130_fd_sc_hd__buf_16 _4091_ (.A(_1677_),
    .X(_1732_));
 sky130_fd_sc_hd__mux4_1 _4092_ (.A0(\rf_reg[266] ),
    .A1(\rf_reg[298] ),
    .A2(\rf_reg[394] ),
    .A3(\rf_reg[426] ),
    .S0(_1675_),
    .S1(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__mux4_1 _4093_ (.A0(\rf_reg[330] ),
    .A1(\rf_reg[362] ),
    .A2(\rf_reg[458] ),
    .A3(\rf_reg[490] ),
    .S0(_1680_),
    .S1(_1681_),
    .X(_1734_));
 sky130_fd_sc_hd__mux2i_1 _4094_ (.A0(_1733_),
    .A1(_1734_),
    .S(_1685_),
    .Y(_1735_));
 sky130_fd_sc_hd__and2_0 _4095_ (.A(_1673_),
    .B(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(\rf_reg[42] ),
    .A1(\rf_reg[106] ),
    .S(_1683_),
    .X(_1737_));
 sky130_fd_sc_hd__nor2b_4 _4097_ (.A(_1675_),
    .B_N(_1683_),
    .Y(_1738_));
 sky130_fd_sc_hd__buf_8 _4098_ (.A(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__a22o_1 _4099_ (.A1(_1705_),
    .A2(_1737_),
    .B1(_1739_),
    .B2(\rf_reg[74] ),
    .X(_1740_));
 sky130_fd_sc_hd__mux2i_1 _4100_ (.A0(\rf_reg[202] ),
    .A1(\rf_reg[234] ),
    .S(_1702_),
    .Y(_1741_));
 sky130_fd_sc_hd__mux2i_1 _4101_ (.A0(\rf_reg[138] ),
    .A1(\rf_reg[170] ),
    .S(_1705_),
    .Y(_1742_));
 sky130_fd_sc_hd__buf_8 _4102_ (.A(_1704_),
    .X(_1743_));
 sky130_fd_sc_hd__o22ai_1 _4103_ (.A1(_1700_),
    .A2(_1741_),
    .B1(_1742_),
    .B2(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__a211oi_1 _4104_ (.A1(_1691_),
    .A2(_1740_),
    .B1(_1744_),
    .C1(_1708_),
    .Y(_1745_));
 sky130_fd_sc_hd__buf_6 _4105_ (.A(_1714_),
    .X(_1746_));
 sky130_fd_sc_hd__buf_16 _4106_ (.A(_1677_),
    .X(_1747_));
 sky130_fd_sc_hd__mux4_1 _4107_ (.A0(\rf_reg[778] ),
    .A1(\rf_reg[810] ),
    .A2(\rf_reg[906] ),
    .A3(\rf_reg[938] ),
    .S0(_1695_),
    .S1(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__mux4_1 _4108_ (.A0(\rf_reg[522] ),
    .A1(\rf_reg[554] ),
    .A2(\rf_reg[650] ),
    .A3(\rf_reg[682] ),
    .S0(_1715_),
    .S1(_1716_),
    .X(_1749_));
 sky130_fd_sc_hd__a22o_1 _4109_ (.A1(_1746_),
    .A2(_1748_),
    .B1(_1749_),
    .B2(_1719_),
    .X(_1750_));
 sky130_fd_sc_hd__buf_6 _4110_ (.A(_1724_),
    .X(_1751_));
 sky130_fd_sc_hd__mux4_1 _4111_ (.A0(\rf_reg[842] ),
    .A1(\rf_reg[874] ),
    .A2(\rf_reg[970] ),
    .A3(\rf_reg[1002] ),
    .S0(_1710_),
    .S1(_1711_),
    .X(_1752_));
 sky130_fd_sc_hd__mux4_1 _4112_ (.A0(\rf_reg[586] ),
    .A1(\rf_reg[618] ),
    .A2(\rf_reg[714] ),
    .A3(\rf_reg[746] ),
    .S0(_1701_),
    .S1(_1689_),
    .X(_1753_));
 sky130_fd_sc_hd__a22o_1 _4113_ (.A1(_1751_),
    .A2(_1752_),
    .B1(_1753_),
    .B2(_1728_),
    .X(_1754_));
 sky130_fd_sc_hd__o21ai_2 _4114_ (.A1(_1750_),
    .A2(_1754_),
    .B1(_1730_),
    .Y(_1755_));
 sky130_fd_sc_hd__o31ai_2 _4115_ (.A1(_1671_),
    .A2(_1736_),
    .A3(_1745_),
    .B1(_1755_),
    .Y(net80));
 sky130_fd_sc_hd__mux4_1 _4116_ (.A0(\rf_reg[267] ),
    .A1(\rf_reg[299] ),
    .A2(\rf_reg[395] ),
    .A3(\rf_reg[427] ),
    .S0(_1675_),
    .S1(_1732_),
    .X(_1756_));
 sky130_fd_sc_hd__mux4_1 _4117_ (.A0(\rf_reg[331] ),
    .A1(\rf_reg[363] ),
    .A2(\rf_reg[459] ),
    .A3(\rf_reg[491] ),
    .S0(_1680_),
    .S1(_1681_),
    .X(_1757_));
 sky130_fd_sc_hd__mux2i_1 _4118_ (.A0(_1756_),
    .A1(_1757_),
    .S(_1685_),
    .Y(_1758_));
 sky130_fd_sc_hd__and2_0 _4119_ (.A(_1673_),
    .B(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__buf_8 _4120_ (.A(_1683_),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_1 _4121_ (.A0(\rf_reg[43] ),
    .A1(\rf_reg[107] ),
    .S(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__a22o_1 _4122_ (.A1(\rf_reg[75] ),
    .A2(_1739_),
    .B1(_1761_),
    .B2(_1697_),
    .X(_1762_));
 sky130_fd_sc_hd__mux2i_1 _4123_ (.A0(\rf_reg[203] ),
    .A1(\rf_reg[235] ),
    .S(_1702_),
    .Y(_1763_));
 sky130_fd_sc_hd__mux2i_1 _4124_ (.A0(\rf_reg[139] ),
    .A1(\rf_reg[171] ),
    .S(_1705_),
    .Y(_1764_));
 sky130_fd_sc_hd__o22ai_1 _4125_ (.A1(_1700_),
    .A2(_1763_),
    .B1(_1764_),
    .B2(_1743_),
    .Y(_1765_));
 sky130_fd_sc_hd__a211oi_1 _4126_ (.A1(_1691_),
    .A2(_1762_),
    .B1(_1765_),
    .C1(_1708_),
    .Y(_1766_));
 sky130_fd_sc_hd__mux4_1 _4127_ (.A0(\rf_reg[779] ),
    .A1(\rf_reg[811] ),
    .A2(\rf_reg[907] ),
    .A3(\rf_reg[939] ),
    .S0(_1695_),
    .S1(_1747_),
    .X(_1767_));
 sky130_fd_sc_hd__mux4_1 _4128_ (.A0(\rf_reg[523] ),
    .A1(\rf_reg[555] ),
    .A2(\rf_reg[651] ),
    .A3(\rf_reg[683] ),
    .S0(_1715_),
    .S1(_1716_),
    .X(_1768_));
 sky130_fd_sc_hd__a22o_1 _4129_ (.A1(_1746_),
    .A2(_1767_),
    .B1(_1768_),
    .B2(_1719_),
    .X(_1769_));
 sky130_fd_sc_hd__mux4_1 _4130_ (.A0(\rf_reg[843] ),
    .A1(\rf_reg[875] ),
    .A2(\rf_reg[971] ),
    .A3(\rf_reg[1003] ),
    .S0(_1710_),
    .S1(_1711_),
    .X(_1770_));
 sky130_fd_sc_hd__mux4_1 _4131_ (.A0(\rf_reg[587] ),
    .A1(\rf_reg[619] ),
    .A2(\rf_reg[715] ),
    .A3(\rf_reg[747] ),
    .S0(_1701_),
    .S1(_1689_),
    .X(_1771_));
 sky130_fd_sc_hd__a22o_1 _4132_ (.A1(_1751_),
    .A2(_1770_),
    .B1(_1771_),
    .B2(_1728_),
    .X(_1772_));
 sky130_fd_sc_hd__o21ai_1 _4133_ (.A1(_1769_),
    .A2(_1772_),
    .B1(_1730_),
    .Y(_1773_));
 sky130_fd_sc_hd__o31ai_1 _4134_ (.A1(_1671_),
    .A2(_1759_),
    .A3(_1766_),
    .B1(_1773_),
    .Y(net81));
 sky130_fd_sc_hd__mux4_1 _4135_ (.A0(\rf_reg[268] ),
    .A1(\rf_reg[300] ),
    .A2(\rf_reg[396] ),
    .A3(\rf_reg[428] ),
    .S0(_1675_),
    .S1(_1732_),
    .X(_1774_));
 sky130_fd_sc_hd__buf_12 _4136_ (.A(_1674_),
    .X(_1775_));
 sky130_fd_sc_hd__mux4_1 _4137_ (.A0(\rf_reg[332] ),
    .A1(\rf_reg[364] ),
    .A2(\rf_reg[460] ),
    .A3(\rf_reg[492] ),
    .S0(_1775_),
    .S1(_1681_),
    .X(_1776_));
 sky130_fd_sc_hd__mux2i_1 _4138_ (.A0(_1774_),
    .A1(_1776_),
    .S(_1685_),
    .Y(_1777_));
 sky130_fd_sc_hd__and2_0 _4139_ (.A(_1673_),
    .B(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__mux2_1 _4140_ (.A0(\rf_reg[44] ),
    .A1(\rf_reg[108] ),
    .S(_1760_),
    .X(_1779_));
 sky130_fd_sc_hd__a22o_1 _4141_ (.A1(\rf_reg[76] ),
    .A2(_1739_),
    .B1(_1779_),
    .B2(_1697_),
    .X(_1780_));
 sky130_fd_sc_hd__mux2i_1 _4142_ (.A0(\rf_reg[204] ),
    .A1(\rf_reg[236] ),
    .S(_1702_),
    .Y(_1781_));
 sky130_fd_sc_hd__mux2i_1 _4143_ (.A0(\rf_reg[140] ),
    .A1(\rf_reg[172] ),
    .S(_1705_),
    .Y(_1782_));
 sky130_fd_sc_hd__o22ai_1 _4144_ (.A1(_1700_),
    .A2(_1781_),
    .B1(_1782_),
    .B2(_1743_),
    .Y(_1783_));
 sky130_fd_sc_hd__a211oi_1 _4145_ (.A1(_1691_),
    .A2(_1780_),
    .B1(_1783_),
    .C1(_1708_),
    .Y(_1784_));
 sky130_fd_sc_hd__buf_8 _4146_ (.A(_1677_),
    .X(_1785_));
 sky130_fd_sc_hd__mux4_1 _4147_ (.A0(\rf_reg[780] ),
    .A1(\rf_reg[812] ),
    .A2(\rf_reg[908] ),
    .A3(\rf_reg[940] ),
    .S0(_1695_),
    .S1(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__buf_8 _4148_ (.A(_1694_),
    .X(_1787_));
 sky130_fd_sc_hd__mux4_1 _4149_ (.A0(\rf_reg[524] ),
    .A1(\rf_reg[556] ),
    .A2(\rf_reg[652] ),
    .A3(\rf_reg[684] ),
    .S0(_1787_),
    .S1(_1716_),
    .X(_1788_));
 sky130_fd_sc_hd__a22o_1 _4150_ (.A1(_1746_),
    .A2(_1786_),
    .B1(_1788_),
    .B2(_1719_),
    .X(_1789_));
 sky130_fd_sc_hd__mux4_1 _4151_ (.A0(\rf_reg[844] ),
    .A1(\rf_reg[876] ),
    .A2(\rf_reg[972] ),
    .A3(\rf_reg[1004] ),
    .S0(_1710_),
    .S1(_1711_),
    .X(_1790_));
 sky130_fd_sc_hd__mux4_1 _4152_ (.A0(\rf_reg[588] ),
    .A1(\rf_reg[620] ),
    .A2(\rf_reg[716] ),
    .A3(\rf_reg[748] ),
    .S0(_1701_),
    .S1(_1689_),
    .X(_1791_));
 sky130_fd_sc_hd__a22o_1 _4153_ (.A1(_1751_),
    .A2(_1790_),
    .B1(_1791_),
    .B2(_1728_),
    .X(_1792_));
 sky130_fd_sc_hd__o21ai_1 _4154_ (.A1(_1789_),
    .A2(_1792_),
    .B1(_1730_),
    .Y(_1793_));
 sky130_fd_sc_hd__o31ai_1 _4155_ (.A1(_1671_),
    .A2(_1778_),
    .A3(_1784_),
    .B1(_1793_),
    .Y(net82));
 sky130_fd_sc_hd__mux4_1 _4156_ (.A0(\rf_reg[269] ),
    .A1(\rf_reg[301] ),
    .A2(\rf_reg[397] ),
    .A3(\rf_reg[429] ),
    .S0(_1675_),
    .S1(_1732_),
    .X(_1794_));
 sky130_fd_sc_hd__mux4_1 _4157_ (.A0(\rf_reg[333] ),
    .A1(\rf_reg[365] ),
    .A2(\rf_reg[461] ),
    .A3(\rf_reg[493] ),
    .S0(_1775_),
    .S1(_1681_),
    .X(_1795_));
 sky130_fd_sc_hd__mux2i_1 _4158_ (.A0(_1794_),
    .A1(_1795_),
    .S(_1685_),
    .Y(_1796_));
 sky130_fd_sc_hd__and2_0 _4159_ (.A(_1673_),
    .B(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__mux2_1 _4160_ (.A0(\rf_reg[45] ),
    .A1(\rf_reg[109] ),
    .S(_1760_),
    .X(_1798_));
 sky130_fd_sc_hd__a22o_1 _4161_ (.A1(\rf_reg[77] ),
    .A2(_1739_),
    .B1(_1798_),
    .B2(_1697_),
    .X(_1799_));
 sky130_fd_sc_hd__mux2i_1 _4162_ (.A0(\rf_reg[205] ),
    .A1(\rf_reg[237] ),
    .S(_1702_),
    .Y(_1800_));
 sky130_fd_sc_hd__mux2i_1 _4163_ (.A0(\rf_reg[141] ),
    .A1(\rf_reg[173] ),
    .S(_1705_),
    .Y(_1801_));
 sky130_fd_sc_hd__o22ai_1 _4164_ (.A1(_1700_),
    .A2(_1800_),
    .B1(_1801_),
    .B2(_1743_),
    .Y(_1802_));
 sky130_fd_sc_hd__a211oi_1 _4165_ (.A1(_1691_),
    .A2(_1799_),
    .B1(_1802_),
    .C1(_1708_),
    .Y(_1803_));
 sky130_fd_sc_hd__mux4_1 _4166_ (.A0(\rf_reg[781] ),
    .A1(\rf_reg[813] ),
    .A2(\rf_reg[909] ),
    .A3(\rf_reg[941] ),
    .S0(_1695_),
    .S1(_1785_),
    .X(_1804_));
 sky130_fd_sc_hd__mux4_1 _4167_ (.A0(\rf_reg[525] ),
    .A1(\rf_reg[557] ),
    .A2(\rf_reg[653] ),
    .A3(\rf_reg[685] ),
    .S0(_1787_),
    .S1(_1716_),
    .X(_1805_));
 sky130_fd_sc_hd__a22o_1 _4168_ (.A1(_1746_),
    .A2(_1804_),
    .B1(_1805_),
    .B2(_1719_),
    .X(_1806_));
 sky130_fd_sc_hd__buf_8 _4169_ (.A(_1677_),
    .X(_1807_));
 sky130_fd_sc_hd__mux4_1 _4170_ (.A0(\rf_reg[845] ),
    .A1(\rf_reg[877] ),
    .A2(\rf_reg[973] ),
    .A3(\rf_reg[1005] ),
    .S0(_1710_),
    .S1(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__mux4_1 _4171_ (.A0(\rf_reg[589] ),
    .A1(\rf_reg[621] ),
    .A2(\rf_reg[717] ),
    .A3(\rf_reg[749] ),
    .S0(_1701_),
    .S1(_1689_),
    .X(_1809_));
 sky130_fd_sc_hd__a22o_1 _4172_ (.A1(_1751_),
    .A2(_1808_),
    .B1(_1809_),
    .B2(_1728_),
    .X(_1810_));
 sky130_fd_sc_hd__o21ai_1 _4173_ (.A1(_1806_),
    .A2(_1810_),
    .B1(_1730_),
    .Y(_1811_));
 sky130_fd_sc_hd__o31ai_1 _4174_ (.A1(_1671_),
    .A2(_1797_),
    .A3(_1803_),
    .B1(_1811_),
    .Y(net83));
 sky130_fd_sc_hd__buf_16 _4175_ (.A(_1674_),
    .X(_1812_));
 sky130_fd_sc_hd__mux4_1 _4176_ (.A0(\rf_reg[270] ),
    .A1(\rf_reg[302] ),
    .A2(\rf_reg[398] ),
    .A3(\rf_reg[430] ),
    .S0(_1812_),
    .S1(_1732_),
    .X(_1813_));
 sky130_fd_sc_hd__mux4_1 _4177_ (.A0(\rf_reg[334] ),
    .A1(\rf_reg[366] ),
    .A2(\rf_reg[462] ),
    .A3(\rf_reg[494] ),
    .S0(_1775_),
    .S1(_1681_),
    .X(_1814_));
 sky130_fd_sc_hd__mux2i_1 _4178_ (.A0(_1813_),
    .A1(_1814_),
    .S(_1685_),
    .Y(_1815_));
 sky130_fd_sc_hd__and2_0 _4179_ (.A(_1673_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(\rf_reg[46] ),
    .A1(\rf_reg[110] ),
    .S(_1760_),
    .X(_1817_));
 sky130_fd_sc_hd__a22o_1 _4181_ (.A1(\rf_reg[78] ),
    .A2(_1739_),
    .B1(_1817_),
    .B2(_1697_),
    .X(_1818_));
 sky130_fd_sc_hd__mux2i_1 _4182_ (.A0(\rf_reg[206] ),
    .A1(\rf_reg[238] ),
    .S(_1702_),
    .Y(_1819_));
 sky130_fd_sc_hd__mux2i_1 _4183_ (.A0(\rf_reg[142] ),
    .A1(\rf_reg[174] ),
    .S(_1705_),
    .Y(_1820_));
 sky130_fd_sc_hd__o22ai_1 _4184_ (.A1(_1700_),
    .A2(_1819_),
    .B1(_1820_),
    .B2(_1743_),
    .Y(_1821_));
 sky130_fd_sc_hd__a211oi_1 _4185_ (.A1(_1691_),
    .A2(_1818_),
    .B1(_1821_),
    .C1(_1708_),
    .Y(_1822_));
 sky130_fd_sc_hd__mux4_1 _4186_ (.A0(\rf_reg[782] ),
    .A1(\rf_reg[814] ),
    .A2(\rf_reg[910] ),
    .A3(\rf_reg[942] ),
    .S0(_1695_),
    .S1(_1785_),
    .X(_1823_));
 sky130_fd_sc_hd__mux4_1 _4187_ (.A0(\rf_reg[526] ),
    .A1(\rf_reg[558] ),
    .A2(\rf_reg[654] ),
    .A3(\rf_reg[686] ),
    .S0(_1787_),
    .S1(_1716_),
    .X(_1824_));
 sky130_fd_sc_hd__a22o_1 _4188_ (.A1(_1746_),
    .A2(_1823_),
    .B1(_1824_),
    .B2(_1719_),
    .X(_1825_));
 sky130_fd_sc_hd__mux4_1 _4189_ (.A0(\rf_reg[846] ),
    .A1(\rf_reg[878] ),
    .A2(\rf_reg[974] ),
    .A3(\rf_reg[1006] ),
    .S0(_1710_),
    .S1(_1807_),
    .X(_1826_));
 sky130_fd_sc_hd__buf_16 _4190_ (.A(_1674_),
    .X(_1827_));
 sky130_fd_sc_hd__buf_8 _4191_ (.A(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__mux4_1 _4192_ (.A0(\rf_reg[590] ),
    .A1(\rf_reg[622] ),
    .A2(\rf_reg[718] ),
    .A3(\rf_reg[750] ),
    .S0(_1828_),
    .S1(_1689_),
    .X(_1829_));
 sky130_fd_sc_hd__a22o_1 _4193_ (.A1(_1751_),
    .A2(_1826_),
    .B1(_1829_),
    .B2(_1728_),
    .X(_1830_));
 sky130_fd_sc_hd__o21ai_1 _4194_ (.A1(_1825_),
    .A2(_1830_),
    .B1(_1730_),
    .Y(_1831_));
 sky130_fd_sc_hd__o31ai_1 _4195_ (.A1(_1671_),
    .A2(_1816_),
    .A3(_1822_),
    .B1(_1831_),
    .Y(net84));
 sky130_fd_sc_hd__mux4_1 _4196_ (.A0(\rf_reg[271] ),
    .A1(\rf_reg[303] ),
    .A2(\rf_reg[399] ),
    .A3(\rf_reg[431] ),
    .S0(_1812_),
    .S1(_1732_),
    .X(_1832_));
 sky130_fd_sc_hd__mux4_1 _4197_ (.A0(\rf_reg[335] ),
    .A1(\rf_reg[367] ),
    .A2(\rf_reg[463] ),
    .A3(\rf_reg[495] ),
    .S0(_1775_),
    .S1(_1681_),
    .X(_1833_));
 sky130_fd_sc_hd__mux2i_1 _4198_ (.A0(_1832_),
    .A1(_1833_),
    .S(_1685_),
    .Y(_1834_));
 sky130_fd_sc_hd__and2_0 _4199_ (.A(_1673_),
    .B(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(\rf_reg[47] ),
    .A1(\rf_reg[111] ),
    .S(_1760_),
    .X(_1836_));
 sky130_fd_sc_hd__a22o_1 _4201_ (.A1(\rf_reg[79] ),
    .A2(_1739_),
    .B1(_1836_),
    .B2(_1697_),
    .X(_1837_));
 sky130_fd_sc_hd__buf_8 _4202_ (.A(_1701_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2i_1 _4203_ (.A0(\rf_reg[207] ),
    .A1(\rf_reg[239] ),
    .S(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__mux2i_1 _4204_ (.A0(\rf_reg[143] ),
    .A1(\rf_reg[175] ),
    .S(_1705_),
    .Y(_1840_));
 sky130_fd_sc_hd__o22ai_1 _4205_ (.A1(_1700_),
    .A2(_1839_),
    .B1(_1840_),
    .B2(_1743_),
    .Y(_1841_));
 sky130_fd_sc_hd__a211oi_1 _4206_ (.A1(_1691_),
    .A2(_1837_),
    .B1(_1841_),
    .C1(_1708_),
    .Y(_1842_));
 sky130_fd_sc_hd__mux4_1 _4207_ (.A0(\rf_reg[783] ),
    .A1(\rf_reg[815] ),
    .A2(\rf_reg[911] ),
    .A3(\rf_reg[943] ),
    .S0(_1695_),
    .S1(_1785_),
    .X(_1843_));
 sky130_fd_sc_hd__mux4_1 _4208_ (.A0(\rf_reg[527] ),
    .A1(\rf_reg[559] ),
    .A2(\rf_reg[655] ),
    .A3(\rf_reg[687] ),
    .S0(_1787_),
    .S1(_1716_),
    .X(_1844_));
 sky130_fd_sc_hd__a22o_1 _4209_ (.A1(_1746_),
    .A2(_1843_),
    .B1(_1844_),
    .B2(_1719_),
    .X(_1845_));
 sky130_fd_sc_hd__mux4_1 _4210_ (.A0(\rf_reg[847] ),
    .A1(\rf_reg[879] ),
    .A2(\rf_reg[975] ),
    .A3(\rf_reg[1007] ),
    .S0(_1710_),
    .S1(_1807_),
    .X(_1846_));
 sky130_fd_sc_hd__mux4_1 _4211_ (.A0(\rf_reg[591] ),
    .A1(\rf_reg[623] ),
    .A2(\rf_reg[719] ),
    .A3(\rf_reg[751] ),
    .S0(_1828_),
    .S1(_1689_),
    .X(_1847_));
 sky130_fd_sc_hd__a22o_1 _4212_ (.A1(_1751_),
    .A2(_1846_),
    .B1(_1847_),
    .B2(_1728_),
    .X(_1848_));
 sky130_fd_sc_hd__o21ai_1 _4213_ (.A1(_1845_),
    .A2(_1848_),
    .B1(_1730_),
    .Y(_1849_));
 sky130_fd_sc_hd__o31ai_1 _4214_ (.A1(_1671_),
    .A2(_1835_),
    .A3(_1842_),
    .B1(_1849_),
    .Y(net85));
 sky130_fd_sc_hd__mux4_1 _4215_ (.A0(\rf_reg[272] ),
    .A1(\rf_reg[304] ),
    .A2(\rf_reg[400] ),
    .A3(\rf_reg[432] ),
    .S0(_1812_),
    .S1(_1732_),
    .X(_1850_));
 sky130_fd_sc_hd__mux4_1 _4216_ (.A0(\rf_reg[336] ),
    .A1(\rf_reg[368] ),
    .A2(\rf_reg[464] ),
    .A3(\rf_reg[496] ),
    .S0(_1775_),
    .S1(_1681_),
    .X(_1851_));
 sky130_fd_sc_hd__mux2i_2 _4217_ (.A0(_1850_),
    .A1(_1851_),
    .S(_1685_),
    .Y(_1852_));
 sky130_fd_sc_hd__and2_0 _4218_ (.A(_1673_),
    .B(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(\rf_reg[48] ),
    .A1(\rf_reg[112] ),
    .S(_1760_),
    .X(_1854_));
 sky130_fd_sc_hd__a22o_1 _4220_ (.A1(\rf_reg[80] ),
    .A2(_1739_),
    .B1(_1854_),
    .B2(_1697_),
    .X(_1855_));
 sky130_fd_sc_hd__mux2i_1 _4221_ (.A0(\rf_reg[208] ),
    .A1(\rf_reg[240] ),
    .S(_1838_),
    .Y(_1856_));
 sky130_fd_sc_hd__mux2i_1 _4222_ (.A0(\rf_reg[144] ),
    .A1(\rf_reg[176] ),
    .S(_1705_),
    .Y(_1857_));
 sky130_fd_sc_hd__o22ai_1 _4223_ (.A1(_1700_),
    .A2(_1856_),
    .B1(_1857_),
    .B2(_1743_),
    .Y(_1858_));
 sky130_fd_sc_hd__a211oi_1 _4224_ (.A1(_1691_),
    .A2(_1855_),
    .B1(_1858_),
    .C1(_1708_),
    .Y(_1859_));
 sky130_fd_sc_hd__mux4_1 _4225_ (.A0(\rf_reg[784] ),
    .A1(\rf_reg[816] ),
    .A2(\rf_reg[912] ),
    .A3(\rf_reg[944] ),
    .S0(_1695_),
    .S1(_1785_),
    .X(_1860_));
 sky130_fd_sc_hd__buf_8 _4226_ (.A(_1688_),
    .X(_1861_));
 sky130_fd_sc_hd__mux4_1 _4227_ (.A0(\rf_reg[528] ),
    .A1(\rf_reg[560] ),
    .A2(\rf_reg[656] ),
    .A3(\rf_reg[688] ),
    .S0(_1787_),
    .S1(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__a22o_1 _4228_ (.A1(_1746_),
    .A2(_1860_),
    .B1(_1862_),
    .B2(_1719_),
    .X(_1863_));
 sky130_fd_sc_hd__mux4_1 _4229_ (.A0(\rf_reg[848] ),
    .A1(\rf_reg[880] ),
    .A2(\rf_reg[976] ),
    .A3(\rf_reg[1008] ),
    .S0(_1710_),
    .S1(_1807_),
    .X(_1864_));
 sky130_fd_sc_hd__mux4_1 _4230_ (.A0(\rf_reg[592] ),
    .A1(\rf_reg[624] ),
    .A2(\rf_reg[720] ),
    .A3(\rf_reg[752] ),
    .S0(_1828_),
    .S1(_1689_),
    .X(_1865_));
 sky130_fd_sc_hd__a22o_1 _4231_ (.A1(_1751_),
    .A2(_1864_),
    .B1(_1865_),
    .B2(_1728_),
    .X(_1866_));
 sky130_fd_sc_hd__o21ai_1 _4232_ (.A1(_1863_),
    .A2(_1866_),
    .B1(_1730_),
    .Y(_1867_));
 sky130_fd_sc_hd__o31ai_1 _4233_ (.A1(_1671_),
    .A2(_1853_),
    .A3(_1859_),
    .B1(_1867_),
    .Y(net86));
 sky130_fd_sc_hd__buf_12 _4234_ (.A(_1670_),
    .X(_1868_));
 sky130_fd_sc_hd__buf_6 _4235_ (.A(_1672_),
    .X(_1869_));
 sky130_fd_sc_hd__mux4_1 _4236_ (.A0(\rf_reg[273] ),
    .A1(\rf_reg[305] ),
    .A2(\rf_reg[401] ),
    .A3(\rf_reg[433] ),
    .S0(_1812_),
    .S1(_1732_),
    .X(_1870_));
 sky130_fd_sc_hd__mux4_1 _4237_ (.A0(\rf_reg[337] ),
    .A1(\rf_reg[369] ),
    .A2(\rf_reg[465] ),
    .A3(\rf_reg[497] ),
    .S0(_1775_),
    .S1(_1681_),
    .X(_1871_));
 sky130_fd_sc_hd__mux2i_1 _4238_ (.A0(_1870_),
    .A1(_1871_),
    .S(_1685_),
    .Y(_1872_));
 sky130_fd_sc_hd__and2_1 _4239_ (.A(_1869_),
    .B(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(\rf_reg[49] ),
    .A1(\rf_reg[113] ),
    .S(_1760_),
    .X(_1874_));
 sky130_fd_sc_hd__a22o_1 _4241_ (.A1(\rf_reg[81] ),
    .A2(_1739_),
    .B1(_1874_),
    .B2(_1697_),
    .X(_1875_));
 sky130_fd_sc_hd__mux2i_1 _4242_ (.A0(\rf_reg[209] ),
    .A1(\rf_reg[241] ),
    .S(_1838_),
    .Y(_1876_));
 sky130_fd_sc_hd__buf_6 _4243_ (.A(_1701_),
    .X(_1877_));
 sky130_fd_sc_hd__mux2i_1 _4244_ (.A0(\rf_reg[145] ),
    .A1(\rf_reg[177] ),
    .S(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__o22ai_1 _4245_ (.A1(_1700_),
    .A2(_1876_),
    .B1(_1878_),
    .B2(_1743_),
    .Y(_1879_));
 sky130_fd_sc_hd__a211oi_2 _4246_ (.A1(_1691_),
    .A2(_1875_),
    .B1(_1879_),
    .C1(_1708_),
    .Y(_1880_));
 sky130_fd_sc_hd__buf_16 _4247_ (.A(_1674_),
    .X(_1881_));
 sky130_fd_sc_hd__mux4_1 _4248_ (.A0(\rf_reg[785] ),
    .A1(\rf_reg[817] ),
    .A2(\rf_reg[913] ),
    .A3(\rf_reg[945] ),
    .S0(_1881_),
    .S1(_1785_),
    .X(_1882_));
 sky130_fd_sc_hd__mux4_1 _4249_ (.A0(\rf_reg[529] ),
    .A1(\rf_reg[561] ),
    .A2(\rf_reg[657] ),
    .A3(\rf_reg[689] ),
    .S0(_1787_),
    .S1(_1861_),
    .X(_1883_));
 sky130_fd_sc_hd__a22o_1 _4250_ (.A1(_1746_),
    .A2(_1882_),
    .B1(_1883_),
    .B2(_1719_),
    .X(_1884_));
 sky130_fd_sc_hd__mux4_1 _4251_ (.A0(\rf_reg[849] ),
    .A1(\rf_reg[881] ),
    .A2(\rf_reg[977] ),
    .A3(\rf_reg[1009] ),
    .S0(_1710_),
    .S1(_1807_),
    .X(_1885_));
 sky130_fd_sc_hd__mux4_1 _4252_ (.A0(\rf_reg[593] ),
    .A1(\rf_reg[625] ),
    .A2(\rf_reg[721] ),
    .A3(\rf_reg[753] ),
    .S0(_1828_),
    .S1(_1689_),
    .X(_1886_));
 sky130_fd_sc_hd__a22o_1 _4253_ (.A1(_1751_),
    .A2(_1885_),
    .B1(_1886_),
    .B2(_1728_),
    .X(_1887_));
 sky130_fd_sc_hd__o21ai_1 _4254_ (.A1(_1884_),
    .A2(_1887_),
    .B1(_1730_),
    .Y(_1888_));
 sky130_fd_sc_hd__o31ai_4 _4255_ (.A1(_1868_),
    .A2(_1873_),
    .A3(_1880_),
    .B1(_1888_),
    .Y(net87));
 sky130_fd_sc_hd__mux4_1 _4256_ (.A0(\rf_reg[274] ),
    .A1(\rf_reg[306] ),
    .A2(\rf_reg[402] ),
    .A3(\rf_reg[434] ),
    .S0(_1812_),
    .S1(_1732_),
    .X(_1889_));
 sky130_fd_sc_hd__buf_8 _4257_ (.A(_1676_),
    .X(_1890_));
 sky130_fd_sc_hd__mux4_1 _4258_ (.A0(\rf_reg[338] ),
    .A1(\rf_reg[370] ),
    .A2(\rf_reg[466] ),
    .A3(\rf_reg[498] ),
    .S0(_1775_),
    .S1(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__buf_16 _4259_ (.A(_1684_),
    .X(_1892_));
 sky130_fd_sc_hd__mux2i_1 _4260_ (.A0(_1889_),
    .A1(_1891_),
    .S(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__and2_1 _4261_ (.A(_1869_),
    .B(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(\rf_reg[50] ),
    .A1(\rf_reg[114] ),
    .S(_1760_),
    .X(_1895_));
 sky130_fd_sc_hd__a22o_1 _4263_ (.A1(\rf_reg[82] ),
    .A2(_1739_),
    .B1(_1895_),
    .B2(_1697_),
    .X(_1896_));
 sky130_fd_sc_hd__mux2i_1 _4264_ (.A0(\rf_reg[210] ),
    .A1(\rf_reg[242] ),
    .S(_1838_),
    .Y(_1897_));
 sky130_fd_sc_hd__mux2i_1 _4265_ (.A0(\rf_reg[146] ),
    .A1(\rf_reg[178] ),
    .S(_1877_),
    .Y(_1898_));
 sky130_fd_sc_hd__o22ai_2 _4266_ (.A1(_1700_),
    .A2(_1897_),
    .B1(_1898_),
    .B2(_1743_),
    .Y(_1899_));
 sky130_fd_sc_hd__a211oi_4 _4267_ (.A1(_1691_),
    .A2(_1896_),
    .B1(_1899_),
    .C1(_1708_),
    .Y(_1900_));
 sky130_fd_sc_hd__mux4_1 _4268_ (.A0(\rf_reg[786] ),
    .A1(\rf_reg[818] ),
    .A2(\rf_reg[914] ),
    .A3(\rf_reg[946] ),
    .S0(_1881_),
    .S1(_1785_),
    .X(_1901_));
 sky130_fd_sc_hd__mux4_1 _4269_ (.A0(\rf_reg[530] ),
    .A1(\rf_reg[562] ),
    .A2(\rf_reg[658] ),
    .A3(\rf_reg[690] ),
    .S0(_1787_),
    .S1(_1861_),
    .X(_1902_));
 sky130_fd_sc_hd__a22o_1 _4270_ (.A1(_1746_),
    .A2(_1901_),
    .B1(_1902_),
    .B2(_1719_),
    .X(_1903_));
 sky130_fd_sc_hd__mux4_1 _4271_ (.A0(\rf_reg[850] ),
    .A1(\rf_reg[882] ),
    .A2(\rf_reg[978] ),
    .A3(\rf_reg[1010] ),
    .S0(_1710_),
    .S1(_1807_),
    .X(_1904_));
 sky130_fd_sc_hd__buf_6 _4272_ (.A(_1688_),
    .X(_1905_));
 sky130_fd_sc_hd__mux4_1 _4273_ (.A0(\rf_reg[594] ),
    .A1(\rf_reg[626] ),
    .A2(\rf_reg[722] ),
    .A3(\rf_reg[754] ),
    .S0(_1828_),
    .S1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__a22o_1 _4274_ (.A1(_1751_),
    .A2(_1904_),
    .B1(_1906_),
    .B2(_1728_),
    .X(_1907_));
 sky130_fd_sc_hd__o21ai_1 _4275_ (.A1(_1903_),
    .A2(_1907_),
    .B1(_1730_),
    .Y(_1908_));
 sky130_fd_sc_hd__o31ai_4 _4276_ (.A1(_1868_),
    .A2(_1894_),
    .A3(_1900_),
    .B1(_1908_),
    .Y(net88));
 sky130_fd_sc_hd__mux4_1 _4277_ (.A0(\rf_reg[275] ),
    .A1(\rf_reg[307] ),
    .A2(\rf_reg[403] ),
    .A3(\rf_reg[435] ),
    .S0(_1812_),
    .S1(_1732_),
    .X(_1909_));
 sky130_fd_sc_hd__mux4_1 _4278_ (.A0(\rf_reg[339] ),
    .A1(\rf_reg[371] ),
    .A2(\rf_reg[467] ),
    .A3(\rf_reg[499] ),
    .S0(_1775_),
    .S1(_1890_),
    .X(_1910_));
 sky130_fd_sc_hd__mux2i_1 _4279_ (.A0(_1909_),
    .A1(_1910_),
    .S(_1892_),
    .Y(_1911_));
 sky130_fd_sc_hd__and2_1 _4280_ (.A(_1869_),
    .B(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__buf_8 _4281_ (.A(_1690_),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(\rf_reg[51] ),
    .A1(\rf_reg[115] ),
    .S(_1760_),
    .X(_1914_));
 sky130_fd_sc_hd__a22o_1 _4283_ (.A1(\rf_reg[83] ),
    .A2(_1739_),
    .B1(_1914_),
    .B2(_1697_),
    .X(_1915_));
 sky130_fd_sc_hd__buf_6 _4284_ (.A(_1699_),
    .X(_1916_));
 sky130_fd_sc_hd__mux2i_1 _4285_ (.A0(\rf_reg[211] ),
    .A1(\rf_reg[243] ),
    .S(_1838_),
    .Y(_1917_));
 sky130_fd_sc_hd__mux2i_1 _4286_ (.A0(\rf_reg[147] ),
    .A1(\rf_reg[179] ),
    .S(_1877_),
    .Y(_1918_));
 sky130_fd_sc_hd__o22ai_2 _4287_ (.A1(_1916_),
    .A2(_1917_),
    .B1(_1918_),
    .B2(_1743_),
    .Y(_1919_));
 sky130_fd_sc_hd__buf_8 _4288_ (.A(_1672_),
    .X(_1920_));
 sky130_fd_sc_hd__a211oi_4 _4289_ (.A1(_1913_),
    .A2(_1915_),
    .B1(_1919_),
    .C1(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__mux4_1 _4290_ (.A0(\rf_reg[787] ),
    .A1(\rf_reg[819] ),
    .A2(\rf_reg[915] ),
    .A3(\rf_reg[947] ),
    .S0(_1881_),
    .S1(_1785_),
    .X(_1922_));
 sky130_fd_sc_hd__mux4_1 _4291_ (.A0(\rf_reg[531] ),
    .A1(\rf_reg[563] ),
    .A2(\rf_reg[659] ),
    .A3(\rf_reg[691] ),
    .S0(_1787_),
    .S1(_1861_),
    .X(_1923_));
 sky130_fd_sc_hd__buf_6 _4292_ (.A(_1718_),
    .X(_1924_));
 sky130_fd_sc_hd__a22o_1 _4293_ (.A1(_1746_),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__buf_16 _4294_ (.A(_1694_),
    .X(_1926_));
 sky130_fd_sc_hd__mux4_1 _4295_ (.A0(\rf_reg[851] ),
    .A1(\rf_reg[883] ),
    .A2(\rf_reg[979] ),
    .A3(\rf_reg[1011] ),
    .S0(_1926_),
    .S1(_1807_),
    .X(_1927_));
 sky130_fd_sc_hd__mux4_1 _4296_ (.A0(\rf_reg[595] ),
    .A1(\rf_reg[627] ),
    .A2(\rf_reg[723] ),
    .A3(\rf_reg[755] ),
    .S0(_1828_),
    .S1(_1905_),
    .X(_1928_));
 sky130_fd_sc_hd__buf_8 _4297_ (.A(_1727_),
    .X(_1929_));
 sky130_fd_sc_hd__a22o_1 _4298_ (.A1(_1751_),
    .A2(_1927_),
    .B1(_1928_),
    .B2(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__buf_8 _4299_ (.A(_1670_),
    .X(_1931_));
 sky130_fd_sc_hd__o21ai_1 _4300_ (.A1(_1925_),
    .A2(_1930_),
    .B1(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__o31ai_4 _4301_ (.A1(_1868_),
    .A2(_1912_),
    .A3(_1921_),
    .B1(_1932_),
    .Y(net89));
 sky130_fd_sc_hd__buf_8 _4302_ (.A(_1677_),
    .X(_1933_));
 sky130_fd_sc_hd__mux4_1 _4303_ (.A0(\rf_reg[257] ),
    .A1(\rf_reg[289] ),
    .A2(\rf_reg[385] ),
    .A3(\rf_reg[417] ),
    .S0(_1812_),
    .S1(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__mux4_1 _4304_ (.A0(\rf_reg[321] ),
    .A1(\rf_reg[353] ),
    .A2(\rf_reg[449] ),
    .A3(\rf_reg[481] ),
    .S0(_1775_),
    .S1(_1890_),
    .X(_1935_));
 sky130_fd_sc_hd__mux2i_1 _4305_ (.A0(_1934_),
    .A1(_1935_),
    .S(_1892_),
    .Y(_1936_));
 sky130_fd_sc_hd__and2_0 _4306_ (.A(_1869_),
    .B(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__buf_6 _4307_ (.A(_1738_),
    .X(_1938_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(\rf_reg[33] ),
    .A1(\rf_reg[97] ),
    .S(_1760_),
    .X(_1939_));
 sky130_fd_sc_hd__buf_6 _4309_ (.A(_1696_),
    .X(_1940_));
 sky130_fd_sc_hd__a22o_1 _4310_ (.A1(\rf_reg[65] ),
    .A2(_1938_),
    .B1(_1939_),
    .B2(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__mux2i_1 _4311_ (.A0(\rf_reg[193] ),
    .A1(\rf_reg[225] ),
    .S(_1838_),
    .Y(_1942_));
 sky130_fd_sc_hd__mux2i_1 _4312_ (.A0(\rf_reg[129] ),
    .A1(\rf_reg[161] ),
    .S(_1877_),
    .Y(_1943_));
 sky130_fd_sc_hd__buf_6 _4313_ (.A(_1704_),
    .X(_1944_));
 sky130_fd_sc_hd__o22ai_1 _4314_ (.A1(_1916_),
    .A2(_1942_),
    .B1(_1943_),
    .B2(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__a211oi_2 _4315_ (.A1(_1913_),
    .A2(_1941_),
    .B1(_1945_),
    .C1(_1920_),
    .Y(_1946_));
 sky130_fd_sc_hd__buf_8 _4316_ (.A(_1714_),
    .X(_1947_));
 sky130_fd_sc_hd__mux4_1 _4317_ (.A0(\rf_reg[769] ),
    .A1(\rf_reg[801] ),
    .A2(\rf_reg[897] ),
    .A3(\rf_reg[929] ),
    .S0(_1881_),
    .S1(_1785_),
    .X(_1948_));
 sky130_fd_sc_hd__mux4_1 _4318_ (.A0(\rf_reg[513] ),
    .A1(\rf_reg[545] ),
    .A2(\rf_reg[641] ),
    .A3(\rf_reg[673] ),
    .S0(_1787_),
    .S1(_1861_),
    .X(_1949_));
 sky130_fd_sc_hd__a22o_1 _4319_ (.A1(_1947_),
    .A2(_1948_),
    .B1(_1949_),
    .B2(_1924_),
    .X(_1950_));
 sky130_fd_sc_hd__buf_8 _4320_ (.A(_1724_),
    .X(_1951_));
 sky130_fd_sc_hd__mux4_1 _4321_ (.A0(\rf_reg[833] ),
    .A1(\rf_reg[865] ),
    .A2(\rf_reg[961] ),
    .A3(\rf_reg[993] ),
    .S0(_1926_),
    .S1(_1807_),
    .X(_1952_));
 sky130_fd_sc_hd__mux4_1 _4322_ (.A0(\rf_reg[577] ),
    .A1(\rf_reg[609] ),
    .A2(\rf_reg[705] ),
    .A3(\rf_reg[737] ),
    .S0(_1828_),
    .S1(_1905_),
    .X(_1953_));
 sky130_fd_sc_hd__a22o_1 _4323_ (.A1(_1951_),
    .A2(_1952_),
    .B1(_1953_),
    .B2(_1929_),
    .X(_1954_));
 sky130_fd_sc_hd__o21ai_1 _4324_ (.A1(_1950_),
    .A2(_1954_),
    .B1(_1931_),
    .Y(_1955_));
 sky130_fd_sc_hd__o31ai_4 _4325_ (.A1(_1868_),
    .A2(_1937_),
    .A3(_1946_),
    .B1(_1955_),
    .Y(net90));
 sky130_fd_sc_hd__mux4_1 _4326_ (.A0(\rf_reg[276] ),
    .A1(\rf_reg[308] ),
    .A2(\rf_reg[404] ),
    .A3(\rf_reg[436] ),
    .S0(_1812_),
    .S1(_1933_),
    .X(_1956_));
 sky130_fd_sc_hd__mux4_1 _4327_ (.A0(\rf_reg[340] ),
    .A1(\rf_reg[372] ),
    .A2(\rf_reg[468] ),
    .A3(\rf_reg[500] ),
    .S0(_1775_),
    .S1(_1890_),
    .X(_1957_));
 sky130_fd_sc_hd__mux2i_1 _4328_ (.A0(_1956_),
    .A1(_1957_),
    .S(_1892_),
    .Y(_1958_));
 sky130_fd_sc_hd__and2_1 _4329_ (.A(_1869_),
    .B(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__buf_8 _4330_ (.A(_1683_),
    .X(_1960_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(\rf_reg[52] ),
    .A1(\rf_reg[116] ),
    .S(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__a22o_1 _4332_ (.A1(\rf_reg[84] ),
    .A2(_1938_),
    .B1(_1961_),
    .B2(_1940_),
    .X(_1962_));
 sky130_fd_sc_hd__mux2i_1 _4333_ (.A0(\rf_reg[212] ),
    .A1(\rf_reg[244] ),
    .S(_1838_),
    .Y(_1963_));
 sky130_fd_sc_hd__mux2i_1 _4334_ (.A0(\rf_reg[148] ),
    .A1(\rf_reg[180] ),
    .S(_1877_),
    .Y(_1964_));
 sky130_fd_sc_hd__o22ai_1 _4335_ (.A1(_1916_),
    .A2(_1963_),
    .B1(_1964_),
    .B2(_1944_),
    .Y(_1965_));
 sky130_fd_sc_hd__a211oi_2 _4336_ (.A1(_1913_),
    .A2(_1962_),
    .B1(_1965_),
    .C1(_1920_),
    .Y(_1966_));
 sky130_fd_sc_hd__mux4_1 _4337_ (.A0(\rf_reg[788] ),
    .A1(\rf_reg[820] ),
    .A2(\rf_reg[916] ),
    .A3(\rf_reg[948] ),
    .S0(_1881_),
    .S1(_1785_),
    .X(_1967_));
 sky130_fd_sc_hd__mux4_1 _4338_ (.A0(\rf_reg[532] ),
    .A1(\rf_reg[564] ),
    .A2(\rf_reg[660] ),
    .A3(\rf_reg[692] ),
    .S0(_1787_),
    .S1(_1861_),
    .X(_1968_));
 sky130_fd_sc_hd__a22o_1 _4339_ (.A1(_1947_),
    .A2(_1967_),
    .B1(_1968_),
    .B2(_1924_),
    .X(_1969_));
 sky130_fd_sc_hd__mux4_1 _4340_ (.A0(\rf_reg[852] ),
    .A1(\rf_reg[884] ),
    .A2(\rf_reg[980] ),
    .A3(\rf_reg[1012] ),
    .S0(_1926_),
    .S1(_1807_),
    .X(_1970_));
 sky130_fd_sc_hd__mux4_1 _4341_ (.A0(\rf_reg[596] ),
    .A1(\rf_reg[628] ),
    .A2(\rf_reg[724] ),
    .A3(\rf_reg[756] ),
    .S0(_1828_),
    .S1(_1905_),
    .X(_1971_));
 sky130_fd_sc_hd__a22o_1 _4342_ (.A1(_1951_),
    .A2(_1970_),
    .B1(_1971_),
    .B2(_1929_),
    .X(_1972_));
 sky130_fd_sc_hd__o21ai_1 _4343_ (.A1(_1969_),
    .A2(_1972_),
    .B1(_1931_),
    .Y(_1973_));
 sky130_fd_sc_hd__o31ai_4 _4344_ (.A1(_1868_),
    .A2(_1959_),
    .A3(_1966_),
    .B1(_1973_),
    .Y(net91));
 sky130_fd_sc_hd__mux4_1 _4345_ (.A0(\rf_reg[277] ),
    .A1(\rf_reg[309] ),
    .A2(\rf_reg[405] ),
    .A3(\rf_reg[437] ),
    .S0(_1812_),
    .S1(_1933_),
    .X(_1974_));
 sky130_fd_sc_hd__buf_8 _4346_ (.A(_1674_),
    .X(_1975_));
 sky130_fd_sc_hd__mux4_1 _4347_ (.A0(\rf_reg[341] ),
    .A1(\rf_reg[373] ),
    .A2(\rf_reg[469] ),
    .A3(\rf_reg[501] ),
    .S0(_1975_),
    .S1(_1890_),
    .X(_1976_));
 sky130_fd_sc_hd__mux2i_1 _4348_ (.A0(_1974_),
    .A1(_1976_),
    .S(_1892_),
    .Y(_1977_));
 sky130_fd_sc_hd__and2_1 _4349_ (.A(_1869_),
    .B(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(\rf_reg[53] ),
    .A1(\rf_reg[117] ),
    .S(_1960_),
    .X(_1979_));
 sky130_fd_sc_hd__a22o_1 _4351_ (.A1(\rf_reg[85] ),
    .A2(_1938_),
    .B1(_1979_),
    .B2(_1940_),
    .X(_1980_));
 sky130_fd_sc_hd__mux2i_1 _4352_ (.A0(\rf_reg[213] ),
    .A1(\rf_reg[245] ),
    .S(_1838_),
    .Y(_1981_));
 sky130_fd_sc_hd__mux2i_1 _4353_ (.A0(\rf_reg[149] ),
    .A1(\rf_reg[181] ),
    .S(_1877_),
    .Y(_1982_));
 sky130_fd_sc_hd__o22ai_1 _4354_ (.A1(_1916_),
    .A2(_1981_),
    .B1(_1982_),
    .B2(_1944_),
    .Y(_1983_));
 sky130_fd_sc_hd__a211oi_2 _4355_ (.A1(_1913_),
    .A2(_1980_),
    .B1(_1983_),
    .C1(_1920_),
    .Y(_1984_));
 sky130_fd_sc_hd__buf_8 _4356_ (.A(_1677_),
    .X(_1985_));
 sky130_fd_sc_hd__mux4_1 _4357_ (.A0(\rf_reg[789] ),
    .A1(\rf_reg[821] ),
    .A2(\rf_reg[917] ),
    .A3(\rf_reg[949] ),
    .S0(_1881_),
    .S1(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__buf_16 _4358_ (.A(_1694_),
    .X(_1987_));
 sky130_fd_sc_hd__mux4_1 _4359_ (.A0(\rf_reg[533] ),
    .A1(\rf_reg[565] ),
    .A2(\rf_reg[661] ),
    .A3(\rf_reg[693] ),
    .S0(_1987_),
    .S1(_1861_),
    .X(_1988_));
 sky130_fd_sc_hd__a22o_1 _4360_ (.A1(_1947_),
    .A2(_1986_),
    .B1(_1988_),
    .B2(_1924_),
    .X(_1989_));
 sky130_fd_sc_hd__mux4_1 _4361_ (.A0(\rf_reg[853] ),
    .A1(\rf_reg[885] ),
    .A2(\rf_reg[981] ),
    .A3(\rf_reg[1013] ),
    .S0(_1926_),
    .S1(_1807_),
    .X(_1990_));
 sky130_fd_sc_hd__mux4_1 _4362_ (.A0(\rf_reg[597] ),
    .A1(\rf_reg[629] ),
    .A2(\rf_reg[725] ),
    .A3(\rf_reg[757] ),
    .S0(_1828_),
    .S1(_1905_),
    .X(_1991_));
 sky130_fd_sc_hd__a22o_1 _4363_ (.A1(_1951_),
    .A2(_1990_),
    .B1(_1991_),
    .B2(_1929_),
    .X(_1992_));
 sky130_fd_sc_hd__o21ai_1 _4364_ (.A1(_1989_),
    .A2(_1992_),
    .B1(_1931_),
    .Y(_1993_));
 sky130_fd_sc_hd__o31ai_4 _4365_ (.A1(_1868_),
    .A2(_1978_),
    .A3(_1984_),
    .B1(_1993_),
    .Y(net92));
 sky130_fd_sc_hd__mux4_1 _4366_ (.A0(\rf_reg[278] ),
    .A1(\rf_reg[310] ),
    .A2(\rf_reg[406] ),
    .A3(\rf_reg[438] ),
    .S0(_1812_),
    .S1(_1933_),
    .X(_1994_));
 sky130_fd_sc_hd__mux4_1 _4367_ (.A0(\rf_reg[342] ),
    .A1(\rf_reg[374] ),
    .A2(\rf_reg[470] ),
    .A3(\rf_reg[502] ),
    .S0(_1975_),
    .S1(_1890_),
    .X(_1995_));
 sky130_fd_sc_hd__mux2i_1 _4368_ (.A0(_1994_),
    .A1(_1995_),
    .S(_1892_),
    .Y(_1996_));
 sky130_fd_sc_hd__and2_1 _4369_ (.A(_1869_),
    .B(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(\rf_reg[54] ),
    .A1(\rf_reg[118] ),
    .S(_1960_),
    .X(_1998_));
 sky130_fd_sc_hd__a22o_1 _4371_ (.A1(\rf_reg[86] ),
    .A2(_1938_),
    .B1(_1998_),
    .B2(_1940_),
    .X(_1999_));
 sky130_fd_sc_hd__mux2i_1 _4372_ (.A0(\rf_reg[214] ),
    .A1(\rf_reg[246] ),
    .S(_1838_),
    .Y(_2000_));
 sky130_fd_sc_hd__mux2i_1 _4373_ (.A0(\rf_reg[150] ),
    .A1(\rf_reg[182] ),
    .S(_1877_),
    .Y(_2001_));
 sky130_fd_sc_hd__o22ai_1 _4374_ (.A1(_1916_),
    .A2(_2000_),
    .B1(_2001_),
    .B2(_1944_),
    .Y(_2002_));
 sky130_fd_sc_hd__a211oi_2 _4375_ (.A1(_1913_),
    .A2(_1999_),
    .B1(_2002_),
    .C1(_1920_),
    .Y(_2003_));
 sky130_fd_sc_hd__mux4_1 _4376_ (.A0(\rf_reg[790] ),
    .A1(\rf_reg[822] ),
    .A2(\rf_reg[918] ),
    .A3(\rf_reg[950] ),
    .S0(_1881_),
    .S1(_1985_),
    .X(_2004_));
 sky130_fd_sc_hd__mux4_1 _4377_ (.A0(\rf_reg[534] ),
    .A1(\rf_reg[566] ),
    .A2(\rf_reg[662] ),
    .A3(\rf_reg[694] ),
    .S0(_1987_),
    .S1(_1861_),
    .X(_2005_));
 sky130_fd_sc_hd__a22o_1 _4378_ (.A1(_1947_),
    .A2(_2004_),
    .B1(_2005_),
    .B2(_1924_),
    .X(_2006_));
 sky130_fd_sc_hd__buf_16 _4379_ (.A(_1677_),
    .X(_2007_));
 sky130_fd_sc_hd__mux4_1 _4380_ (.A0(\rf_reg[854] ),
    .A1(\rf_reg[886] ),
    .A2(\rf_reg[982] ),
    .A3(\rf_reg[1014] ),
    .S0(_1926_),
    .S1(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__mux4_1 _4381_ (.A0(\rf_reg[598] ),
    .A1(\rf_reg[630] ),
    .A2(\rf_reg[726] ),
    .A3(\rf_reg[758] ),
    .S0(_1828_),
    .S1(_1905_),
    .X(_2009_));
 sky130_fd_sc_hd__a22o_1 _4382_ (.A1(_1951_),
    .A2(_2008_),
    .B1(_2009_),
    .B2(_1929_),
    .X(_2010_));
 sky130_fd_sc_hd__o21ai_1 _4383_ (.A1(_2006_),
    .A2(_2010_),
    .B1(_1931_),
    .Y(_2011_));
 sky130_fd_sc_hd__o31ai_4 _4384_ (.A1(_1868_),
    .A2(_1997_),
    .A3(_2003_),
    .B1(_2011_),
    .Y(net93));
 sky130_fd_sc_hd__buf_8 _4385_ (.A(_1674_),
    .X(_2012_));
 sky130_fd_sc_hd__mux4_1 _4386_ (.A0(\rf_reg[279] ),
    .A1(\rf_reg[311] ),
    .A2(\rf_reg[407] ),
    .A3(\rf_reg[439] ),
    .S0(_2012_),
    .S1(_1933_),
    .X(_2013_));
 sky130_fd_sc_hd__mux4_1 _4387_ (.A0(\rf_reg[343] ),
    .A1(\rf_reg[375] ),
    .A2(\rf_reg[471] ),
    .A3(\rf_reg[503] ),
    .S0(_1975_),
    .S1(_1890_),
    .X(_2014_));
 sky130_fd_sc_hd__mux2i_1 _4388_ (.A0(_2013_),
    .A1(_2014_),
    .S(_1892_),
    .Y(_2015_));
 sky130_fd_sc_hd__and2_1 _4389_ (.A(_1869_),
    .B(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__mux2_1 _4390_ (.A0(\rf_reg[55] ),
    .A1(\rf_reg[119] ),
    .S(_1960_),
    .X(_2017_));
 sky130_fd_sc_hd__a22o_1 _4391_ (.A1(\rf_reg[87] ),
    .A2(_1938_),
    .B1(_2017_),
    .B2(_1940_),
    .X(_2018_));
 sky130_fd_sc_hd__mux2i_1 _4392_ (.A0(\rf_reg[215] ),
    .A1(\rf_reg[247] ),
    .S(_1838_),
    .Y(_2019_));
 sky130_fd_sc_hd__mux2i_1 _4393_ (.A0(\rf_reg[151] ),
    .A1(\rf_reg[183] ),
    .S(_1877_),
    .Y(_2020_));
 sky130_fd_sc_hd__o22ai_2 _4394_ (.A1(_1916_),
    .A2(_2019_),
    .B1(_2020_),
    .B2(_1944_),
    .Y(_2021_));
 sky130_fd_sc_hd__a211oi_4 _4395_ (.A1(_1913_),
    .A2(_2018_),
    .B1(_2021_),
    .C1(_1920_),
    .Y(_2022_));
 sky130_fd_sc_hd__mux4_1 _4396_ (.A0(\rf_reg[791] ),
    .A1(\rf_reg[823] ),
    .A2(\rf_reg[919] ),
    .A3(\rf_reg[951] ),
    .S0(_1881_),
    .S1(_1985_),
    .X(_2023_));
 sky130_fd_sc_hd__mux4_1 _4397_ (.A0(\rf_reg[535] ),
    .A1(\rf_reg[567] ),
    .A2(\rf_reg[663] ),
    .A3(\rf_reg[695] ),
    .S0(_1987_),
    .S1(_1861_),
    .X(_2024_));
 sky130_fd_sc_hd__a22o_1 _4398_ (.A1(_1947_),
    .A2(_2023_),
    .B1(_2024_),
    .B2(_1924_),
    .X(_2025_));
 sky130_fd_sc_hd__mux4_1 _4399_ (.A0(\rf_reg[855] ),
    .A1(\rf_reg[887] ),
    .A2(\rf_reg[983] ),
    .A3(\rf_reg[1015] ),
    .S0(_1926_),
    .S1(_2007_),
    .X(_2026_));
 sky130_fd_sc_hd__buf_8 _4400_ (.A(_1694_),
    .X(_2027_));
 sky130_fd_sc_hd__mux4_1 _4401_ (.A0(\rf_reg[599] ),
    .A1(\rf_reg[631] ),
    .A2(\rf_reg[727] ),
    .A3(\rf_reg[759] ),
    .S0(_2027_),
    .S1(_1905_),
    .X(_2028_));
 sky130_fd_sc_hd__a22o_1 _4402_ (.A1(_1951_),
    .A2(_2026_),
    .B1(_2028_),
    .B2(_1929_),
    .X(_2029_));
 sky130_fd_sc_hd__o21ai_1 _4403_ (.A1(_2025_),
    .A2(_2029_),
    .B1(_1931_),
    .Y(_2030_));
 sky130_fd_sc_hd__o31ai_4 _4404_ (.A1(_1868_),
    .A2(_2016_),
    .A3(_2022_),
    .B1(_2030_),
    .Y(net94));
 sky130_fd_sc_hd__mux4_1 _4405_ (.A0(\rf_reg[280] ),
    .A1(\rf_reg[312] ),
    .A2(\rf_reg[408] ),
    .A3(\rf_reg[440] ),
    .S0(_2012_),
    .S1(_1933_),
    .X(_2031_));
 sky130_fd_sc_hd__mux4_1 _4406_ (.A0(\rf_reg[344] ),
    .A1(\rf_reg[376] ),
    .A2(\rf_reg[472] ),
    .A3(\rf_reg[504] ),
    .S0(_1975_),
    .S1(_1890_),
    .X(_2032_));
 sky130_fd_sc_hd__mux2i_1 _4407_ (.A0(_2031_),
    .A1(_2032_),
    .S(_1892_),
    .Y(_2033_));
 sky130_fd_sc_hd__and2_1 _4408_ (.A(_1869_),
    .B(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__mux2_1 _4409_ (.A0(\rf_reg[56] ),
    .A1(\rf_reg[120] ),
    .S(_1960_),
    .X(_2035_));
 sky130_fd_sc_hd__a22o_1 _4410_ (.A1(\rf_reg[88] ),
    .A2(_1938_),
    .B1(_2035_),
    .B2(_1940_),
    .X(_2036_));
 sky130_fd_sc_hd__buf_8 _4411_ (.A(_1701_),
    .X(_2037_));
 sky130_fd_sc_hd__mux2i_2 _4412_ (.A0(\rf_reg[216] ),
    .A1(\rf_reg[248] ),
    .S(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__mux2i_2 _4413_ (.A0(\rf_reg[152] ),
    .A1(\rf_reg[184] ),
    .S(_1877_),
    .Y(_2039_));
 sky130_fd_sc_hd__o22ai_4 _4414_ (.A1(_1916_),
    .A2(_2038_),
    .B1(_2039_),
    .B2(_1944_),
    .Y(_2040_));
 sky130_fd_sc_hd__a211oi_4 _4415_ (.A1(_1913_),
    .A2(_2036_),
    .B1(_2040_),
    .C1(_1920_),
    .Y(_2041_));
 sky130_fd_sc_hd__mux4_1 _4416_ (.A0(\rf_reg[792] ),
    .A1(\rf_reg[824] ),
    .A2(\rf_reg[920] ),
    .A3(\rf_reg[952] ),
    .S0(_1881_),
    .S1(_1985_),
    .X(_2042_));
 sky130_fd_sc_hd__mux4_1 _4417_ (.A0(\rf_reg[536] ),
    .A1(\rf_reg[568] ),
    .A2(\rf_reg[664] ),
    .A3(\rf_reg[696] ),
    .S0(_1987_),
    .S1(_1861_),
    .X(_2043_));
 sky130_fd_sc_hd__a22o_1 _4418_ (.A1(_1947_),
    .A2(_2042_),
    .B1(_2043_),
    .B2(_1924_),
    .X(_2044_));
 sky130_fd_sc_hd__mux4_1 _4419_ (.A0(\rf_reg[856] ),
    .A1(\rf_reg[888] ),
    .A2(\rf_reg[984] ),
    .A3(\rf_reg[1016] ),
    .S0(_1926_),
    .S1(_2007_),
    .X(_2045_));
 sky130_fd_sc_hd__mux4_1 _4420_ (.A0(\rf_reg[600] ),
    .A1(\rf_reg[632] ),
    .A2(\rf_reg[728] ),
    .A3(\rf_reg[760] ),
    .S0(_2027_),
    .S1(_1905_),
    .X(_2046_));
 sky130_fd_sc_hd__a22o_1 _4421_ (.A1(_1951_),
    .A2(_2045_),
    .B1(_2046_),
    .B2(_1929_),
    .X(_2047_));
 sky130_fd_sc_hd__o21ai_2 _4422_ (.A1(_2044_),
    .A2(_2047_),
    .B1(_1931_),
    .Y(_2048_));
 sky130_fd_sc_hd__o31ai_4 _4423_ (.A1(_1868_),
    .A2(_2034_),
    .A3(_2041_),
    .B1(_2048_),
    .Y(net95));
 sky130_fd_sc_hd__mux4_1 _4424_ (.A0(\rf_reg[281] ),
    .A1(\rf_reg[313] ),
    .A2(\rf_reg[409] ),
    .A3(\rf_reg[441] ),
    .S0(_2012_),
    .S1(_1933_),
    .X(_2049_));
 sky130_fd_sc_hd__mux4_1 _4425_ (.A0(\rf_reg[345] ),
    .A1(\rf_reg[377] ),
    .A2(\rf_reg[473] ),
    .A3(\rf_reg[505] ),
    .S0(_1975_),
    .S1(_1890_),
    .X(_2050_));
 sky130_fd_sc_hd__mux2i_1 _4426_ (.A0(_2049_),
    .A1(_2050_),
    .S(_1892_),
    .Y(_2051_));
 sky130_fd_sc_hd__and2_0 _4427_ (.A(_1869_),
    .B(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__mux2_1 _4428_ (.A0(\rf_reg[57] ),
    .A1(\rf_reg[121] ),
    .S(_1960_),
    .X(_2053_));
 sky130_fd_sc_hd__a22o_1 _4429_ (.A1(\rf_reg[89] ),
    .A2(_1938_),
    .B1(_2053_),
    .B2(_1940_),
    .X(_2054_));
 sky130_fd_sc_hd__mux2i_1 _4430_ (.A0(\rf_reg[217] ),
    .A1(\rf_reg[249] ),
    .S(_2037_),
    .Y(_2055_));
 sky130_fd_sc_hd__mux2i_1 _4431_ (.A0(\rf_reg[153] ),
    .A1(\rf_reg[185] ),
    .S(_1877_),
    .Y(_2056_));
 sky130_fd_sc_hd__o22ai_2 _4432_ (.A1(_1916_),
    .A2(_2055_),
    .B1(_2056_),
    .B2(_1944_),
    .Y(_2057_));
 sky130_fd_sc_hd__a211oi_4 _4433_ (.A1(_1913_),
    .A2(_2054_),
    .B1(_2057_),
    .C1(_1920_),
    .Y(_2058_));
 sky130_fd_sc_hd__mux4_1 _4434_ (.A0(\rf_reg[793] ),
    .A1(\rf_reg[825] ),
    .A2(\rf_reg[921] ),
    .A3(\rf_reg[953] ),
    .S0(_1881_),
    .S1(_1985_),
    .X(_2059_));
 sky130_fd_sc_hd__buf_8 _4435_ (.A(_1688_),
    .X(_2060_));
 sky130_fd_sc_hd__mux4_1 _4436_ (.A0(\rf_reg[537] ),
    .A1(\rf_reg[569] ),
    .A2(\rf_reg[665] ),
    .A3(\rf_reg[697] ),
    .S0(_1987_),
    .S1(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__a22o_1 _4437_ (.A1(_1947_),
    .A2(_2059_),
    .B1(_2061_),
    .B2(_1924_),
    .X(_2062_));
 sky130_fd_sc_hd__mux4_1 _4438_ (.A0(\rf_reg[857] ),
    .A1(\rf_reg[889] ),
    .A2(\rf_reg[985] ),
    .A3(\rf_reg[1017] ),
    .S0(_1926_),
    .S1(_2007_),
    .X(_2063_));
 sky130_fd_sc_hd__mux4_1 _4439_ (.A0(\rf_reg[601] ),
    .A1(\rf_reg[633] ),
    .A2(\rf_reg[729] ),
    .A3(\rf_reg[761] ),
    .S0(_2027_),
    .S1(_1905_),
    .X(_2064_));
 sky130_fd_sc_hd__a22o_1 _4440_ (.A1(_1951_),
    .A2(_2063_),
    .B1(_2064_),
    .B2(_1929_),
    .X(_2065_));
 sky130_fd_sc_hd__o21ai_2 _4441_ (.A1(_2062_),
    .A2(_2065_),
    .B1(_1931_),
    .Y(_2066_));
 sky130_fd_sc_hd__o31ai_4 _4442_ (.A1(_1868_),
    .A2(_2052_),
    .A3(_2058_),
    .B1(_2066_),
    .Y(net96));
 sky130_fd_sc_hd__buf_12 _4443_ (.A(_1670_),
    .X(_2067_));
 sky130_fd_sc_hd__buf_6 _4444_ (.A(_1672_),
    .X(_2068_));
 sky130_fd_sc_hd__mux4_1 _4445_ (.A0(\rf_reg[282] ),
    .A1(\rf_reg[314] ),
    .A2(\rf_reg[410] ),
    .A3(\rf_reg[442] ),
    .S0(_2012_),
    .S1(_1933_),
    .X(_2069_));
 sky130_fd_sc_hd__mux4_1 _4446_ (.A0(\rf_reg[346] ),
    .A1(\rf_reg[378] ),
    .A2(\rf_reg[474] ),
    .A3(\rf_reg[506] ),
    .S0(_1975_),
    .S1(_1890_),
    .X(_2070_));
 sky130_fd_sc_hd__mux2i_1 _4447_ (.A0(_2069_),
    .A1(_2070_),
    .S(_1892_),
    .Y(_2071_));
 sky130_fd_sc_hd__and2_0 _4448_ (.A(_2068_),
    .B(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(\rf_reg[58] ),
    .A1(\rf_reg[122] ),
    .S(_1960_),
    .X(_2073_));
 sky130_fd_sc_hd__a22o_1 _4450_ (.A1(\rf_reg[90] ),
    .A2(_1938_),
    .B1(_2073_),
    .B2(_1940_),
    .X(_2074_));
 sky130_fd_sc_hd__mux2i_1 _4451_ (.A0(\rf_reg[218] ),
    .A1(\rf_reg[250] ),
    .S(_2037_),
    .Y(_2075_));
 sky130_fd_sc_hd__buf_8 _4452_ (.A(_1701_),
    .X(_2076_));
 sky130_fd_sc_hd__mux2i_1 _4453_ (.A0(\rf_reg[154] ),
    .A1(\rf_reg[186] ),
    .S(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__o22ai_1 _4454_ (.A1(_1916_),
    .A2(_2075_),
    .B1(_2077_),
    .B2(_1944_),
    .Y(_2078_));
 sky130_fd_sc_hd__a211oi_2 _4455_ (.A1(_1913_),
    .A2(_2074_),
    .B1(_2078_),
    .C1(_1920_),
    .Y(_2079_));
 sky130_fd_sc_hd__buf_16 _4456_ (.A(_1674_),
    .X(_2080_));
 sky130_fd_sc_hd__mux4_1 _4457_ (.A0(\rf_reg[794] ),
    .A1(\rf_reg[826] ),
    .A2(\rf_reg[922] ),
    .A3(\rf_reg[954] ),
    .S0(_2080_),
    .S1(_1985_),
    .X(_2081_));
 sky130_fd_sc_hd__mux4_1 _4458_ (.A0(\rf_reg[538] ),
    .A1(\rf_reg[570] ),
    .A2(\rf_reg[666] ),
    .A3(\rf_reg[698] ),
    .S0(_1987_),
    .S1(_2060_),
    .X(_2082_));
 sky130_fd_sc_hd__a22o_1 _4459_ (.A1(_1947_),
    .A2(_2081_),
    .B1(_2082_),
    .B2(_1924_),
    .X(_2083_));
 sky130_fd_sc_hd__mux4_1 _4460_ (.A0(\rf_reg[858] ),
    .A1(\rf_reg[890] ),
    .A2(\rf_reg[986] ),
    .A3(\rf_reg[1018] ),
    .S0(_1926_),
    .S1(_2007_),
    .X(_2084_));
 sky130_fd_sc_hd__mux4_1 _4461_ (.A0(\rf_reg[602] ),
    .A1(\rf_reg[634] ),
    .A2(\rf_reg[730] ),
    .A3(\rf_reg[762] ),
    .S0(_2027_),
    .S1(_1905_),
    .X(_2085_));
 sky130_fd_sc_hd__a22o_1 _4462_ (.A1(_1951_),
    .A2(_2084_),
    .B1(_2085_),
    .B2(_1929_),
    .X(_2086_));
 sky130_fd_sc_hd__o21ai_2 _4463_ (.A1(_2083_),
    .A2(_2086_),
    .B1(_1931_),
    .Y(_2087_));
 sky130_fd_sc_hd__o31ai_4 _4464_ (.A1(_2067_),
    .A2(_2072_),
    .A3(_2079_),
    .B1(_2087_),
    .Y(net97));
 sky130_fd_sc_hd__mux4_1 _4465_ (.A0(\rf_reg[283] ),
    .A1(\rf_reg[315] ),
    .A2(\rf_reg[411] ),
    .A3(\rf_reg[443] ),
    .S0(_2012_),
    .S1(_1933_),
    .X(_2088_));
 sky130_fd_sc_hd__buf_8 _4466_ (.A(_1676_),
    .X(_2089_));
 sky130_fd_sc_hd__mux4_1 _4467_ (.A0(\rf_reg[347] ),
    .A1(\rf_reg[379] ),
    .A2(\rf_reg[475] ),
    .A3(\rf_reg[507] ),
    .S0(_1975_),
    .S1(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__clkbuf_16 _4468_ (.A(_1684_),
    .X(_2091_));
 sky130_fd_sc_hd__mux2i_1 _4469_ (.A0(_2088_),
    .A1(_2090_),
    .S(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__and2_0 _4470_ (.A(_2068_),
    .B(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(\rf_reg[59] ),
    .A1(\rf_reg[123] ),
    .S(_1960_),
    .X(_2094_));
 sky130_fd_sc_hd__a22o_1 _4472_ (.A1(\rf_reg[91] ),
    .A2(_1938_),
    .B1(_2094_),
    .B2(_1940_),
    .X(_2095_));
 sky130_fd_sc_hd__mux2i_1 _4473_ (.A0(\rf_reg[219] ),
    .A1(\rf_reg[251] ),
    .S(_2037_),
    .Y(_2096_));
 sky130_fd_sc_hd__mux2i_1 _4474_ (.A0(\rf_reg[155] ),
    .A1(\rf_reg[187] ),
    .S(_2076_),
    .Y(_2097_));
 sky130_fd_sc_hd__o22ai_1 _4475_ (.A1(_1916_),
    .A2(_2096_),
    .B1(_2097_),
    .B2(_1944_),
    .Y(_2098_));
 sky130_fd_sc_hd__a211oi_2 _4476_ (.A1(_1913_),
    .A2(_2095_),
    .B1(_2098_),
    .C1(_1920_),
    .Y(_2099_));
 sky130_fd_sc_hd__mux4_1 _4477_ (.A0(\rf_reg[795] ),
    .A1(\rf_reg[827] ),
    .A2(\rf_reg[923] ),
    .A3(\rf_reg[955] ),
    .S0(_2080_),
    .S1(_1985_),
    .X(_2100_));
 sky130_fd_sc_hd__mux4_1 _4478_ (.A0(\rf_reg[539] ),
    .A1(\rf_reg[571] ),
    .A2(\rf_reg[667] ),
    .A3(\rf_reg[699] ),
    .S0(_1987_),
    .S1(_2060_),
    .X(_2101_));
 sky130_fd_sc_hd__a22o_1 _4479_ (.A1(_1947_),
    .A2(_2100_),
    .B1(_2101_),
    .B2(_1924_),
    .X(_2102_));
 sky130_fd_sc_hd__mux4_1 _4480_ (.A0(\rf_reg[859] ),
    .A1(\rf_reg[891] ),
    .A2(\rf_reg[987] ),
    .A3(\rf_reg[1019] ),
    .S0(_1926_),
    .S1(_2007_),
    .X(_2103_));
 sky130_fd_sc_hd__buf_8 _4481_ (.A(_1688_),
    .X(_2104_));
 sky130_fd_sc_hd__mux4_1 _4482_ (.A0(\rf_reg[603] ),
    .A1(\rf_reg[635] ),
    .A2(\rf_reg[731] ),
    .A3(\rf_reg[763] ),
    .S0(_2027_),
    .S1(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__a22o_1 _4483_ (.A1(_1951_),
    .A2(_2103_),
    .B1(_2105_),
    .B2(_1929_),
    .X(_2106_));
 sky130_fd_sc_hd__o21ai_2 _4484_ (.A1(_2102_),
    .A2(_2106_),
    .B1(_1931_),
    .Y(_2107_));
 sky130_fd_sc_hd__o31ai_4 _4485_ (.A1(_2067_),
    .A2(_2093_),
    .A3(_2099_),
    .B1(_2107_),
    .Y(net98));
 sky130_fd_sc_hd__mux4_1 _4486_ (.A0(\rf_reg[284] ),
    .A1(\rf_reg[316] ),
    .A2(\rf_reg[412] ),
    .A3(\rf_reg[444] ),
    .S0(_2012_),
    .S1(_1933_),
    .X(_2108_));
 sky130_fd_sc_hd__mux4_1 _4487_ (.A0(\rf_reg[348] ),
    .A1(\rf_reg[380] ),
    .A2(\rf_reg[476] ),
    .A3(\rf_reg[508] ),
    .S0(_1975_),
    .S1(_2089_),
    .X(_2109_));
 sky130_fd_sc_hd__mux2i_1 _4488_ (.A0(_2108_),
    .A1(_2109_),
    .S(_2091_),
    .Y(_2110_));
 sky130_fd_sc_hd__and2_0 _4489_ (.A(_2068_),
    .B(_2110_),
    .X(_2111_));
 sky130_fd_sc_hd__buf_6 _4490_ (.A(_1690_),
    .X(_2112_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(\rf_reg[60] ),
    .A1(\rf_reg[124] ),
    .S(_1960_),
    .X(_2113_));
 sky130_fd_sc_hd__a22o_1 _4492_ (.A1(\rf_reg[92] ),
    .A2(_1938_),
    .B1(_2113_),
    .B2(_1940_),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_8 _4493_ (.A(_1699_),
    .X(_2115_));
 sky130_fd_sc_hd__mux2i_1 _4494_ (.A0(\rf_reg[220] ),
    .A1(\rf_reg[252] ),
    .S(_2037_),
    .Y(_2116_));
 sky130_fd_sc_hd__mux2i_1 _4495_ (.A0(\rf_reg[156] ),
    .A1(\rf_reg[188] ),
    .S(_2076_),
    .Y(_2117_));
 sky130_fd_sc_hd__o22ai_1 _4496_ (.A1(_2115_),
    .A2(_2116_),
    .B1(_2117_),
    .B2(_1944_),
    .Y(_2118_));
 sky130_fd_sc_hd__buf_8 _4497_ (.A(_1672_),
    .X(_2119_));
 sky130_fd_sc_hd__a211oi_2 _4498_ (.A1(_2112_),
    .A2(_2114_),
    .B1(_2118_),
    .C1(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__mux4_1 _4499_ (.A0(\rf_reg[796] ),
    .A1(\rf_reg[828] ),
    .A2(\rf_reg[924] ),
    .A3(\rf_reg[956] ),
    .S0(_2080_),
    .S1(_1985_),
    .X(_2121_));
 sky130_fd_sc_hd__mux4_1 _4500_ (.A0(\rf_reg[540] ),
    .A1(\rf_reg[572] ),
    .A2(\rf_reg[668] ),
    .A3(\rf_reg[700] ),
    .S0(_1987_),
    .S1(_2060_),
    .X(_2122_));
 sky130_fd_sc_hd__buf_8 _4501_ (.A(_1718_),
    .X(_2123_));
 sky130_fd_sc_hd__a22o_1 _4502_ (.A1(_1947_),
    .A2(_2121_),
    .B1(_2122_),
    .B2(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__buf_16 _4503_ (.A(_1694_),
    .X(_2125_));
 sky130_fd_sc_hd__mux4_1 _4504_ (.A0(\rf_reg[860] ),
    .A1(\rf_reg[892] ),
    .A2(\rf_reg[988] ),
    .A3(\rf_reg[1020] ),
    .S0(_2125_),
    .S1(_2007_),
    .X(_2126_));
 sky130_fd_sc_hd__mux4_1 _4505_ (.A0(\rf_reg[604] ),
    .A1(\rf_reg[636] ),
    .A2(\rf_reg[732] ),
    .A3(\rf_reg[764] ),
    .S0(_2027_),
    .S1(_2104_),
    .X(_2127_));
 sky130_fd_sc_hd__buf_8 _4506_ (.A(_1727_),
    .X(_2128_));
 sky130_fd_sc_hd__a22o_1 _4507_ (.A1(_1951_),
    .A2(_2126_),
    .B1(_2127_),
    .B2(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__buf_8 _4508_ (.A(_1670_),
    .X(_2130_));
 sky130_fd_sc_hd__o21ai_2 _4509_ (.A1(_2124_),
    .A2(_2129_),
    .B1(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__o31ai_4 _4510_ (.A1(_2067_),
    .A2(_2111_),
    .A3(_2120_),
    .B1(_2131_),
    .Y(net99));
 sky130_fd_sc_hd__buf_8 _4511_ (.A(_1676_),
    .X(_2132_));
 sky130_fd_sc_hd__mux4_1 _4512_ (.A0(\rf_reg[285] ),
    .A1(\rf_reg[317] ),
    .A2(\rf_reg[413] ),
    .A3(\rf_reg[445] ),
    .S0(_2012_),
    .S1(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__mux4_1 _4513_ (.A0(\rf_reg[349] ),
    .A1(\rf_reg[381] ),
    .A2(\rf_reg[477] ),
    .A3(\rf_reg[509] ),
    .S0(_1975_),
    .S1(_2089_),
    .X(_2134_));
 sky130_fd_sc_hd__mux2i_1 _4514_ (.A0(_2133_),
    .A1(_2134_),
    .S(_2091_),
    .Y(_2135_));
 sky130_fd_sc_hd__and2_0 _4515_ (.A(_2068_),
    .B(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__buf_6 _4516_ (.A(_1738_),
    .X(_2137_));
 sky130_fd_sc_hd__mux2_1 _4517_ (.A0(\rf_reg[61] ),
    .A1(\rf_reg[125] ),
    .S(_1960_),
    .X(_2138_));
 sky130_fd_sc_hd__clkbuf_8 _4518_ (.A(_1696_),
    .X(_2139_));
 sky130_fd_sc_hd__a22o_1 _4519_ (.A1(\rf_reg[93] ),
    .A2(_2137_),
    .B1(_2138_),
    .B2(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__mux2i_1 _4520_ (.A0(\rf_reg[221] ),
    .A1(\rf_reg[253] ),
    .S(_2037_),
    .Y(_2141_));
 sky130_fd_sc_hd__mux2i_1 _4521_ (.A0(\rf_reg[157] ),
    .A1(\rf_reg[189] ),
    .S(_2076_),
    .Y(_2142_));
 sky130_fd_sc_hd__clkbuf_8 _4522_ (.A(_1704_),
    .X(_2143_));
 sky130_fd_sc_hd__o22ai_1 _4523_ (.A1(_2115_),
    .A2(_2141_),
    .B1(_2142_),
    .B2(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__a211oi_2 _4524_ (.A1(_2112_),
    .A2(_2140_),
    .B1(_2144_),
    .C1(_2119_),
    .Y(_2145_));
 sky130_fd_sc_hd__buf_8 _4525_ (.A(_1714_),
    .X(_2146_));
 sky130_fd_sc_hd__mux4_1 _4526_ (.A0(\rf_reg[797] ),
    .A1(\rf_reg[829] ),
    .A2(\rf_reg[925] ),
    .A3(\rf_reg[957] ),
    .S0(_2080_),
    .S1(_1985_),
    .X(_2147_));
 sky130_fd_sc_hd__mux4_1 _4527_ (.A0(\rf_reg[541] ),
    .A1(\rf_reg[573] ),
    .A2(\rf_reg[669] ),
    .A3(\rf_reg[701] ),
    .S0(_1987_),
    .S1(_2060_),
    .X(_2148_));
 sky130_fd_sc_hd__a22o_1 _4528_ (.A1(_2146_),
    .A2(_2147_),
    .B1(_2148_),
    .B2(_2123_),
    .X(_2149_));
 sky130_fd_sc_hd__buf_8 _4529_ (.A(_1724_),
    .X(_2150_));
 sky130_fd_sc_hd__mux4_1 _4530_ (.A0(\rf_reg[861] ),
    .A1(\rf_reg[893] ),
    .A2(\rf_reg[989] ),
    .A3(\rf_reg[1021] ),
    .S0(_2125_),
    .S1(_2007_),
    .X(_2151_));
 sky130_fd_sc_hd__mux4_1 _4531_ (.A0(\rf_reg[605] ),
    .A1(\rf_reg[637] ),
    .A2(\rf_reg[733] ),
    .A3(\rf_reg[765] ),
    .S0(_2027_),
    .S1(_2104_),
    .X(_2152_));
 sky130_fd_sc_hd__a22o_1 _4532_ (.A1(_2150_),
    .A2(_2151_),
    .B1(_2152_),
    .B2(_2128_),
    .X(_2153_));
 sky130_fd_sc_hd__o21ai_2 _4533_ (.A1(_2149_),
    .A2(_2153_),
    .B1(_2130_),
    .Y(_2154_));
 sky130_fd_sc_hd__o31ai_4 _4534_ (.A1(_2067_),
    .A2(_2136_),
    .A3(_2145_),
    .B1(_2154_),
    .Y(net100));
 sky130_fd_sc_hd__mux4_1 _4535_ (.A0(\rf_reg[258] ),
    .A1(\rf_reg[290] ),
    .A2(\rf_reg[386] ),
    .A3(\rf_reg[418] ),
    .S0(_2012_),
    .S1(_2132_),
    .X(_2155_));
 sky130_fd_sc_hd__mux4_1 _4536_ (.A0(\rf_reg[322] ),
    .A1(\rf_reg[354] ),
    .A2(\rf_reg[450] ),
    .A3(\rf_reg[482] ),
    .S0(_1975_),
    .S1(_2089_),
    .X(_2156_));
 sky130_fd_sc_hd__mux2i_1 _4537_ (.A0(_2155_),
    .A1(_2156_),
    .S(_2091_),
    .Y(_2157_));
 sky130_fd_sc_hd__and2_0 _4538_ (.A(_2068_),
    .B(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__buf_6 _4539_ (.A(_1683_),
    .X(_2159_));
 sky130_fd_sc_hd__mux2_1 _4540_ (.A0(\rf_reg[34] ),
    .A1(\rf_reg[98] ),
    .S(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__a22o_1 _4541_ (.A1(\rf_reg[66] ),
    .A2(_2137_),
    .B1(_2160_),
    .B2(_2139_),
    .X(_2161_));
 sky130_fd_sc_hd__mux2i_1 _4542_ (.A0(\rf_reg[194] ),
    .A1(\rf_reg[226] ),
    .S(_2037_),
    .Y(_2162_));
 sky130_fd_sc_hd__mux2i_1 _4543_ (.A0(\rf_reg[130] ),
    .A1(\rf_reg[162] ),
    .S(_2076_),
    .Y(_2163_));
 sky130_fd_sc_hd__o22ai_1 _4544_ (.A1(_2115_),
    .A2(_2162_),
    .B1(_2163_),
    .B2(_2143_),
    .Y(_2164_));
 sky130_fd_sc_hd__a211oi_2 _4545_ (.A1(_2112_),
    .A2(_2161_),
    .B1(_2164_),
    .C1(_2119_),
    .Y(_2165_));
 sky130_fd_sc_hd__mux4_1 _4546_ (.A0(\rf_reg[770] ),
    .A1(\rf_reg[802] ),
    .A2(\rf_reg[898] ),
    .A3(\rf_reg[930] ),
    .S0(_2080_),
    .S1(_1985_),
    .X(_2166_));
 sky130_fd_sc_hd__mux4_1 _4547_ (.A0(\rf_reg[514] ),
    .A1(\rf_reg[546] ),
    .A2(\rf_reg[642] ),
    .A3(\rf_reg[674] ),
    .S0(_1987_),
    .S1(_2060_),
    .X(_2167_));
 sky130_fd_sc_hd__a22o_1 _4548_ (.A1(_2146_),
    .A2(_2166_),
    .B1(_2167_),
    .B2(_2123_),
    .X(_2168_));
 sky130_fd_sc_hd__mux4_1 _4549_ (.A0(\rf_reg[834] ),
    .A1(\rf_reg[866] ),
    .A2(\rf_reg[962] ),
    .A3(\rf_reg[994] ),
    .S0(_2125_),
    .S1(_2007_),
    .X(_2169_));
 sky130_fd_sc_hd__mux4_1 _4550_ (.A0(\rf_reg[578] ),
    .A1(\rf_reg[610] ),
    .A2(\rf_reg[706] ),
    .A3(\rf_reg[738] ),
    .S0(_2027_),
    .S1(_2104_),
    .X(_2170_));
 sky130_fd_sc_hd__a22o_1 _4551_ (.A1(_2150_),
    .A2(_2169_),
    .B1(_2170_),
    .B2(_2128_),
    .X(_2171_));
 sky130_fd_sc_hd__o21ai_2 _4552_ (.A1(_2168_),
    .A2(_2171_),
    .B1(_2130_),
    .Y(_2172_));
 sky130_fd_sc_hd__o31ai_4 _4553_ (.A1(_2067_),
    .A2(_2158_),
    .A3(_2165_),
    .B1(_2172_),
    .Y(net101));
 sky130_fd_sc_hd__mux4_1 _4554_ (.A0(\rf_reg[286] ),
    .A1(\rf_reg[318] ),
    .A2(\rf_reg[414] ),
    .A3(\rf_reg[446] ),
    .S0(_2012_),
    .S1(_2132_),
    .X(_2173_));
 sky130_fd_sc_hd__mux4_1 _4555_ (.A0(\rf_reg[350] ),
    .A1(\rf_reg[382] ),
    .A2(\rf_reg[478] ),
    .A3(\rf_reg[510] ),
    .S0(_1827_),
    .S1(_2089_),
    .X(_2174_));
 sky130_fd_sc_hd__mux2i_2 _4556_ (.A0(_2173_),
    .A1(_2174_),
    .S(_2091_),
    .Y(_2175_));
 sky130_fd_sc_hd__and2_0 _4557_ (.A(_2068_),
    .B(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__mux2_1 _4558_ (.A0(\rf_reg[62] ),
    .A1(\rf_reg[126] ),
    .S(_2159_),
    .X(_2177_));
 sky130_fd_sc_hd__a22o_1 _4559_ (.A1(\rf_reg[94] ),
    .A2(_2137_),
    .B1(_2177_),
    .B2(_2139_),
    .X(_2178_));
 sky130_fd_sc_hd__mux2i_1 _4560_ (.A0(\rf_reg[222] ),
    .A1(\rf_reg[254] ),
    .S(_2037_),
    .Y(_2179_));
 sky130_fd_sc_hd__mux2i_1 _4561_ (.A0(\rf_reg[158] ),
    .A1(\rf_reg[190] ),
    .S(_2076_),
    .Y(_2180_));
 sky130_fd_sc_hd__o22ai_1 _4562_ (.A1(_2115_),
    .A2(_2179_),
    .B1(_2180_),
    .B2(_2143_),
    .Y(_2181_));
 sky130_fd_sc_hd__a211oi_2 _4563_ (.A1(_2112_),
    .A2(_2178_),
    .B1(_2181_),
    .C1(_2119_),
    .Y(_2182_));
 sky130_fd_sc_hd__mux4_1 _4564_ (.A0(\rf_reg[798] ),
    .A1(\rf_reg[830] ),
    .A2(\rf_reg[926] ),
    .A3(\rf_reg[958] ),
    .S0(_2080_),
    .S1(_1678_),
    .X(_2183_));
 sky130_fd_sc_hd__mux4_1 _4565_ (.A0(\rf_reg[542] ),
    .A1(\rf_reg[574] ),
    .A2(\rf_reg[670] ),
    .A3(\rf_reg[702] ),
    .S0(_1721_),
    .S1(_2060_),
    .X(_2184_));
 sky130_fd_sc_hd__a22o_1 _4566_ (.A1(_2146_),
    .A2(_2183_),
    .B1(_2184_),
    .B2(_2123_),
    .X(_2185_));
 sky130_fd_sc_hd__mux4_1 _4567_ (.A0(\rf_reg[862] ),
    .A1(\rf_reg[894] ),
    .A2(\rf_reg[990] ),
    .A3(\rf_reg[1022] ),
    .S0(_2125_),
    .S1(_2007_),
    .X(_2186_));
 sky130_fd_sc_hd__mux4_1 _4568_ (.A0(\rf_reg[606] ),
    .A1(\rf_reg[638] ),
    .A2(\rf_reg[734] ),
    .A3(\rf_reg[766] ),
    .S0(_2027_),
    .S1(_2104_),
    .X(_2187_));
 sky130_fd_sc_hd__a22o_1 _4569_ (.A1(_2150_),
    .A2(_2186_),
    .B1(_2187_),
    .B2(_2128_),
    .X(_2188_));
 sky130_fd_sc_hd__o21ai_2 _4570_ (.A1(_2185_),
    .A2(_2188_),
    .B1(_2130_),
    .Y(_2189_));
 sky130_fd_sc_hd__o31ai_4 _4571_ (.A1(_2067_),
    .A2(_2176_),
    .A3(_2182_),
    .B1(_2189_),
    .Y(net102));
 sky130_fd_sc_hd__mux4_1 _4572_ (.A0(\rf_reg[287] ),
    .A1(\rf_reg[319] ),
    .A2(\rf_reg[415] ),
    .A3(\rf_reg[447] ),
    .S0(_2012_),
    .S1(_2132_),
    .X(_2190_));
 sky130_fd_sc_hd__mux4_1 _4573_ (.A0(\rf_reg[351] ),
    .A1(\rf_reg[383] ),
    .A2(\rf_reg[479] ),
    .A3(\rf_reg[511] ),
    .S0(_1827_),
    .S1(_2089_),
    .X(_2191_));
 sky130_fd_sc_hd__mux2i_2 _4574_ (.A0(_2190_),
    .A1(_2191_),
    .S(_2091_),
    .Y(_2192_));
 sky130_fd_sc_hd__and2_0 _4575_ (.A(_2068_),
    .B(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__mux2_1 _4576_ (.A0(\rf_reg[63] ),
    .A1(\rf_reg[127] ),
    .S(_2159_),
    .X(_2194_));
 sky130_fd_sc_hd__a22o_1 _4577_ (.A1(\rf_reg[95] ),
    .A2(_2137_),
    .B1(_2194_),
    .B2(_2139_),
    .X(_2195_));
 sky130_fd_sc_hd__mux2i_1 _4578_ (.A0(\rf_reg[223] ),
    .A1(\rf_reg[255] ),
    .S(_2037_),
    .Y(_2196_));
 sky130_fd_sc_hd__mux2i_1 _4579_ (.A0(\rf_reg[159] ),
    .A1(\rf_reg[191] ),
    .S(_2076_),
    .Y(_2197_));
 sky130_fd_sc_hd__o22ai_1 _4580_ (.A1(_2115_),
    .A2(_2196_),
    .B1(_2197_),
    .B2(_2143_),
    .Y(_2198_));
 sky130_fd_sc_hd__a211oi_2 _4581_ (.A1(_2112_),
    .A2(_2195_),
    .B1(_2198_),
    .C1(_2119_),
    .Y(_2199_));
 sky130_fd_sc_hd__mux4_1 _4582_ (.A0(\rf_reg[799] ),
    .A1(\rf_reg[831] ),
    .A2(\rf_reg[927] ),
    .A3(\rf_reg[959] ),
    .S0(_2080_),
    .S1(_1678_),
    .X(_2200_));
 sky130_fd_sc_hd__mux4_1 _4583_ (.A0(\rf_reg[543] ),
    .A1(\rf_reg[575] ),
    .A2(\rf_reg[671] ),
    .A3(\rf_reg[703] ),
    .S0(_1721_),
    .S1(_2060_),
    .X(_2201_));
 sky130_fd_sc_hd__a22o_1 _4584_ (.A1(_2146_),
    .A2(_2200_),
    .B1(_2201_),
    .B2(_2123_),
    .X(_2202_));
 sky130_fd_sc_hd__mux4_1 _4585_ (.A0(\rf_reg[863] ),
    .A1(\rf_reg[895] ),
    .A2(\rf_reg[991] ),
    .A3(\rf_reg[1023] ),
    .S0(_2125_),
    .S1(_1747_),
    .X(_2203_));
 sky130_fd_sc_hd__mux4_1 _4586_ (.A0(\rf_reg[607] ),
    .A1(\rf_reg[639] ),
    .A2(\rf_reg[735] ),
    .A3(\rf_reg[767] ),
    .S0(_2027_),
    .S1(_2104_),
    .X(_2204_));
 sky130_fd_sc_hd__a22o_1 _4587_ (.A1(_2150_),
    .A2(_2203_),
    .B1(_2204_),
    .B2(_2128_),
    .X(_2205_));
 sky130_fd_sc_hd__o21ai_2 _4588_ (.A1(_2202_),
    .A2(_2205_),
    .B1(_2130_),
    .Y(_2206_));
 sky130_fd_sc_hd__o31ai_4 _4589_ (.A1(_2067_),
    .A2(_2193_),
    .A3(_2199_),
    .B1(_2206_),
    .Y(net103));
 sky130_fd_sc_hd__mux4_1 _4590_ (.A0(\rf_reg[259] ),
    .A1(\rf_reg[291] ),
    .A2(\rf_reg[387] ),
    .A3(\rf_reg[419] ),
    .S0(_1680_),
    .S1(_2132_),
    .X(_2207_));
 sky130_fd_sc_hd__mux4_1 _4591_ (.A0(\rf_reg[323] ),
    .A1(\rf_reg[355] ),
    .A2(\rf_reg[451] ),
    .A3(\rf_reg[483] ),
    .S0(_1827_),
    .S1(_2089_),
    .X(_2208_));
 sky130_fd_sc_hd__mux2i_1 _4592_ (.A0(_2207_),
    .A1(_2208_),
    .S(_2091_),
    .Y(_2209_));
 sky130_fd_sc_hd__and2_0 _4593_ (.A(_2068_),
    .B(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__mux2_1 _4594_ (.A0(\rf_reg[35] ),
    .A1(\rf_reg[99] ),
    .S(_2159_),
    .X(_2211_));
 sky130_fd_sc_hd__a22o_1 _4595_ (.A1(\rf_reg[67] ),
    .A2(_2137_),
    .B1(_2211_),
    .B2(_2139_),
    .X(_2212_));
 sky130_fd_sc_hd__mux2i_1 _4596_ (.A0(\rf_reg[195] ),
    .A1(\rf_reg[227] ),
    .S(_2037_),
    .Y(_2213_));
 sky130_fd_sc_hd__mux2i_1 _4597_ (.A0(\rf_reg[131] ),
    .A1(\rf_reg[163] ),
    .S(_2076_),
    .Y(_2214_));
 sky130_fd_sc_hd__o22ai_1 _4598_ (.A1(_2115_),
    .A2(_2213_),
    .B1(_2214_),
    .B2(_2143_),
    .Y(_2215_));
 sky130_fd_sc_hd__a211oi_2 _4599_ (.A1(_2112_),
    .A2(_2212_),
    .B1(_2215_),
    .C1(_2119_),
    .Y(_2216_));
 sky130_fd_sc_hd__mux4_1 _4600_ (.A0(\rf_reg[771] ),
    .A1(\rf_reg[803] ),
    .A2(\rf_reg[899] ),
    .A3(\rf_reg[931] ),
    .S0(_2080_),
    .S1(_1678_),
    .X(_2217_));
 sky130_fd_sc_hd__mux4_1 _4601_ (.A0(\rf_reg[515] ),
    .A1(\rf_reg[547] ),
    .A2(\rf_reg[643] ),
    .A3(\rf_reg[675] ),
    .S0(_1721_),
    .S1(_2060_),
    .X(_2218_));
 sky130_fd_sc_hd__a22o_1 _4602_ (.A1(_2146_),
    .A2(_2217_),
    .B1(_2218_),
    .B2(_2123_),
    .X(_2219_));
 sky130_fd_sc_hd__mux4_1 _4603_ (.A0(\rf_reg[835] ),
    .A1(\rf_reg[867] ),
    .A2(\rf_reg[963] ),
    .A3(\rf_reg[995] ),
    .S0(_2125_),
    .S1(_1747_),
    .X(_2220_));
 sky130_fd_sc_hd__mux4_1 _4604_ (.A0(\rf_reg[579] ),
    .A1(\rf_reg[611] ),
    .A2(\rf_reg[707] ),
    .A3(\rf_reg[739] ),
    .S0(_1715_),
    .S1(_2104_),
    .X(_2221_));
 sky130_fd_sc_hd__a22o_1 _4605_ (.A1(_2150_),
    .A2(_2220_),
    .B1(_2221_),
    .B2(_2128_),
    .X(_2222_));
 sky130_fd_sc_hd__o21ai_2 _4606_ (.A1(_2219_),
    .A2(_2222_),
    .B1(_2130_),
    .Y(_2223_));
 sky130_fd_sc_hd__o31ai_4 _4607_ (.A1(_2067_),
    .A2(_2210_),
    .A3(_2216_),
    .B1(_2223_),
    .Y(net104));
 sky130_fd_sc_hd__mux4_1 _4608_ (.A0(\rf_reg[260] ),
    .A1(\rf_reg[292] ),
    .A2(\rf_reg[388] ),
    .A3(\rf_reg[420] ),
    .S0(_1680_),
    .S1(_2132_),
    .X(_2224_));
 sky130_fd_sc_hd__mux4_1 _4609_ (.A0(\rf_reg[324] ),
    .A1(\rf_reg[356] ),
    .A2(\rf_reg[452] ),
    .A3(\rf_reg[484] ),
    .S0(_1827_),
    .S1(_2089_),
    .X(_2225_));
 sky130_fd_sc_hd__mux2i_1 _4610_ (.A0(_2224_),
    .A1(_2225_),
    .S(_2091_),
    .Y(_2226_));
 sky130_fd_sc_hd__and2_0 _4611_ (.A(_2068_),
    .B(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__mux2_1 _4612_ (.A0(\rf_reg[36] ),
    .A1(\rf_reg[100] ),
    .S(_2159_),
    .X(_2228_));
 sky130_fd_sc_hd__a22o_1 _4613_ (.A1(\rf_reg[68] ),
    .A2(_2137_),
    .B1(_2228_),
    .B2(_2139_),
    .X(_2229_));
 sky130_fd_sc_hd__mux2i_1 _4614_ (.A0(\rf_reg[196] ),
    .A1(\rf_reg[228] ),
    .S(_1696_),
    .Y(_2230_));
 sky130_fd_sc_hd__mux2i_1 _4615_ (.A0(\rf_reg[132] ),
    .A1(\rf_reg[164] ),
    .S(_2076_),
    .Y(_2231_));
 sky130_fd_sc_hd__o22ai_2 _4616_ (.A1(_2115_),
    .A2(_2230_),
    .B1(_2231_),
    .B2(_2143_),
    .Y(_2232_));
 sky130_fd_sc_hd__a211oi_2 _4617_ (.A1(_2112_),
    .A2(_2229_),
    .B1(_2232_),
    .C1(_2119_),
    .Y(_2233_));
 sky130_fd_sc_hd__mux4_1 _4618_ (.A0(\rf_reg[772] ),
    .A1(\rf_reg[804] ),
    .A2(\rf_reg[900] ),
    .A3(\rf_reg[932] ),
    .S0(_2080_),
    .S1(_1678_),
    .X(_2234_));
 sky130_fd_sc_hd__mux4_1 _4619_ (.A0(\rf_reg[516] ),
    .A1(\rf_reg[548] ),
    .A2(\rf_reg[644] ),
    .A3(\rf_reg[676] ),
    .S0(_1721_),
    .S1(_2060_),
    .X(_2235_));
 sky130_fd_sc_hd__a22o_1 _4620_ (.A1(_2146_),
    .A2(_2234_),
    .B1(_2235_),
    .B2(_2123_),
    .X(_2236_));
 sky130_fd_sc_hd__mux4_1 _4621_ (.A0(\rf_reg[836] ),
    .A1(\rf_reg[868] ),
    .A2(\rf_reg[964] ),
    .A3(\rf_reg[996] ),
    .S0(_2125_),
    .S1(_1747_),
    .X(_2237_));
 sky130_fd_sc_hd__mux4_1 _4622_ (.A0(\rf_reg[580] ),
    .A1(\rf_reg[612] ),
    .A2(\rf_reg[708] ),
    .A3(\rf_reg[740] ),
    .S0(_1715_),
    .S1(_2104_),
    .X(_2238_));
 sky130_fd_sc_hd__a22o_1 _4623_ (.A1(_2150_),
    .A2(_2237_),
    .B1(_2238_),
    .B2(_2128_),
    .X(_2239_));
 sky130_fd_sc_hd__o21ai_2 _4624_ (.A1(_2236_),
    .A2(_2239_),
    .B1(_2130_),
    .Y(_2240_));
 sky130_fd_sc_hd__o31ai_4 _4625_ (.A1(_2067_),
    .A2(_2227_),
    .A3(_2233_),
    .B1(_2240_),
    .Y(net105));
 sky130_fd_sc_hd__mux4_1 _4626_ (.A0(\rf_reg[261] ),
    .A1(\rf_reg[293] ),
    .A2(\rf_reg[389] ),
    .A3(\rf_reg[421] ),
    .S0(_1680_),
    .S1(_2132_),
    .X(_2241_));
 sky130_fd_sc_hd__mux4_1 _4627_ (.A0(\rf_reg[325] ),
    .A1(\rf_reg[357] ),
    .A2(\rf_reg[453] ),
    .A3(\rf_reg[485] ),
    .S0(_1827_),
    .S1(_2089_),
    .X(_2242_));
 sky130_fd_sc_hd__mux2i_1 _4628_ (.A0(_2241_),
    .A1(_2242_),
    .S(_2091_),
    .Y(_2243_));
 sky130_fd_sc_hd__and2_0 _4629_ (.A(_2068_),
    .B(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(\rf_reg[37] ),
    .A1(\rf_reg[101] ),
    .S(_2159_),
    .X(_2245_));
 sky130_fd_sc_hd__a22o_1 _4631_ (.A1(\rf_reg[69] ),
    .A2(_2137_),
    .B1(_2245_),
    .B2(_2139_),
    .X(_2246_));
 sky130_fd_sc_hd__mux2i_1 _4632_ (.A0(\rf_reg[197] ),
    .A1(\rf_reg[229] ),
    .S(_1696_),
    .Y(_2247_));
 sky130_fd_sc_hd__mux2i_1 _4633_ (.A0(\rf_reg[133] ),
    .A1(\rf_reg[165] ),
    .S(_2076_),
    .Y(_2248_));
 sky130_fd_sc_hd__o22ai_1 _4634_ (.A1(_2115_),
    .A2(_2247_),
    .B1(_2248_),
    .B2(_2143_),
    .Y(_2249_));
 sky130_fd_sc_hd__a211oi_2 _4635_ (.A1(_2112_),
    .A2(_2246_),
    .B1(_2249_),
    .C1(_2119_),
    .Y(_2250_));
 sky130_fd_sc_hd__mux4_1 _4636_ (.A0(\rf_reg[773] ),
    .A1(\rf_reg[805] ),
    .A2(\rf_reg[901] ),
    .A3(\rf_reg[933] ),
    .S0(_2080_),
    .S1(_1678_),
    .X(_2251_));
 sky130_fd_sc_hd__mux4_1 _4637_ (.A0(\rf_reg[517] ),
    .A1(\rf_reg[549] ),
    .A2(\rf_reg[645] ),
    .A3(\rf_reg[677] ),
    .S0(_1721_),
    .S1(_1711_),
    .X(_2252_));
 sky130_fd_sc_hd__a22o_1 _4638_ (.A1(_2146_),
    .A2(_2251_),
    .B1(_2252_),
    .B2(_2123_),
    .X(_2253_));
 sky130_fd_sc_hd__mux4_1 _4639_ (.A0(\rf_reg[837] ),
    .A1(\rf_reg[869] ),
    .A2(\rf_reg[965] ),
    .A3(\rf_reg[997] ),
    .S0(_2125_),
    .S1(_1747_),
    .X(_2254_));
 sky130_fd_sc_hd__mux4_1 _4640_ (.A0(\rf_reg[581] ),
    .A1(\rf_reg[613] ),
    .A2(\rf_reg[709] ),
    .A3(\rf_reg[741] ),
    .S0(_1715_),
    .S1(_2104_),
    .X(_2255_));
 sky130_fd_sc_hd__a22o_1 _4641_ (.A1(_2150_),
    .A2(_2254_),
    .B1(_2255_),
    .B2(_2128_),
    .X(_2256_));
 sky130_fd_sc_hd__o21ai_2 _4642_ (.A1(_2253_),
    .A2(_2256_),
    .B1(_2130_),
    .Y(_2257_));
 sky130_fd_sc_hd__o31ai_4 _4643_ (.A1(_2067_),
    .A2(_2244_),
    .A3(_2250_),
    .B1(_2257_),
    .Y(net106));
 sky130_fd_sc_hd__mux4_1 _4644_ (.A0(\rf_reg[262] ),
    .A1(\rf_reg[294] ),
    .A2(\rf_reg[390] ),
    .A3(\rf_reg[422] ),
    .S0(_1680_),
    .S1(_2132_),
    .X(_2258_));
 sky130_fd_sc_hd__mux4_1 _4645_ (.A0(\rf_reg[326] ),
    .A1(\rf_reg[358] ),
    .A2(\rf_reg[454] ),
    .A3(\rf_reg[486] ),
    .S0(_1827_),
    .S1(_2089_),
    .X(_2259_));
 sky130_fd_sc_hd__mux2i_1 _4646_ (.A0(_2258_),
    .A1(_2259_),
    .S(_2091_),
    .Y(_2260_));
 sky130_fd_sc_hd__and2_0 _4647_ (.A(_1672_),
    .B(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(\rf_reg[38] ),
    .A1(\rf_reg[102] ),
    .S(_2159_),
    .X(_2262_));
 sky130_fd_sc_hd__a22o_1 _4649_ (.A1(\rf_reg[70] ),
    .A2(_2137_),
    .B1(_2262_),
    .B2(_2139_),
    .X(_2263_));
 sky130_fd_sc_hd__mux2i_1 _4650_ (.A0(\rf_reg[198] ),
    .A1(\rf_reg[230] ),
    .S(_1696_),
    .Y(_2264_));
 sky130_fd_sc_hd__mux2i_1 _4651_ (.A0(\rf_reg[134] ),
    .A1(\rf_reg[166] ),
    .S(_1702_),
    .Y(_2265_));
 sky130_fd_sc_hd__o22ai_1 _4652_ (.A1(_2115_),
    .A2(_2264_),
    .B1(_2265_),
    .B2(_2143_),
    .Y(_2266_));
 sky130_fd_sc_hd__a211oi_2 _4653_ (.A1(_2112_),
    .A2(_2263_),
    .B1(_2266_),
    .C1(_2119_),
    .Y(_2267_));
 sky130_fd_sc_hd__mux4_1 _4654_ (.A0(\rf_reg[774] ),
    .A1(\rf_reg[806] ),
    .A2(\rf_reg[902] ),
    .A3(\rf_reg[934] ),
    .S0(_1675_),
    .S1(_1678_),
    .X(_2268_));
 sky130_fd_sc_hd__mux4_1 _4655_ (.A0(\rf_reg[518] ),
    .A1(\rf_reg[550] ),
    .A2(\rf_reg[646] ),
    .A3(\rf_reg[678] ),
    .S0(_1721_),
    .S1(_1711_),
    .X(_2269_));
 sky130_fd_sc_hd__a22o_1 _4656_ (.A1(_2146_),
    .A2(_2268_),
    .B1(_2269_),
    .B2(_2123_),
    .X(_2270_));
 sky130_fd_sc_hd__mux4_1 _4657_ (.A0(\rf_reg[838] ),
    .A1(\rf_reg[870] ),
    .A2(\rf_reg[966] ),
    .A3(\rf_reg[998] ),
    .S0(_2125_),
    .S1(_1747_),
    .X(_2271_));
 sky130_fd_sc_hd__mux4_1 _4658_ (.A0(\rf_reg[582] ),
    .A1(\rf_reg[614] ),
    .A2(\rf_reg[710] ),
    .A3(\rf_reg[742] ),
    .S0(_1715_),
    .S1(_2104_),
    .X(_2272_));
 sky130_fd_sc_hd__a22o_1 _4659_ (.A1(_2150_),
    .A2(_2271_),
    .B1(_2272_),
    .B2(_2128_),
    .X(_2273_));
 sky130_fd_sc_hd__o21ai_2 _4660_ (.A1(_2270_),
    .A2(_2273_),
    .B1(_2130_),
    .Y(_2274_));
 sky130_fd_sc_hd__o31ai_4 _4661_ (.A1(_1670_),
    .A2(_2261_),
    .A3(_2267_),
    .B1(_2274_),
    .Y(net107));
 sky130_fd_sc_hd__mux4_1 _4662_ (.A0(\rf_reg[263] ),
    .A1(\rf_reg[295] ),
    .A2(\rf_reg[391] ),
    .A3(\rf_reg[423] ),
    .S0(_1680_),
    .S1(_2132_),
    .X(_2275_));
 sky130_fd_sc_hd__mux4_1 _4663_ (.A0(\rf_reg[327] ),
    .A1(\rf_reg[359] ),
    .A2(\rf_reg[455] ),
    .A3(\rf_reg[487] ),
    .S0(_1827_),
    .S1(_1688_),
    .X(_2276_));
 sky130_fd_sc_hd__mux2i_1 _4664_ (.A0(_2275_),
    .A1(_2276_),
    .S(_1684_),
    .Y(_2277_));
 sky130_fd_sc_hd__and2_0 _4665_ (.A(_1672_),
    .B(_2277_),
    .X(_2278_));
 sky130_fd_sc_hd__mux2_1 _4666_ (.A0(\rf_reg[39] ),
    .A1(\rf_reg[103] ),
    .S(_2159_),
    .X(_2279_));
 sky130_fd_sc_hd__a22o_1 _4667_ (.A1(\rf_reg[71] ),
    .A2(_2137_),
    .B1(_2279_),
    .B2(_2139_),
    .X(_2280_));
 sky130_fd_sc_hd__mux2i_1 _4668_ (.A0(\rf_reg[199] ),
    .A1(\rf_reg[231] ),
    .S(_1696_),
    .Y(_2281_));
 sky130_fd_sc_hd__mux2i_1 _4669_ (.A0(\rf_reg[135] ),
    .A1(\rf_reg[167] ),
    .S(_1702_),
    .Y(_2282_));
 sky130_fd_sc_hd__o22ai_1 _4670_ (.A1(_2115_),
    .A2(_2281_),
    .B1(_2282_),
    .B2(_2143_),
    .Y(_2283_));
 sky130_fd_sc_hd__a211oi_2 _4671_ (.A1(_2112_),
    .A2(_2280_),
    .B1(_2283_),
    .C1(_2119_),
    .Y(_2284_));
 sky130_fd_sc_hd__mux4_1 _4672_ (.A0(\rf_reg[775] ),
    .A1(\rf_reg[807] ),
    .A2(\rf_reg[903] ),
    .A3(\rf_reg[935] ),
    .S0(_1675_),
    .S1(_1678_),
    .X(_2285_));
 sky130_fd_sc_hd__mux4_1 _4673_ (.A0(\rf_reg[519] ),
    .A1(\rf_reg[551] ),
    .A2(\rf_reg[647] ),
    .A3(\rf_reg[679] ),
    .S0(_1721_),
    .S1(_1711_),
    .X(_2286_));
 sky130_fd_sc_hd__a22o_1 _4674_ (.A1(_2146_),
    .A2(_2285_),
    .B1(_2286_),
    .B2(_2123_),
    .X(_2287_));
 sky130_fd_sc_hd__mux4_1 _4675_ (.A0(\rf_reg[839] ),
    .A1(\rf_reg[871] ),
    .A2(\rf_reg[967] ),
    .A3(\rf_reg[999] ),
    .S0(_2125_),
    .S1(_1747_),
    .X(_2288_));
 sky130_fd_sc_hd__mux4_1 _4676_ (.A0(\rf_reg[583] ),
    .A1(\rf_reg[615] ),
    .A2(\rf_reg[711] ),
    .A3(\rf_reg[743] ),
    .S0(_1715_),
    .S1(_1716_),
    .X(_2289_));
 sky130_fd_sc_hd__a22o_1 _4677_ (.A1(_2150_),
    .A2(_2288_),
    .B1(_2289_),
    .B2(_2128_),
    .X(_2290_));
 sky130_fd_sc_hd__o21ai_2 _4678_ (.A1(_2287_),
    .A2(_2290_),
    .B1(_2130_),
    .Y(_2291_));
 sky130_fd_sc_hd__o31ai_4 _4679_ (.A1(_1670_),
    .A2(_2278_),
    .A3(_2284_),
    .B1(_2291_),
    .Y(net108));
 sky130_fd_sc_hd__mux4_1 _4680_ (.A0(\rf_reg[264] ),
    .A1(\rf_reg[296] ),
    .A2(\rf_reg[392] ),
    .A3(\rf_reg[424] ),
    .S0(_1680_),
    .S1(_2132_),
    .X(_2292_));
 sky130_fd_sc_hd__mux4_1 _4681_ (.A0(\rf_reg[328] ),
    .A1(\rf_reg[360] ),
    .A2(\rf_reg[456] ),
    .A3(\rf_reg[488] ),
    .S0(_1827_),
    .S1(_1688_),
    .X(_2293_));
 sky130_fd_sc_hd__mux2i_1 _4682_ (.A0(_2292_),
    .A1(_2293_),
    .S(_1684_),
    .Y(_2294_));
 sky130_fd_sc_hd__and2_0 _4683_ (.A(_1672_),
    .B(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__mux2_1 _4684_ (.A0(\rf_reg[40] ),
    .A1(\rf_reg[104] ),
    .S(_2159_),
    .X(_2296_));
 sky130_fd_sc_hd__a22o_1 _4685_ (.A1(\rf_reg[72] ),
    .A2(_2137_),
    .B1(_2296_),
    .B2(_2139_),
    .X(_2297_));
 sky130_fd_sc_hd__mux2i_1 _4686_ (.A0(\rf_reg[200] ),
    .A1(\rf_reg[232] ),
    .S(_1696_),
    .Y(_2298_));
 sky130_fd_sc_hd__mux2i_1 _4687_ (.A0(\rf_reg[136] ),
    .A1(\rf_reg[168] ),
    .S(_1702_),
    .Y(_2299_));
 sky130_fd_sc_hd__o22ai_1 _4688_ (.A1(_1699_),
    .A2(_2298_),
    .B1(_2299_),
    .B2(_2143_),
    .Y(_2300_));
 sky130_fd_sc_hd__a211oi_2 _4689_ (.A1(_1690_),
    .A2(_2297_),
    .B1(_2300_),
    .C1(_1673_),
    .Y(_2301_));
 sky130_fd_sc_hd__mux4_1 _4690_ (.A0(\rf_reg[776] ),
    .A1(\rf_reg[808] ),
    .A2(\rf_reg[904] ),
    .A3(\rf_reg[936] ),
    .S0(_1675_),
    .S1(_1678_),
    .X(_2302_));
 sky130_fd_sc_hd__mux4_1 _4691_ (.A0(\rf_reg[520] ),
    .A1(\rf_reg[552] ),
    .A2(\rf_reg[648] ),
    .A3(\rf_reg[680] ),
    .S0(_1721_),
    .S1(_1711_),
    .X(_2303_));
 sky130_fd_sc_hd__a22o_1 _4692_ (.A1(_2146_),
    .A2(_2302_),
    .B1(_2303_),
    .B2(_1718_),
    .X(_2304_));
 sky130_fd_sc_hd__mux4_1 _4693_ (.A0(\rf_reg[840] ),
    .A1(\rf_reg[872] ),
    .A2(\rf_reg[968] ),
    .A3(\rf_reg[1000] ),
    .S0(_1695_),
    .S1(_1747_),
    .X(_2305_));
 sky130_fd_sc_hd__mux4_1 _4694_ (.A0(\rf_reg[584] ),
    .A1(\rf_reg[616] ),
    .A2(\rf_reg[712] ),
    .A3(\rf_reg[744] ),
    .S0(_1715_),
    .S1(_1716_),
    .X(_2306_));
 sky130_fd_sc_hd__a22o_1 _4695_ (.A1(_2150_),
    .A2(_2305_),
    .B1(_2306_),
    .B2(_1727_),
    .X(_2307_));
 sky130_fd_sc_hd__o21ai_2 _4696_ (.A1(_2304_),
    .A2(_2307_),
    .B1(_1671_),
    .Y(_2308_));
 sky130_fd_sc_hd__o31ai_4 _4697_ (.A1(_1670_),
    .A2(_2295_),
    .A3(_2301_),
    .B1(_2308_),
    .Y(net109));
 sky130_fd_sc_hd__mux4_1 _4698_ (.A0(\rf_reg[265] ),
    .A1(\rf_reg[297] ),
    .A2(\rf_reg[393] ),
    .A3(\rf_reg[425] ),
    .S0(_1680_),
    .S1(_1681_),
    .X(_2309_));
 sky130_fd_sc_hd__mux4_1 _4699_ (.A0(\rf_reg[329] ),
    .A1(\rf_reg[361] ),
    .A2(\rf_reg[457] ),
    .A3(\rf_reg[489] ),
    .S0(_1827_),
    .S1(_1688_),
    .X(_2310_));
 sky130_fd_sc_hd__mux2i_1 _4700_ (.A0(_2309_),
    .A1(_2310_),
    .S(_1684_),
    .Y(_2311_));
 sky130_fd_sc_hd__and2_0 _4701_ (.A(_1672_),
    .B(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__mux2_1 _4702_ (.A0(\rf_reg[41] ),
    .A1(\rf_reg[105] ),
    .S(_2159_),
    .X(_2313_));
 sky130_fd_sc_hd__a22o_1 _4703_ (.A1(\rf_reg[73] ),
    .A2(_1738_),
    .B1(_2313_),
    .B2(_1705_),
    .X(_2314_));
 sky130_fd_sc_hd__mux2i_1 _4704_ (.A0(\rf_reg[201] ),
    .A1(\rf_reg[233] ),
    .S(_1696_),
    .Y(_2315_));
 sky130_fd_sc_hd__mux2i_1 _4705_ (.A0(\rf_reg[137] ),
    .A1(\rf_reg[169] ),
    .S(_1702_),
    .Y(_2316_));
 sky130_fd_sc_hd__o22ai_2 _4706_ (.A1(_1699_),
    .A2(_2315_),
    .B1(_2316_),
    .B2(_1704_),
    .Y(_2317_));
 sky130_fd_sc_hd__a211oi_4 _4707_ (.A1(_1690_),
    .A2(_2314_),
    .B1(_2317_),
    .C1(_1673_),
    .Y(_2318_));
 sky130_fd_sc_hd__mux4_1 _4708_ (.A0(\rf_reg[777] ),
    .A1(\rf_reg[809] ),
    .A2(\rf_reg[905] ),
    .A3(\rf_reg[937] ),
    .S0(_1675_),
    .S1(_1678_),
    .X(_2319_));
 sky130_fd_sc_hd__mux4_1 _4709_ (.A0(\rf_reg[521] ),
    .A1(\rf_reg[553] ),
    .A2(\rf_reg[649] ),
    .A3(\rf_reg[681] ),
    .S0(_1721_),
    .S1(_1711_),
    .X(_2320_));
 sky130_fd_sc_hd__a22o_1 _4710_ (.A1(_1714_),
    .A2(_2319_),
    .B1(_2320_),
    .B2(_1718_),
    .X(_2321_));
 sky130_fd_sc_hd__mux4_1 _4711_ (.A0(\rf_reg[841] ),
    .A1(\rf_reg[873] ),
    .A2(\rf_reg[969] ),
    .A3(\rf_reg[1001] ),
    .S0(_1695_),
    .S1(_1747_),
    .X(_2322_));
 sky130_fd_sc_hd__mux4_1 _4712_ (.A0(\rf_reg[585] ),
    .A1(\rf_reg[617] ),
    .A2(\rf_reg[713] ),
    .A3(\rf_reg[745] ),
    .S0(_1715_),
    .S1(_1716_),
    .X(_2323_));
 sky130_fd_sc_hd__a22o_1 _4713_ (.A1(_1724_),
    .A2(_2322_),
    .B1(_2323_),
    .B2(_1727_),
    .X(_2324_));
 sky130_fd_sc_hd__o21ai_2 _4714_ (.A1(_2321_),
    .A2(_2324_),
    .B1(_1671_),
    .Y(_2325_));
 sky130_fd_sc_hd__o31ai_4 _4715_ (.A1(_1670_),
    .A2(_2312_),
    .A3(_2318_),
    .B1(_2325_),
    .Y(net110));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[0]$_DFFE_PN0P_  (.D(_0000_),
    .Q(\rf_reg[32] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[100]$_DFFE_PN0P_  (.D(_0001_),
    .Q(\rf_reg[132] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[101]$_DFFE_PN0P_  (.D(_0002_),
    .Q(\rf_reg[133] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[102]$_DFFE_PN0P_  (.D(_0003_),
    .Q(\rf_reg[134] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[103]$_DFFE_PN0P_  (.D(_0004_),
    .Q(\rf_reg[135] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[104]$_DFFE_PN0P_  (.D(_0005_),
    .Q(\rf_reg[136] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[105]$_DFFE_PN0P_  (.D(_0006_),
    .Q(\rf_reg[137] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[106]$_DFFE_PN0P_  (.D(_0007_),
    .Q(\rf_reg[138] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[107]$_DFFE_PN0P_  (.D(_0008_),
    .Q(\rf_reg[139] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[108]$_DFFE_PN0P_  (.D(_0009_),
    .Q(\rf_reg[140] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[109]$_DFFE_PN0P_  (.D(_0010_),
    .Q(\rf_reg[141] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[10]$_DFFE_PN0P_  (.D(_0011_),
    .Q(\rf_reg[42] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[110]$_DFFE_PN0P_  (.D(_0012_),
    .Q(\rf_reg[142] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[111]$_DFFE_PN0P_  (.D(_0013_),
    .Q(\rf_reg[143] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[112]$_DFFE_PN0P_  (.D(_0014_),
    .Q(\rf_reg[144] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[113]$_DFFE_PN0P_  (.D(_0015_),
    .Q(\rf_reg[145] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[114]$_DFFE_PN0P_  (.D(_0016_),
    .Q(\rf_reg[146] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[115]$_DFFE_PN0P_  (.D(_0017_),
    .Q(\rf_reg[147] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[116]$_DFFE_PN0P_  (.D(_0018_),
    .Q(\rf_reg[148] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[117]$_DFFE_PN0P_  (.D(_0019_),
    .Q(\rf_reg[149] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[118]$_DFFE_PN0P_  (.D(_0020_),
    .Q(\rf_reg[150] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[119]$_DFFE_PN0P_  (.D(_0021_),
    .Q(\rf_reg[151] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[11]$_DFFE_PN0P_  (.D(_0022_),
    .Q(\rf_reg[43] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[120]$_DFFE_PN0P_  (.D(_0023_),
    .Q(\rf_reg[152] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[121]$_DFFE_PN0P_  (.D(_0024_),
    .Q(\rf_reg[153] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[122]$_DFFE_PN0P_  (.D(_0025_),
    .Q(\rf_reg[154] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[123]$_DFFE_PN0P_  (.D(_0026_),
    .Q(\rf_reg[155] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[124]$_DFFE_PN0P_  (.D(_0027_),
    .Q(\rf_reg[156] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[125]$_DFFE_PN0P_  (.D(_0028_),
    .Q(\rf_reg[157] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[126]$_DFFE_PN0P_  (.D(_0029_),
    .Q(\rf_reg[158] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[127]$_DFFE_PN0P_  (.D(_0030_),
    .Q(\rf_reg[159] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[128]$_DFFE_PN0P_  (.D(_0031_),
    .Q(\rf_reg[160] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[129]$_DFFE_PN0P_  (.D(_0032_),
    .Q(\rf_reg[161] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[12]$_DFFE_PN0P_  (.D(_0033_),
    .Q(\rf_reg[44] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[130]$_DFFE_PN0P_  (.D(_0034_),
    .Q(\rf_reg[162] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[131]$_DFFE_PN0P_  (.D(_0035_),
    .Q(\rf_reg[163] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[132]$_DFFE_PN0P_  (.D(_0036_),
    .Q(\rf_reg[164] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[133]$_DFFE_PN0P_  (.D(_0037_),
    .Q(\rf_reg[165] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[134]$_DFFE_PN0P_  (.D(_0038_),
    .Q(\rf_reg[166] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[135]$_DFFE_PN0P_  (.D(_0039_),
    .Q(\rf_reg[167] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[136]$_DFFE_PN0P_  (.D(_0040_),
    .Q(\rf_reg[168] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[137]$_DFFE_PN0P_  (.D(_0041_),
    .Q(\rf_reg[169] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[138]$_DFFE_PN0P_  (.D(_0042_),
    .Q(\rf_reg[170] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[139]$_DFFE_PN0P_  (.D(_0043_),
    .Q(\rf_reg[171] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[13]$_DFFE_PN0P_  (.D(_0044_),
    .Q(\rf_reg[45] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[140]$_DFFE_PN0P_  (.D(_0045_),
    .Q(\rf_reg[172] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[141]$_DFFE_PN0P_  (.D(_0046_),
    .Q(\rf_reg[173] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[142]$_DFFE_PN0P_  (.D(_0047_),
    .Q(\rf_reg[174] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[143]$_DFFE_PN0P_  (.D(_0048_),
    .Q(\rf_reg[175] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[144]$_DFFE_PN0P_  (.D(_0049_),
    .Q(\rf_reg[176] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[145]$_DFFE_PN0P_  (.D(_0050_),
    .Q(\rf_reg[177] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[146]$_DFFE_PN0P_  (.D(_0051_),
    .Q(\rf_reg[178] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[147]$_DFFE_PN0P_  (.D(_0052_),
    .Q(\rf_reg[179] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[148]$_DFFE_PN0P_  (.D(_0053_),
    .Q(\rf_reg[180] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[149]$_DFFE_PN0P_  (.D(_0054_),
    .Q(\rf_reg[181] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[14]$_DFFE_PN0P_  (.D(_0055_),
    .Q(\rf_reg[46] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[150]$_DFFE_PN0P_  (.D(_0056_),
    .Q(\rf_reg[182] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[151]$_DFFE_PN0P_  (.D(_0057_),
    .Q(\rf_reg[183] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[152]$_DFFE_PN0P_  (.D(_0058_),
    .Q(\rf_reg[184] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[153]$_DFFE_PN0P_  (.D(_0059_),
    .Q(\rf_reg[185] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[154]$_DFFE_PN0P_  (.D(_0060_),
    .Q(\rf_reg[186] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[155]$_DFFE_PN0P_  (.D(_0061_),
    .Q(\rf_reg[187] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[156]$_DFFE_PN0P_  (.D(_0062_),
    .Q(\rf_reg[188] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[157]$_DFFE_PN0P_  (.D(_0063_),
    .Q(\rf_reg[189] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[158]$_DFFE_PN0P_  (.D(_0064_),
    .Q(\rf_reg[190] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[159]$_DFFE_PN0P_  (.D(_0065_),
    .Q(\rf_reg[191] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[15]$_DFFE_PN0P_  (.D(_0066_),
    .Q(\rf_reg[47] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[160]$_DFFE_PN0P_  (.D(_0067_),
    .Q(\rf_reg[192] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[161]$_DFFE_PN0P_  (.D(_0068_),
    .Q(\rf_reg[193] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[162]$_DFFE_PN0P_  (.D(_0069_),
    .Q(\rf_reg[194] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[163]$_DFFE_PN0P_  (.D(_0070_),
    .Q(\rf_reg[195] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[164]$_DFFE_PN0P_  (.D(_0071_),
    .Q(\rf_reg[196] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[165]$_DFFE_PN0P_  (.D(_0072_),
    .Q(\rf_reg[197] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[166]$_DFFE_PN0P_  (.D(_0073_),
    .Q(\rf_reg[198] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[167]$_DFFE_PN0P_  (.D(_0074_),
    .Q(\rf_reg[199] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[168]$_DFFE_PN0P_  (.D(_0075_),
    .Q(\rf_reg[200] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[169]$_DFFE_PN0P_  (.D(_0076_),
    .Q(\rf_reg[201] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[16]$_DFFE_PN0P_  (.D(_0077_),
    .Q(\rf_reg[48] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[170]$_DFFE_PN0P_  (.D(_0078_),
    .Q(\rf_reg[202] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[171]$_DFFE_PN0P_  (.D(_0079_),
    .Q(\rf_reg[203] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[172]$_DFFE_PN0P_  (.D(_0080_),
    .Q(\rf_reg[204] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[173]$_DFFE_PN0P_  (.D(_0081_),
    .Q(\rf_reg[205] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[174]$_DFFE_PN0P_  (.D(_0082_),
    .Q(\rf_reg[206] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[175]$_DFFE_PN0P_  (.D(_0083_),
    .Q(\rf_reg[207] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[176]$_DFFE_PN0P_  (.D(_0084_),
    .Q(\rf_reg[208] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[177]$_DFFE_PN0P_  (.D(_0085_),
    .Q(\rf_reg[209] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[178]$_DFFE_PN0P_  (.D(_0086_),
    .Q(\rf_reg[210] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[179]$_DFFE_PN0P_  (.D(_0087_),
    .Q(\rf_reg[211] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[17]$_DFFE_PN0P_  (.D(_0088_),
    .Q(\rf_reg[49] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[180]$_DFFE_PN0P_  (.D(_0089_),
    .Q(\rf_reg[212] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[181]$_DFFE_PN0P_  (.D(_0090_),
    .Q(\rf_reg[213] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[182]$_DFFE_PN0P_  (.D(_0091_),
    .Q(\rf_reg[214] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[183]$_DFFE_PN0P_  (.D(_0092_),
    .Q(\rf_reg[215] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[184]$_DFFE_PN0P_  (.D(_0093_),
    .Q(\rf_reg[216] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[185]$_DFFE_PN0P_  (.D(_0094_),
    .Q(\rf_reg[217] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[186]$_DFFE_PN0P_  (.D(_0095_),
    .Q(\rf_reg[218] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[187]$_DFFE_PN0P_  (.D(_0096_),
    .Q(\rf_reg[219] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[188]$_DFFE_PN0P_  (.D(_0097_),
    .Q(\rf_reg[220] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[189]$_DFFE_PN0P_  (.D(_0098_),
    .Q(\rf_reg[221] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[18]$_DFFE_PN0P_  (.D(_0099_),
    .Q(\rf_reg[50] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[190]$_DFFE_PN0P_  (.D(_0100_),
    .Q(\rf_reg[222] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[191]$_DFFE_PN0P_  (.D(_0101_),
    .Q(\rf_reg[223] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[192]$_DFFE_PN0P_  (.D(_0102_),
    .Q(\rf_reg[224] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[193]$_DFFE_PN0P_  (.D(_0103_),
    .Q(\rf_reg[225] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[194]$_DFFE_PN0P_  (.D(_0104_),
    .Q(\rf_reg[226] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[195]$_DFFE_PN0P_  (.D(_0105_),
    .Q(\rf_reg[227] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[196]$_DFFE_PN0P_  (.D(_0106_),
    .Q(\rf_reg[228] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[197]$_DFFE_PN0P_  (.D(_0107_),
    .Q(\rf_reg[229] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[198]$_DFFE_PN0P_  (.D(_0108_),
    .Q(\rf_reg[230] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[199]$_DFFE_PN0P_  (.D(_0109_),
    .Q(\rf_reg[231] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[19]$_DFFE_PN0P_  (.D(_0110_),
    .Q(\rf_reg[51] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[1]$_DFFE_PN0P_  (.D(_0111_),
    .Q(\rf_reg[33] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[200]$_DFFE_PN0P_  (.D(_0112_),
    .Q(\rf_reg[232] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[201]$_DFFE_PN0P_  (.D(_0113_),
    .Q(\rf_reg[233] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[202]$_DFFE_PN0P_  (.D(_0114_),
    .Q(\rf_reg[234] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[203]$_DFFE_PN0P_  (.D(_0115_),
    .Q(\rf_reg[235] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[204]$_DFFE_PN0P_  (.D(_0116_),
    .Q(\rf_reg[236] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[205]$_DFFE_PN0P_  (.D(_0117_),
    .Q(\rf_reg[237] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[206]$_DFFE_PN0P_  (.D(_0118_),
    .Q(\rf_reg[238] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[207]$_DFFE_PN0P_  (.D(_0119_),
    .Q(\rf_reg[239] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[208]$_DFFE_PN0P_  (.D(_0120_),
    .Q(\rf_reg[240] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[209]$_DFFE_PN0P_  (.D(_0121_),
    .Q(\rf_reg[241] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[20]$_DFFE_PN0P_  (.D(_0122_),
    .Q(\rf_reg[52] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[210]$_DFFE_PN0P_  (.D(_0123_),
    .Q(\rf_reg[242] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[211]$_DFFE_PN0P_  (.D(_0124_),
    .Q(\rf_reg[243] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[212]$_DFFE_PN0P_  (.D(_0125_),
    .Q(\rf_reg[244] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[213]$_DFFE_PN0P_  (.D(_0126_),
    .Q(\rf_reg[245] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[214]$_DFFE_PN0P_  (.D(_0127_),
    .Q(\rf_reg[246] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[215]$_DFFE_PN0P_  (.D(_0128_),
    .Q(\rf_reg[247] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[216]$_DFFE_PN0P_  (.D(_0129_),
    .Q(\rf_reg[248] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[217]$_DFFE_PN0P_  (.D(_0130_),
    .Q(\rf_reg[249] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[218]$_DFFE_PN0P_  (.D(_0131_),
    .Q(\rf_reg[250] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[219]$_DFFE_PN0P_  (.D(_0132_),
    .Q(\rf_reg[251] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[21]$_DFFE_PN0P_  (.D(_0133_),
    .Q(\rf_reg[53] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[220]$_DFFE_PN0P_  (.D(_0134_),
    .Q(\rf_reg[252] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[221]$_DFFE_PN0P_  (.D(_0135_),
    .Q(\rf_reg[253] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[222]$_DFFE_PN0P_  (.D(_0136_),
    .Q(\rf_reg[254] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[223]$_DFFE_PN0P_  (.D(_0137_),
    .Q(\rf_reg[255] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[224]$_DFFE_PN0P_  (.D(_0138_),
    .Q(\rf_reg[256] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[225]$_DFFE_PN0P_  (.D(_0139_),
    .Q(\rf_reg[257] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[226]$_DFFE_PN0P_  (.D(_0140_),
    .Q(\rf_reg[258] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[227]$_DFFE_PN0P_  (.D(_0141_),
    .Q(\rf_reg[259] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[228]$_DFFE_PN0P_  (.D(_0142_),
    .Q(\rf_reg[260] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[229]$_DFFE_PN0P_  (.D(_0143_),
    .Q(\rf_reg[261] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[22]$_DFFE_PN0P_  (.D(_0144_),
    .Q(\rf_reg[54] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[230]$_DFFE_PN0P_  (.D(_0145_),
    .Q(\rf_reg[262] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[231]$_DFFE_PN0P_  (.D(_0146_),
    .Q(\rf_reg[263] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[232]$_DFFE_PN0P_  (.D(_0147_),
    .Q(\rf_reg[264] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[233]$_DFFE_PN0P_  (.D(_0148_),
    .Q(\rf_reg[265] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[234]$_DFFE_PN0P_  (.D(_0149_),
    .Q(\rf_reg[266] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[235]$_DFFE_PN0P_  (.D(_0150_),
    .Q(\rf_reg[267] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[236]$_DFFE_PN0P_  (.D(_0151_),
    .Q(\rf_reg[268] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[237]$_DFFE_PN0P_  (.D(_0152_),
    .Q(\rf_reg[269] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[238]$_DFFE_PN0P_  (.D(_0153_),
    .Q(\rf_reg[270] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[239]$_DFFE_PN0P_  (.D(_0154_),
    .Q(\rf_reg[271] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[23]$_DFFE_PN0P_  (.D(_0155_),
    .Q(\rf_reg[55] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[240]$_DFFE_PN0P_  (.D(_0156_),
    .Q(\rf_reg[272] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[241]$_DFFE_PN0P_  (.D(_0157_),
    .Q(\rf_reg[273] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[242]$_DFFE_PN0P_  (.D(_0158_),
    .Q(\rf_reg[274] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[243]$_DFFE_PN0P_  (.D(_0159_),
    .Q(\rf_reg[275] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[244]$_DFFE_PN0P_  (.D(_0160_),
    .Q(\rf_reg[276] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[245]$_DFFE_PN0P_  (.D(_0161_),
    .Q(\rf_reg[277] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[246]$_DFFE_PN0P_  (.D(_0162_),
    .Q(\rf_reg[278] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[247]$_DFFE_PN0P_  (.D(_0163_),
    .Q(\rf_reg[279] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[248]$_DFFE_PN0P_  (.D(_0164_),
    .Q(\rf_reg[280] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[249]$_DFFE_PN0P_  (.D(_0165_),
    .Q(\rf_reg[281] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[24]$_DFFE_PN0P_  (.D(_0166_),
    .Q(\rf_reg[56] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[250]$_DFFE_PN0P_  (.D(_0167_),
    .Q(\rf_reg[282] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[251]$_DFFE_PN0P_  (.D(_0168_),
    .Q(\rf_reg[283] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[252]$_DFFE_PN0P_  (.D(_0169_),
    .Q(\rf_reg[284] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[253]$_DFFE_PN0P_  (.D(_0170_),
    .Q(\rf_reg[285] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[254]$_DFFE_PN0P_  (.D(_0171_),
    .Q(\rf_reg[286] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[255]$_DFFE_PN0P_  (.D(_0172_),
    .Q(\rf_reg[287] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[256]$_DFFE_PN0P_  (.D(_0173_),
    .Q(\rf_reg[288] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[257]$_DFFE_PN0P_  (.D(_0174_),
    .Q(\rf_reg[289] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[258]$_DFFE_PN0P_  (.D(_0175_),
    .Q(\rf_reg[290] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[259]$_DFFE_PN0P_  (.D(_0176_),
    .Q(\rf_reg[291] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[25]$_DFFE_PN0P_  (.D(_0177_),
    .Q(\rf_reg[57] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[260]$_DFFE_PN0P_  (.D(_0178_),
    .Q(\rf_reg[292] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[261]$_DFFE_PN0P_  (.D(_0179_),
    .Q(\rf_reg[293] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[262]$_DFFE_PN0P_  (.D(_0180_),
    .Q(\rf_reg[294] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[263]$_DFFE_PN0P_  (.D(_0181_),
    .Q(\rf_reg[295] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[264]$_DFFE_PN0P_  (.D(_0182_),
    .Q(\rf_reg[296] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[265]$_DFFE_PN0P_  (.D(_0183_),
    .Q(\rf_reg[297] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[266]$_DFFE_PN0P_  (.D(_0184_),
    .Q(\rf_reg[298] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[267]$_DFFE_PN0P_  (.D(_0185_),
    .Q(\rf_reg[299] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[268]$_DFFE_PN0P_  (.D(_0186_),
    .Q(\rf_reg[300] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[269]$_DFFE_PN0P_  (.D(_0187_),
    .Q(\rf_reg[301] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[26]$_DFFE_PN0P_  (.D(_0188_),
    .Q(\rf_reg[58] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[270]$_DFFE_PN0P_  (.D(_0189_),
    .Q(\rf_reg[302] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[271]$_DFFE_PN0P_  (.D(_0190_),
    .Q(\rf_reg[303] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[272]$_DFFE_PN0P_  (.D(_0191_),
    .Q(\rf_reg[304] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[273]$_DFFE_PN0P_  (.D(_0192_),
    .Q(\rf_reg[305] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[274]$_DFFE_PN0P_  (.D(_0193_),
    .Q(\rf_reg[306] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[275]$_DFFE_PN0P_  (.D(_0194_),
    .Q(\rf_reg[307] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[276]$_DFFE_PN0P_  (.D(_0195_),
    .Q(\rf_reg[308] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[277]$_DFFE_PN0P_  (.D(_0196_),
    .Q(\rf_reg[309] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[278]$_DFFE_PN0P_  (.D(_0197_),
    .Q(\rf_reg[310] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[279]$_DFFE_PN0P_  (.D(_0198_),
    .Q(\rf_reg[311] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[27]$_DFFE_PN0P_  (.D(_0199_),
    .Q(\rf_reg[59] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[280]$_DFFE_PN0P_  (.D(_0200_),
    .Q(\rf_reg[312] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[281]$_DFFE_PN0P_  (.D(_0201_),
    .Q(\rf_reg[313] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[282]$_DFFE_PN0P_  (.D(_0202_),
    .Q(\rf_reg[314] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[283]$_DFFE_PN0P_  (.D(_0203_),
    .Q(\rf_reg[315] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[284]$_DFFE_PN0P_  (.D(_0204_),
    .Q(\rf_reg[316] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[285]$_DFFE_PN0P_  (.D(_0205_),
    .Q(\rf_reg[317] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[286]$_DFFE_PN0P_  (.D(_0206_),
    .Q(\rf_reg[318] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[287]$_DFFE_PN0P_  (.D(_0207_),
    .Q(\rf_reg[319] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[288]$_DFFE_PN0P_  (.D(_0208_),
    .Q(\rf_reg[320] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[289]$_DFFE_PN0P_  (.D(_0209_),
    .Q(\rf_reg[321] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[28]$_DFFE_PN0P_  (.D(_0210_),
    .Q(\rf_reg[60] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[290]$_DFFE_PN0P_  (.D(_0211_),
    .Q(\rf_reg[322] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[291]$_DFFE_PN0P_  (.D(_0212_),
    .Q(\rf_reg[323] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[292]$_DFFE_PN0P_  (.D(_0213_),
    .Q(\rf_reg[324] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[293]$_DFFE_PN0P_  (.D(_0214_),
    .Q(\rf_reg[325] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[294]$_DFFE_PN0P_  (.D(_0215_),
    .Q(\rf_reg[326] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[295]$_DFFE_PN0P_  (.D(_0216_),
    .Q(\rf_reg[327] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[296]$_DFFE_PN0P_  (.D(_0217_),
    .Q(\rf_reg[328] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[297]$_DFFE_PN0P_  (.D(_0218_),
    .Q(\rf_reg[329] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[298]$_DFFE_PN0P_  (.D(_0219_),
    .Q(\rf_reg[330] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[299]$_DFFE_PN0P_  (.D(_0220_),
    .Q(\rf_reg[331] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[29]$_DFFE_PN0P_  (.D(_0221_),
    .Q(\rf_reg[61] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[2]$_DFFE_PN0P_  (.D(_0222_),
    .Q(\rf_reg[34] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[300]$_DFFE_PN0P_  (.D(_0223_),
    .Q(\rf_reg[332] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[301]$_DFFE_PN0P_  (.D(_0224_),
    .Q(\rf_reg[333] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[302]$_DFFE_PN0P_  (.D(_0225_),
    .Q(\rf_reg[334] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[303]$_DFFE_PN0P_  (.D(_0226_),
    .Q(\rf_reg[335] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[304]$_DFFE_PN0P_  (.D(_0227_),
    .Q(\rf_reg[336] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[305]$_DFFE_PN0P_  (.D(_0228_),
    .Q(\rf_reg[337] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[306]$_DFFE_PN0P_  (.D(_0229_),
    .Q(\rf_reg[338] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[307]$_DFFE_PN0P_  (.D(_0230_),
    .Q(\rf_reg[339] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[308]$_DFFE_PN0P_  (.D(_0231_),
    .Q(\rf_reg[340] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[309]$_DFFE_PN0P_  (.D(_0232_),
    .Q(\rf_reg[341] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[30]$_DFFE_PN0P_  (.D(_0233_),
    .Q(\rf_reg[62] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[310]$_DFFE_PN0P_  (.D(_0234_),
    .Q(\rf_reg[342] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[311]$_DFFE_PN0P_  (.D(_0235_),
    .Q(\rf_reg[343] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[312]$_DFFE_PN0P_  (.D(_0236_),
    .Q(\rf_reg[344] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[313]$_DFFE_PN0P_  (.D(_0237_),
    .Q(\rf_reg[345] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[314]$_DFFE_PN0P_  (.D(_0238_),
    .Q(\rf_reg[346] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[315]$_DFFE_PN0P_  (.D(_0239_),
    .Q(\rf_reg[347] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[316]$_DFFE_PN0P_  (.D(_0240_),
    .Q(\rf_reg[348] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[317]$_DFFE_PN0P_  (.D(_0241_),
    .Q(\rf_reg[349] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[318]$_DFFE_PN0P_  (.D(_0242_),
    .Q(\rf_reg[350] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[319]$_DFFE_PN0P_  (.D(_0243_),
    .Q(\rf_reg[351] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[31]$_DFFE_PN0P_  (.D(_0244_),
    .Q(\rf_reg[63] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[320]$_DFFE_PN0P_  (.D(_0245_),
    .Q(\rf_reg[352] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[321]$_DFFE_PN0P_  (.D(_0246_),
    .Q(\rf_reg[353] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[322]$_DFFE_PN0P_  (.D(_0247_),
    .Q(\rf_reg[354] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[323]$_DFFE_PN0P_  (.D(_0248_),
    .Q(\rf_reg[355] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[324]$_DFFE_PN0P_  (.D(_0249_),
    .Q(\rf_reg[356] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[325]$_DFFE_PN0P_  (.D(_0250_),
    .Q(\rf_reg[357] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[326]$_DFFE_PN0P_  (.D(_0251_),
    .Q(\rf_reg[358] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[327]$_DFFE_PN0P_  (.D(_0252_),
    .Q(\rf_reg[359] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[328]$_DFFE_PN0P_  (.D(_0253_),
    .Q(\rf_reg[360] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[329]$_DFFE_PN0P_  (.D(_0254_),
    .Q(\rf_reg[361] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[32]$_DFFE_PN0P_  (.D(_0255_),
    .Q(\rf_reg[64] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[330]$_DFFE_PN0P_  (.D(_0256_),
    .Q(\rf_reg[362] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[331]$_DFFE_PN0P_  (.D(_0257_),
    .Q(\rf_reg[363] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[332]$_DFFE_PN0P_  (.D(_0258_),
    .Q(\rf_reg[364] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[333]$_DFFE_PN0P_  (.D(_0259_),
    .Q(\rf_reg[365] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[334]$_DFFE_PN0P_  (.D(_0260_),
    .Q(\rf_reg[366] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[335]$_DFFE_PN0P_  (.D(_0261_),
    .Q(\rf_reg[367] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[336]$_DFFE_PN0P_  (.D(_0262_),
    .Q(\rf_reg[368] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[337]$_DFFE_PN0P_  (.D(_0263_),
    .Q(\rf_reg[369] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[338]$_DFFE_PN0P_  (.D(_0264_),
    .Q(\rf_reg[370] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[339]$_DFFE_PN0P_  (.D(_0265_),
    .Q(\rf_reg[371] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[33]$_DFFE_PN0P_  (.D(_0266_),
    .Q(\rf_reg[65] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[340]$_DFFE_PN0P_  (.D(_0267_),
    .Q(\rf_reg[372] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[341]$_DFFE_PN0P_  (.D(_0268_),
    .Q(\rf_reg[373] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[342]$_DFFE_PN0P_  (.D(_0269_),
    .Q(\rf_reg[374] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[343]$_DFFE_PN0P_  (.D(_0270_),
    .Q(\rf_reg[375] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[344]$_DFFE_PN0P_  (.D(_0271_),
    .Q(\rf_reg[376] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[345]$_DFFE_PN0P_  (.D(_0272_),
    .Q(\rf_reg[377] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[346]$_DFFE_PN0P_  (.D(_0273_),
    .Q(\rf_reg[378] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[347]$_DFFE_PN0P_  (.D(_0274_),
    .Q(\rf_reg[379] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[348]$_DFFE_PN0P_  (.D(_0275_),
    .Q(\rf_reg[380] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[349]$_DFFE_PN0P_  (.D(_0276_),
    .Q(\rf_reg[381] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[34]$_DFFE_PN0P_  (.D(_0277_),
    .Q(\rf_reg[66] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[350]$_DFFE_PN0P_  (.D(_0278_),
    .Q(\rf_reg[382] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[351]$_DFFE_PN0P_  (.D(_0279_),
    .Q(\rf_reg[383] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[352]$_DFFE_PN0P_  (.D(_0280_),
    .Q(\rf_reg[384] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[353]$_DFFE_PN0P_  (.D(_0281_),
    .Q(\rf_reg[385] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[354]$_DFFE_PN0P_  (.D(_0282_),
    .Q(\rf_reg[386] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[355]$_DFFE_PN0P_  (.D(_0283_),
    .Q(\rf_reg[387] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[356]$_DFFE_PN0P_  (.D(_0284_),
    .Q(\rf_reg[388] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[357]$_DFFE_PN0P_  (.D(_0285_),
    .Q(\rf_reg[389] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[358]$_DFFE_PN0P_  (.D(_0286_),
    .Q(\rf_reg[390] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[359]$_DFFE_PN0P_  (.D(_0287_),
    .Q(\rf_reg[391] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[35]$_DFFE_PN0P_  (.D(_0288_),
    .Q(\rf_reg[67] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[360]$_DFFE_PN0P_  (.D(_0289_),
    .Q(\rf_reg[392] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[361]$_DFFE_PN0P_  (.D(_0290_),
    .Q(\rf_reg[393] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[362]$_DFFE_PN0P_  (.D(_0291_),
    .Q(\rf_reg[394] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[363]$_DFFE_PN0P_  (.D(_0292_),
    .Q(\rf_reg[395] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[364]$_DFFE_PN0P_  (.D(_0293_),
    .Q(\rf_reg[396] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[365]$_DFFE_PN0P_  (.D(_0294_),
    .Q(\rf_reg[397] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[366]$_DFFE_PN0P_  (.D(_0295_),
    .Q(\rf_reg[398] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[367]$_DFFE_PN0P_  (.D(_0296_),
    .Q(\rf_reg[399] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[368]$_DFFE_PN0P_  (.D(_0297_),
    .Q(\rf_reg[400] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[369]$_DFFE_PN0P_  (.D(_0298_),
    .Q(\rf_reg[401] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[36]$_DFFE_PN0P_  (.D(_0299_),
    .Q(\rf_reg[68] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[370]$_DFFE_PN0P_  (.D(_0300_),
    .Q(\rf_reg[402] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[371]$_DFFE_PN0P_  (.D(_0301_),
    .Q(\rf_reg[403] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[372]$_DFFE_PN0P_  (.D(_0302_),
    .Q(\rf_reg[404] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[373]$_DFFE_PN0P_  (.D(_0303_),
    .Q(\rf_reg[405] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[374]$_DFFE_PN0P_  (.D(_0304_),
    .Q(\rf_reg[406] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[375]$_DFFE_PN0P_  (.D(_0305_),
    .Q(\rf_reg[407] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[376]$_DFFE_PN0P_  (.D(_0306_),
    .Q(\rf_reg[408] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[377]$_DFFE_PN0P_  (.D(_0307_),
    .Q(\rf_reg[409] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[378]$_DFFE_PN0P_  (.D(_0308_),
    .Q(\rf_reg[410] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[379]$_DFFE_PN0P_  (.D(_0309_),
    .Q(\rf_reg[411] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[37]$_DFFE_PN0P_  (.D(_0310_),
    .Q(\rf_reg[69] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[380]$_DFFE_PN0P_  (.D(_0311_),
    .Q(\rf_reg[412] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[381]$_DFFE_PN0P_  (.D(_0312_),
    .Q(\rf_reg[413] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[382]$_DFFE_PN0P_  (.D(_0313_),
    .Q(\rf_reg[414] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[383]$_DFFE_PN0P_  (.D(_0314_),
    .Q(\rf_reg[415] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[384]$_DFFE_PN0P_  (.D(_0315_),
    .Q(\rf_reg[416] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[385]$_DFFE_PN0P_  (.D(_0316_),
    .Q(\rf_reg[417] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[386]$_DFFE_PN0P_  (.D(_0317_),
    .Q(\rf_reg[418] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[387]$_DFFE_PN0P_  (.D(_0318_),
    .Q(\rf_reg[419] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[388]$_DFFE_PN0P_  (.D(_0319_),
    .Q(\rf_reg[420] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[389]$_DFFE_PN0P_  (.D(_0320_),
    .Q(\rf_reg[421] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[38]$_DFFE_PN0P_  (.D(_0321_),
    .Q(\rf_reg[70] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[390]$_DFFE_PN0P_  (.D(_0322_),
    .Q(\rf_reg[422] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[391]$_DFFE_PN0P_  (.D(_0323_),
    .Q(\rf_reg[423] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[392]$_DFFE_PN0P_  (.D(_0324_),
    .Q(\rf_reg[424] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[393]$_DFFE_PN0P_  (.D(_0325_),
    .Q(\rf_reg[425] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[394]$_DFFE_PN0P_  (.D(_0326_),
    .Q(\rf_reg[426] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[395]$_DFFE_PN0P_  (.D(_0327_),
    .Q(\rf_reg[427] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[396]$_DFFE_PN0P_  (.D(_0328_),
    .Q(\rf_reg[428] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[397]$_DFFE_PN0P_  (.D(_0329_),
    .Q(\rf_reg[429] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[398]$_DFFE_PN0P_  (.D(_0330_),
    .Q(\rf_reg[430] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[399]$_DFFE_PN0P_  (.D(_0331_),
    .Q(\rf_reg[431] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[39]$_DFFE_PN0P_  (.D(_0332_),
    .Q(\rf_reg[71] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[3]$_DFFE_PN0P_  (.D(_0333_),
    .Q(\rf_reg[35] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[400]$_DFFE_PN0P_  (.D(_0334_),
    .Q(\rf_reg[432] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[401]$_DFFE_PN0P_  (.D(_0335_),
    .Q(\rf_reg[433] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[402]$_DFFE_PN0P_  (.D(_0336_),
    .Q(\rf_reg[434] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[403]$_DFFE_PN0P_  (.D(_0337_),
    .Q(\rf_reg[435] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[404]$_DFFE_PN0P_  (.D(_0338_),
    .Q(\rf_reg[436] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[405]$_DFFE_PN0P_  (.D(_0339_),
    .Q(\rf_reg[437] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[406]$_DFFE_PN0P_  (.D(_0340_),
    .Q(\rf_reg[438] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[407]$_DFFE_PN0P_  (.D(_0341_),
    .Q(\rf_reg[439] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[408]$_DFFE_PN0P_  (.D(_0342_),
    .Q(\rf_reg[440] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[409]$_DFFE_PN0P_  (.D(_0343_),
    .Q(\rf_reg[441] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[40]$_DFFE_PN0P_  (.D(_0344_),
    .Q(\rf_reg[72] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[410]$_DFFE_PN0P_  (.D(_0345_),
    .Q(\rf_reg[442] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[411]$_DFFE_PN0P_  (.D(_0346_),
    .Q(\rf_reg[443] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[412]$_DFFE_PN0P_  (.D(_0347_),
    .Q(\rf_reg[444] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[413]$_DFFE_PN0P_  (.D(_0348_),
    .Q(\rf_reg[445] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[414]$_DFFE_PN0P_  (.D(_0349_),
    .Q(\rf_reg[446] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[415]$_DFFE_PN0P_  (.D(_0350_),
    .Q(\rf_reg[447] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[416]$_DFFE_PN0P_  (.D(_0351_),
    .Q(\rf_reg[448] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[417]$_DFFE_PN0P_  (.D(_0352_),
    .Q(\rf_reg[449] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[418]$_DFFE_PN0P_  (.D(_0353_),
    .Q(\rf_reg[450] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[419]$_DFFE_PN0P_  (.D(_0354_),
    .Q(\rf_reg[451] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[41]$_DFFE_PN0P_  (.D(_0355_),
    .Q(\rf_reg[73] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[420]$_DFFE_PN0P_  (.D(_0356_),
    .Q(\rf_reg[452] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[421]$_DFFE_PN0P_  (.D(_0357_),
    .Q(\rf_reg[453] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[422]$_DFFE_PN0P_  (.D(_0358_),
    .Q(\rf_reg[454] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[423]$_DFFE_PN0P_  (.D(_0359_),
    .Q(\rf_reg[455] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[424]$_DFFE_PN0P_  (.D(_0360_),
    .Q(\rf_reg[456] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[425]$_DFFE_PN0P_  (.D(_0361_),
    .Q(\rf_reg[457] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[426]$_DFFE_PN0P_  (.D(_0362_),
    .Q(\rf_reg[458] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[427]$_DFFE_PN0P_  (.D(_0363_),
    .Q(\rf_reg[459] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[428]$_DFFE_PN0P_  (.D(_0364_),
    .Q(\rf_reg[460] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[429]$_DFFE_PN0P_  (.D(_0365_),
    .Q(\rf_reg[461] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[42]$_DFFE_PN0P_  (.D(_0366_),
    .Q(\rf_reg[74] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[430]$_DFFE_PN0P_  (.D(_0367_),
    .Q(\rf_reg[462] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[431]$_DFFE_PN0P_  (.D(_0368_),
    .Q(\rf_reg[463] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[432]$_DFFE_PN0P_  (.D(_0369_),
    .Q(\rf_reg[464] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[433]$_DFFE_PN0P_  (.D(_0370_),
    .Q(\rf_reg[465] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[434]$_DFFE_PN0P_  (.D(_0371_),
    .Q(\rf_reg[466] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[435]$_DFFE_PN0P_  (.D(_0372_),
    .Q(\rf_reg[467] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[436]$_DFFE_PN0P_  (.D(_0373_),
    .Q(\rf_reg[468] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[437]$_DFFE_PN0P_  (.D(_0374_),
    .Q(\rf_reg[469] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[438]$_DFFE_PN0P_  (.D(_0375_),
    .Q(\rf_reg[470] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[439]$_DFFE_PN0P_  (.D(_0376_),
    .Q(\rf_reg[471] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[43]$_DFFE_PN0P_  (.D(_0377_),
    .Q(\rf_reg[75] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[440]$_DFFE_PN0P_  (.D(_0378_),
    .Q(\rf_reg[472] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[441]$_DFFE_PN0P_  (.D(_0379_),
    .Q(\rf_reg[473] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[442]$_DFFE_PN0P_  (.D(_0380_),
    .Q(\rf_reg[474] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[443]$_DFFE_PN0P_  (.D(_0381_),
    .Q(\rf_reg[475] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[444]$_DFFE_PN0P_  (.D(_0382_),
    .Q(\rf_reg[476] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[445]$_DFFE_PN0P_  (.D(_0383_),
    .Q(\rf_reg[477] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[446]$_DFFE_PN0P_  (.D(_0384_),
    .Q(\rf_reg[478] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[447]$_DFFE_PN0P_  (.D(_0385_),
    .Q(\rf_reg[479] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[448]$_DFFE_PN0P_  (.D(_0386_),
    .Q(\rf_reg[480] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[449]$_DFFE_PN0P_  (.D(_0387_),
    .Q(\rf_reg[481] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[44]$_DFFE_PN0P_  (.D(_0388_),
    .Q(\rf_reg[76] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[450]$_DFFE_PN0P_  (.D(_0389_),
    .Q(\rf_reg[482] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[451]$_DFFE_PN0P_  (.D(_0390_),
    .Q(\rf_reg[483] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[452]$_DFFE_PN0P_  (.D(_0391_),
    .Q(\rf_reg[484] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[453]$_DFFE_PN0P_  (.D(_0392_),
    .Q(\rf_reg[485] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[454]$_DFFE_PN0P_  (.D(_0393_),
    .Q(\rf_reg[486] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[455]$_DFFE_PN0P_  (.D(_0394_),
    .Q(\rf_reg[487] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[456]$_DFFE_PN0P_  (.D(_0395_),
    .Q(\rf_reg[488] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[457]$_DFFE_PN0P_  (.D(_0396_),
    .Q(\rf_reg[489] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[458]$_DFFE_PN0P_  (.D(_0397_),
    .Q(\rf_reg[490] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[459]$_DFFE_PN0P_  (.D(_0398_),
    .Q(\rf_reg[491] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[45]$_DFFE_PN0P_  (.D(_0399_),
    .Q(\rf_reg[77] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[460]$_DFFE_PN0P_  (.D(_0400_),
    .Q(\rf_reg[492] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[461]$_DFFE_PN0P_  (.D(_0401_),
    .Q(\rf_reg[493] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[462]$_DFFE_PN0P_  (.D(_0402_),
    .Q(\rf_reg[494] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[463]$_DFFE_PN0P_  (.D(_0403_),
    .Q(\rf_reg[495] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[464]$_DFFE_PN0P_  (.D(_0404_),
    .Q(\rf_reg[496] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[465]$_DFFE_PN0P_  (.D(_0405_),
    .Q(\rf_reg[497] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[466]$_DFFE_PN0P_  (.D(_0406_),
    .Q(\rf_reg[498] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[467]$_DFFE_PN0P_  (.D(_0407_),
    .Q(\rf_reg[499] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[468]$_DFFE_PN0P_  (.D(_0408_),
    .Q(\rf_reg[500] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[469]$_DFFE_PN0P_  (.D(_0409_),
    .Q(\rf_reg[501] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[46]$_DFFE_PN0P_  (.D(_0410_),
    .Q(\rf_reg[78] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[470]$_DFFE_PN0P_  (.D(_0411_),
    .Q(\rf_reg[502] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[471]$_DFFE_PN0P_  (.D(_0412_),
    .Q(\rf_reg[503] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[472]$_DFFE_PN0P_  (.D(_0413_),
    .Q(\rf_reg[504] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[473]$_DFFE_PN0P_  (.D(_0414_),
    .Q(\rf_reg[505] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[474]$_DFFE_PN0P_  (.D(_0415_),
    .Q(\rf_reg[506] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[475]$_DFFE_PN0P_  (.D(_0416_),
    .Q(\rf_reg[507] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[476]$_DFFE_PN0P_  (.D(_0417_),
    .Q(\rf_reg[508] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[477]$_DFFE_PN0P_  (.D(_0418_),
    .Q(\rf_reg[509] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[478]$_DFFE_PN0P_  (.D(_0419_),
    .Q(\rf_reg[510] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[479]$_DFFE_PN0P_  (.D(_0420_),
    .Q(\rf_reg[511] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[47]$_DFFE_PN0P_  (.D(_0421_),
    .Q(\rf_reg[79] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[480]$_DFFE_PN0P_  (.D(_0422_),
    .Q(\rf_reg[512] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[481]$_DFFE_PN0P_  (.D(_0423_),
    .Q(\rf_reg[513] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[482]$_DFFE_PN0P_  (.D(_0424_),
    .Q(\rf_reg[514] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[483]$_DFFE_PN0P_  (.D(_0425_),
    .Q(\rf_reg[515] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[484]$_DFFE_PN0P_  (.D(_0426_),
    .Q(\rf_reg[516] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[485]$_DFFE_PN0P_  (.D(_0427_),
    .Q(\rf_reg[517] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[486]$_DFFE_PN0P_  (.D(_0428_),
    .Q(\rf_reg[518] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[487]$_DFFE_PN0P_  (.D(_0429_),
    .Q(\rf_reg[519] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[488]$_DFFE_PN0P_  (.D(_0430_),
    .Q(\rf_reg[520] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[489]$_DFFE_PN0P_  (.D(_0431_),
    .Q(\rf_reg[521] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[48]$_DFFE_PN0P_  (.D(_0432_),
    .Q(\rf_reg[80] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[490]$_DFFE_PN0P_  (.D(_0433_),
    .Q(\rf_reg[522] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[491]$_DFFE_PN0P_  (.D(_0434_),
    .Q(\rf_reg[523] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[492]$_DFFE_PN0P_  (.D(_0435_),
    .Q(\rf_reg[524] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[493]$_DFFE_PN0P_  (.D(_0436_),
    .Q(\rf_reg[525] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[494]$_DFFE_PN0P_  (.D(_0437_),
    .Q(\rf_reg[526] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[495]$_DFFE_PN0P_  (.D(_0438_),
    .Q(\rf_reg[527] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[496]$_DFFE_PN0P_  (.D(_0439_),
    .Q(\rf_reg[528] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[497]$_DFFE_PN0P_  (.D(_0440_),
    .Q(\rf_reg[529] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[498]$_DFFE_PN0P_  (.D(_0441_),
    .Q(\rf_reg[530] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[499]$_DFFE_PN0P_  (.D(_0442_),
    .Q(\rf_reg[531] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[49]$_DFFE_PN0P_  (.D(_0443_),
    .Q(\rf_reg[81] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[4]$_DFFE_PN0P_  (.D(_0444_),
    .Q(\rf_reg[36] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[500]$_DFFE_PN0P_  (.D(_0445_),
    .Q(\rf_reg[532] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[501]$_DFFE_PN0P_  (.D(_0446_),
    .Q(\rf_reg[533] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[502]$_DFFE_PN0P_  (.D(_0447_),
    .Q(\rf_reg[534] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[503]$_DFFE_PN0P_  (.D(_0448_),
    .Q(\rf_reg[535] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[504]$_DFFE_PN0P_  (.D(_0449_),
    .Q(\rf_reg[536] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[505]$_DFFE_PN0P_  (.D(_0450_),
    .Q(\rf_reg[537] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[506]$_DFFE_PN0P_  (.D(_0451_),
    .Q(\rf_reg[538] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[507]$_DFFE_PN0P_  (.D(_0452_),
    .Q(\rf_reg[539] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[508]$_DFFE_PN0P_  (.D(_0453_),
    .Q(\rf_reg[540] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[509]$_DFFE_PN0P_  (.D(_0454_),
    .Q(\rf_reg[541] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[50]$_DFFE_PN0P_  (.D(_0455_),
    .Q(\rf_reg[82] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[510]$_DFFE_PN0P_  (.D(_0456_),
    .Q(\rf_reg[542] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[511]$_DFFE_PN0P_  (.D(_0457_),
    .Q(\rf_reg[543] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[512]$_DFFE_PN0P_  (.D(_0458_),
    .Q(\rf_reg[544] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[513]$_DFFE_PN0P_  (.D(_0459_),
    .Q(\rf_reg[545] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[514]$_DFFE_PN0P_  (.D(_0460_),
    .Q(\rf_reg[546] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[515]$_DFFE_PN0P_  (.D(_0461_),
    .Q(\rf_reg[547] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[516]$_DFFE_PN0P_  (.D(_0462_),
    .Q(\rf_reg[548] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[517]$_DFFE_PN0P_  (.D(_0463_),
    .Q(\rf_reg[549] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[518]$_DFFE_PN0P_  (.D(_0464_),
    .Q(\rf_reg[550] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[519]$_DFFE_PN0P_  (.D(_0465_),
    .Q(\rf_reg[551] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[51]$_DFFE_PN0P_  (.D(_0466_),
    .Q(\rf_reg[83] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[520]$_DFFE_PN0P_  (.D(_0467_),
    .Q(\rf_reg[552] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[521]$_DFFE_PN0P_  (.D(_0468_),
    .Q(\rf_reg[553] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[522]$_DFFE_PN0P_  (.D(_0469_),
    .Q(\rf_reg[554] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[523]$_DFFE_PN0P_  (.D(_0470_),
    .Q(\rf_reg[555] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[524]$_DFFE_PN0P_  (.D(_0471_),
    .Q(\rf_reg[556] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[525]$_DFFE_PN0P_  (.D(_0472_),
    .Q(\rf_reg[557] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[526]$_DFFE_PN0P_  (.D(_0473_),
    .Q(\rf_reg[558] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[527]$_DFFE_PN0P_  (.D(_0474_),
    .Q(\rf_reg[559] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[528]$_DFFE_PN0P_  (.D(_0475_),
    .Q(\rf_reg[560] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[529]$_DFFE_PN0P_  (.D(_0476_),
    .Q(\rf_reg[561] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[52]$_DFFE_PN0P_  (.D(_0477_),
    .Q(\rf_reg[84] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[530]$_DFFE_PN0P_  (.D(_0478_),
    .Q(\rf_reg[562] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[531]$_DFFE_PN0P_  (.D(_0479_),
    .Q(\rf_reg[563] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[532]$_DFFE_PN0P_  (.D(_0480_),
    .Q(\rf_reg[564] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[533]$_DFFE_PN0P_  (.D(_0481_),
    .Q(\rf_reg[565] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[534]$_DFFE_PN0P_  (.D(_0482_),
    .Q(\rf_reg[566] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[535]$_DFFE_PN0P_  (.D(_0483_),
    .Q(\rf_reg[567] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[536]$_DFFE_PN0P_  (.D(_0484_),
    .Q(\rf_reg[568] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[537]$_DFFE_PN0P_  (.D(_0485_),
    .Q(\rf_reg[569] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[538]$_DFFE_PN0P_  (.D(_0486_),
    .Q(\rf_reg[570] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[539]$_DFFE_PN0P_  (.D(_0487_),
    .Q(\rf_reg[571] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[53]$_DFFE_PN0P_  (.D(_0488_),
    .Q(\rf_reg[85] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[540]$_DFFE_PN0P_  (.D(_0489_),
    .Q(\rf_reg[572] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[541]$_DFFE_PN0P_  (.D(_0490_),
    .Q(\rf_reg[573] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[542]$_DFFE_PN0P_  (.D(_0491_),
    .Q(\rf_reg[574] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[543]$_DFFE_PN0P_  (.D(_0492_),
    .Q(\rf_reg[575] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[544]$_DFFE_PN0P_  (.D(_0493_),
    .Q(\rf_reg[576] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[545]$_DFFE_PN0P_  (.D(_0494_),
    .Q(\rf_reg[577] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[546]$_DFFE_PN0P_  (.D(_0495_),
    .Q(\rf_reg[578] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[547]$_DFFE_PN0P_  (.D(_0496_),
    .Q(\rf_reg[579] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[548]$_DFFE_PN0P_  (.D(_0497_),
    .Q(\rf_reg[580] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[549]$_DFFE_PN0P_  (.D(_0498_),
    .Q(\rf_reg[581] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[54]$_DFFE_PN0P_  (.D(_0499_),
    .Q(\rf_reg[86] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[550]$_DFFE_PN0P_  (.D(_0500_),
    .Q(\rf_reg[582] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[551]$_DFFE_PN0P_  (.D(_0501_),
    .Q(\rf_reg[583] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[552]$_DFFE_PN0P_  (.D(_0502_),
    .Q(\rf_reg[584] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[553]$_DFFE_PN0P_  (.D(_0503_),
    .Q(\rf_reg[585] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[554]$_DFFE_PN0P_  (.D(_0504_),
    .Q(\rf_reg[586] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[555]$_DFFE_PN0P_  (.D(_0505_),
    .Q(\rf_reg[587] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[556]$_DFFE_PN0P_  (.D(_0506_),
    .Q(\rf_reg[588] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[557]$_DFFE_PN0P_  (.D(_0507_),
    .Q(\rf_reg[589] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[558]$_DFFE_PN0P_  (.D(_0508_),
    .Q(\rf_reg[590] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[559]$_DFFE_PN0P_  (.D(_0509_),
    .Q(\rf_reg[591] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[55]$_DFFE_PN0P_  (.D(_0510_),
    .Q(\rf_reg[87] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[560]$_DFFE_PN0P_  (.D(_0511_),
    .Q(\rf_reg[592] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[561]$_DFFE_PN0P_  (.D(_0512_),
    .Q(\rf_reg[593] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[562]$_DFFE_PN0P_  (.D(_0513_),
    .Q(\rf_reg[594] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[563]$_DFFE_PN0P_  (.D(_0514_),
    .Q(\rf_reg[595] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[564]$_DFFE_PN0P_  (.D(_0515_),
    .Q(\rf_reg[596] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[565]$_DFFE_PN0P_  (.D(_0516_),
    .Q(\rf_reg[597] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[566]$_DFFE_PN0P_  (.D(_0517_),
    .Q(\rf_reg[598] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[567]$_DFFE_PN0P_  (.D(_0518_),
    .Q(\rf_reg[599] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[568]$_DFFE_PN0P_  (.D(_0519_),
    .Q(\rf_reg[600] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[569]$_DFFE_PN0P_  (.D(_0520_),
    .Q(\rf_reg[601] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[56]$_DFFE_PN0P_  (.D(_0521_),
    .Q(\rf_reg[88] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[570]$_DFFE_PN0P_  (.D(_0522_),
    .Q(\rf_reg[602] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[571]$_DFFE_PN0P_  (.D(_0523_),
    .Q(\rf_reg[603] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[572]$_DFFE_PN0P_  (.D(_0524_),
    .Q(\rf_reg[604] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[573]$_DFFE_PN0P_  (.D(_0525_),
    .Q(\rf_reg[605] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[574]$_DFFE_PN0P_  (.D(_0526_),
    .Q(\rf_reg[606] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[575]$_DFFE_PN0P_  (.D(_0527_),
    .Q(\rf_reg[607] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[576]$_DFFE_PN0P_  (.D(_0528_),
    .Q(\rf_reg[608] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[577]$_DFFE_PN0P_  (.D(_0529_),
    .Q(\rf_reg[609] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[578]$_DFFE_PN0P_  (.D(_0530_),
    .Q(\rf_reg[610] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[579]$_DFFE_PN0P_  (.D(_0531_),
    .Q(\rf_reg[611] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[57]$_DFFE_PN0P_  (.D(_0532_),
    .Q(\rf_reg[89] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[580]$_DFFE_PN0P_  (.D(_0533_),
    .Q(\rf_reg[612] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[581]$_DFFE_PN0P_  (.D(_0534_),
    .Q(\rf_reg[613] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[582]$_DFFE_PN0P_  (.D(_0535_),
    .Q(\rf_reg[614] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[583]$_DFFE_PN0P_  (.D(_0536_),
    .Q(\rf_reg[615] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[584]$_DFFE_PN0P_  (.D(_0537_),
    .Q(\rf_reg[616] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[585]$_DFFE_PN0P_  (.D(_0538_),
    .Q(\rf_reg[617] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[586]$_DFFE_PN0P_  (.D(_0539_),
    .Q(\rf_reg[618] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[587]$_DFFE_PN0P_  (.D(_0540_),
    .Q(\rf_reg[619] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[588]$_DFFE_PN0P_  (.D(_0541_),
    .Q(\rf_reg[620] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[589]$_DFFE_PN0P_  (.D(_0542_),
    .Q(\rf_reg[621] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[58]$_DFFE_PN0P_  (.D(_0543_),
    .Q(\rf_reg[90] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[590]$_DFFE_PN0P_  (.D(_0544_),
    .Q(\rf_reg[622] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[591]$_DFFE_PN0P_  (.D(_0545_),
    .Q(\rf_reg[623] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[592]$_DFFE_PN0P_  (.D(_0546_),
    .Q(\rf_reg[624] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[593]$_DFFE_PN0P_  (.D(_0547_),
    .Q(\rf_reg[625] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[594]$_DFFE_PN0P_  (.D(_0548_),
    .Q(\rf_reg[626] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[595]$_DFFE_PN0P_  (.D(_0549_),
    .Q(\rf_reg[627] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[596]$_DFFE_PN0P_  (.D(_0550_),
    .Q(\rf_reg[628] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[597]$_DFFE_PN0P_  (.D(_0551_),
    .Q(\rf_reg[629] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[598]$_DFFE_PN0P_  (.D(_0552_),
    .Q(\rf_reg[630] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[599]$_DFFE_PN0P_  (.D(_0553_),
    .Q(\rf_reg[631] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[59]$_DFFE_PN0P_  (.D(_0554_),
    .Q(\rf_reg[91] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[5]$_DFFE_PN0P_  (.D(_0555_),
    .Q(\rf_reg[37] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[600]$_DFFE_PN0P_  (.D(_0556_),
    .Q(\rf_reg[632] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[601]$_DFFE_PN0P_  (.D(_0557_),
    .Q(\rf_reg[633] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[602]$_DFFE_PN0P_  (.D(_0558_),
    .Q(\rf_reg[634] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[603]$_DFFE_PN0P_  (.D(_0559_),
    .Q(\rf_reg[635] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[604]$_DFFE_PN0P_  (.D(_0560_),
    .Q(\rf_reg[636] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[605]$_DFFE_PN0P_  (.D(_0561_),
    .Q(\rf_reg[637] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[606]$_DFFE_PN0P_  (.D(_0562_),
    .Q(\rf_reg[638] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[607]$_DFFE_PN0P_  (.D(_0563_),
    .Q(\rf_reg[639] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[608]$_DFFE_PN0P_  (.D(_0564_),
    .Q(\rf_reg[640] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[609]$_DFFE_PN0P_  (.D(_0565_),
    .Q(\rf_reg[641] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[60]$_DFFE_PN0P_  (.D(_0566_),
    .Q(\rf_reg[92] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[610]$_DFFE_PN0P_  (.D(_0567_),
    .Q(\rf_reg[642] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[611]$_DFFE_PN0P_  (.D(_0568_),
    .Q(\rf_reg[643] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[612]$_DFFE_PN0P_  (.D(_0569_),
    .Q(\rf_reg[644] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[613]$_DFFE_PN0P_  (.D(_0570_),
    .Q(\rf_reg[645] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[614]$_DFFE_PN0P_  (.D(_0571_),
    .Q(\rf_reg[646] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[615]$_DFFE_PN0P_  (.D(_0572_),
    .Q(\rf_reg[647] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[616]$_DFFE_PN0P_  (.D(_0573_),
    .Q(\rf_reg[648] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[617]$_DFFE_PN0P_  (.D(_0574_),
    .Q(\rf_reg[649] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[618]$_DFFE_PN0P_  (.D(_0575_),
    .Q(\rf_reg[650] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[619]$_DFFE_PN0P_  (.D(_0576_),
    .Q(\rf_reg[651] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[61]$_DFFE_PN0P_  (.D(_0577_),
    .Q(\rf_reg[93] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[620]$_DFFE_PN0P_  (.D(_0578_),
    .Q(\rf_reg[652] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[621]$_DFFE_PN0P_  (.D(_0579_),
    .Q(\rf_reg[653] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[622]$_DFFE_PN0P_  (.D(_0580_),
    .Q(\rf_reg[654] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[623]$_DFFE_PN0P_  (.D(_0581_),
    .Q(\rf_reg[655] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[624]$_DFFE_PN0P_  (.D(_0582_),
    .Q(\rf_reg[656] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[625]$_DFFE_PN0P_  (.D(_0583_),
    .Q(\rf_reg[657] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[626]$_DFFE_PN0P_  (.D(_0584_),
    .Q(\rf_reg[658] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[627]$_DFFE_PN0P_  (.D(_0585_),
    .Q(\rf_reg[659] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[628]$_DFFE_PN0P_  (.D(_0586_),
    .Q(\rf_reg[660] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[629]$_DFFE_PN0P_  (.D(_0587_),
    .Q(\rf_reg[661] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[62]$_DFFE_PN0P_  (.D(_0588_),
    .Q(\rf_reg[94] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[630]$_DFFE_PN0P_  (.D(_0589_),
    .Q(\rf_reg[662] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[631]$_DFFE_PN0P_  (.D(_0590_),
    .Q(\rf_reg[663] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[632]$_DFFE_PN0P_  (.D(_0591_),
    .Q(\rf_reg[664] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[633]$_DFFE_PN0P_  (.D(_0592_),
    .Q(\rf_reg[665] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[634]$_DFFE_PN0P_  (.D(_0593_),
    .Q(\rf_reg[666] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[635]$_DFFE_PN0P_  (.D(_0594_),
    .Q(\rf_reg[667] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[636]$_DFFE_PN0P_  (.D(_0595_),
    .Q(\rf_reg[668] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[637]$_DFFE_PN0P_  (.D(_0596_),
    .Q(\rf_reg[669] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[638]$_DFFE_PN0P_  (.D(_0597_),
    .Q(\rf_reg[670] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[639]$_DFFE_PN0P_  (.D(_0598_),
    .Q(\rf_reg[671] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[63]$_DFFE_PN0P_  (.D(_0599_),
    .Q(\rf_reg[95] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[640]$_DFFE_PN0P_  (.D(_0600_),
    .Q(\rf_reg[672] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[641]$_DFFE_PN0P_  (.D(_0601_),
    .Q(\rf_reg[673] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[642]$_DFFE_PN0P_  (.D(_0602_),
    .Q(\rf_reg[674] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[643]$_DFFE_PN0P_  (.D(_0603_),
    .Q(\rf_reg[675] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[644]$_DFFE_PN0P_  (.D(_0604_),
    .Q(\rf_reg[676] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[645]$_DFFE_PN0P_  (.D(_0605_),
    .Q(\rf_reg[677] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[646]$_DFFE_PN0P_  (.D(_0606_),
    .Q(\rf_reg[678] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[647]$_DFFE_PN0P_  (.D(_0607_),
    .Q(\rf_reg[679] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[648]$_DFFE_PN0P_  (.D(_0608_),
    .Q(\rf_reg[680] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[649]$_DFFE_PN0P_  (.D(_0609_),
    .Q(\rf_reg[681] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[64]$_DFFE_PN0P_  (.D(_0610_),
    .Q(\rf_reg[96] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[650]$_DFFE_PN0P_  (.D(_0611_),
    .Q(\rf_reg[682] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[651]$_DFFE_PN0P_  (.D(_0612_),
    .Q(\rf_reg[683] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[652]$_DFFE_PN0P_  (.D(_0613_),
    .Q(\rf_reg[684] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[653]$_DFFE_PN0P_  (.D(_0614_),
    .Q(\rf_reg[685] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[654]$_DFFE_PN0P_  (.D(_0615_),
    .Q(\rf_reg[686] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[655]$_DFFE_PN0P_  (.D(_0616_),
    .Q(\rf_reg[687] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[656]$_DFFE_PN0P_  (.D(_0617_),
    .Q(\rf_reg[688] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[657]$_DFFE_PN0P_  (.D(_0618_),
    .Q(\rf_reg[689] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[658]$_DFFE_PN0P_  (.D(_0619_),
    .Q(\rf_reg[690] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[659]$_DFFE_PN0P_  (.D(_0620_),
    .Q(\rf_reg[691] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[65]$_DFFE_PN0P_  (.D(_0621_),
    .Q(\rf_reg[97] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[660]$_DFFE_PN0P_  (.D(_0622_),
    .Q(\rf_reg[692] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[661]$_DFFE_PN0P_  (.D(_0623_),
    .Q(\rf_reg[693] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[662]$_DFFE_PN0P_  (.D(_0624_),
    .Q(\rf_reg[694] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[663]$_DFFE_PN0P_  (.D(_0625_),
    .Q(\rf_reg[695] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[664]$_DFFE_PN0P_  (.D(_0626_),
    .Q(\rf_reg[696] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[665]$_DFFE_PN0P_  (.D(_0627_),
    .Q(\rf_reg[697] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[666]$_DFFE_PN0P_  (.D(_0628_),
    .Q(\rf_reg[698] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[667]$_DFFE_PN0P_  (.D(_0629_),
    .Q(\rf_reg[699] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[668]$_DFFE_PN0P_  (.D(_0630_),
    .Q(\rf_reg[700] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[669]$_DFFE_PN0P_  (.D(_0631_),
    .Q(\rf_reg[701] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[66]$_DFFE_PN0P_  (.D(_0632_),
    .Q(\rf_reg[98] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[670]$_DFFE_PN0P_  (.D(_0633_),
    .Q(\rf_reg[702] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[671]$_DFFE_PN0P_  (.D(_0634_),
    .Q(\rf_reg[703] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[672]$_DFFE_PN0P_  (.D(_0635_),
    .Q(\rf_reg[704] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[673]$_DFFE_PN0P_  (.D(_0636_),
    .Q(\rf_reg[705] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[674]$_DFFE_PN0P_  (.D(_0637_),
    .Q(\rf_reg[706] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[675]$_DFFE_PN0P_  (.D(_0638_),
    .Q(\rf_reg[707] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[676]$_DFFE_PN0P_  (.D(_0639_),
    .Q(\rf_reg[708] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[677]$_DFFE_PN0P_  (.D(_0640_),
    .Q(\rf_reg[709] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[678]$_DFFE_PN0P_  (.D(_0641_),
    .Q(\rf_reg[710] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[679]$_DFFE_PN0P_  (.D(_0642_),
    .Q(\rf_reg[711] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[67]$_DFFE_PN0P_  (.D(_0643_),
    .Q(\rf_reg[99] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[680]$_DFFE_PN0P_  (.D(_0644_),
    .Q(\rf_reg[712] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[681]$_DFFE_PN0P_  (.D(_0645_),
    .Q(\rf_reg[713] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[682]$_DFFE_PN0P_  (.D(_0646_),
    .Q(\rf_reg[714] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[683]$_DFFE_PN0P_  (.D(_0647_),
    .Q(\rf_reg[715] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[684]$_DFFE_PN0P_  (.D(_0648_),
    .Q(\rf_reg[716] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[685]$_DFFE_PN0P_  (.D(_0649_),
    .Q(\rf_reg[717] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[686]$_DFFE_PN0P_  (.D(_0650_),
    .Q(\rf_reg[718] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[687]$_DFFE_PN0P_  (.D(_0651_),
    .Q(\rf_reg[719] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[688]$_DFFE_PN0P_  (.D(_0652_),
    .Q(\rf_reg[720] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[689]$_DFFE_PN0P_  (.D(_0653_),
    .Q(\rf_reg[721] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[68]$_DFFE_PN0P_  (.D(_0654_),
    .Q(\rf_reg[100] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[690]$_DFFE_PN0P_  (.D(_0655_),
    .Q(\rf_reg[722] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[691]$_DFFE_PN0P_  (.D(_0656_),
    .Q(\rf_reg[723] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[692]$_DFFE_PN0P_  (.D(_0657_),
    .Q(\rf_reg[724] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[693]$_DFFE_PN0P_  (.D(_0658_),
    .Q(\rf_reg[725] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[694]$_DFFE_PN0P_  (.D(_0659_),
    .Q(\rf_reg[726] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[695]$_DFFE_PN0P_  (.D(_0660_),
    .Q(\rf_reg[727] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[696]$_DFFE_PN0P_  (.D(_0661_),
    .Q(\rf_reg[728] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[697]$_DFFE_PN0P_  (.D(_0662_),
    .Q(\rf_reg[729] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[698]$_DFFE_PN0P_  (.D(_0663_),
    .Q(\rf_reg[730] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[699]$_DFFE_PN0P_  (.D(_0664_),
    .Q(\rf_reg[731] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[69]$_DFFE_PN0P_  (.D(_0665_),
    .Q(\rf_reg[101] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[6]$_DFFE_PN0P_  (.D(_0666_),
    .Q(\rf_reg[38] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[700]$_DFFE_PN0P_  (.D(_0667_),
    .Q(\rf_reg[732] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[701]$_DFFE_PN0P_  (.D(_0668_),
    .Q(\rf_reg[733] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[702]$_DFFE_PN0P_  (.D(_0669_),
    .Q(\rf_reg[734] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[703]$_DFFE_PN0P_  (.D(_0670_),
    .Q(\rf_reg[735] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[704]$_DFFE_PN0P_  (.D(_0671_),
    .Q(\rf_reg[736] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[705]$_DFFE_PN0P_  (.D(_0672_),
    .Q(\rf_reg[737] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[706]$_DFFE_PN0P_  (.D(_0673_),
    .Q(\rf_reg[738] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[707]$_DFFE_PN0P_  (.D(_0674_),
    .Q(\rf_reg[739] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[708]$_DFFE_PN0P_  (.D(_0675_),
    .Q(\rf_reg[740] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[709]$_DFFE_PN0P_  (.D(_0676_),
    .Q(\rf_reg[741] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[70]$_DFFE_PN0P_  (.D(_0677_),
    .Q(\rf_reg[102] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[710]$_DFFE_PN0P_  (.D(_0678_),
    .Q(\rf_reg[742] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[711]$_DFFE_PN0P_  (.D(_0679_),
    .Q(\rf_reg[743] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[712]$_DFFE_PN0P_  (.D(_0680_),
    .Q(\rf_reg[744] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[713]$_DFFE_PN0P_  (.D(_0681_),
    .Q(\rf_reg[745] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[714]$_DFFE_PN0P_  (.D(_0682_),
    .Q(\rf_reg[746] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[715]$_DFFE_PN0P_  (.D(_0683_),
    .Q(\rf_reg[747] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[716]$_DFFE_PN0P_  (.D(_0684_),
    .Q(\rf_reg[748] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[717]$_DFFE_PN0P_  (.D(_0685_),
    .Q(\rf_reg[749] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[718]$_DFFE_PN0P_  (.D(_0686_),
    .Q(\rf_reg[750] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[719]$_DFFE_PN0P_  (.D(_0687_),
    .Q(\rf_reg[751] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[71]$_DFFE_PN0P_  (.D(_0688_),
    .Q(\rf_reg[103] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[720]$_DFFE_PN0P_  (.D(_0689_),
    .Q(\rf_reg[752] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[721]$_DFFE_PN0P_  (.D(_0690_),
    .Q(\rf_reg[753] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[722]$_DFFE_PN0P_  (.D(_0691_),
    .Q(\rf_reg[754] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[723]$_DFFE_PN0P_  (.D(_0692_),
    .Q(\rf_reg[755] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[724]$_DFFE_PN0P_  (.D(_0693_),
    .Q(\rf_reg[756] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[725]$_DFFE_PN0P_  (.D(_0694_),
    .Q(\rf_reg[757] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[726]$_DFFE_PN0P_  (.D(_0695_),
    .Q(\rf_reg[758] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[727]$_DFFE_PN0P_  (.D(_0696_),
    .Q(\rf_reg[759] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[728]$_DFFE_PN0P_  (.D(_0697_),
    .Q(\rf_reg[760] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[729]$_DFFE_PN0P_  (.D(_0698_),
    .Q(\rf_reg[761] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[72]$_DFFE_PN0P_  (.D(_0699_),
    .Q(\rf_reg[104] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[730]$_DFFE_PN0P_  (.D(_0700_),
    .Q(\rf_reg[762] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[731]$_DFFE_PN0P_  (.D(_0701_),
    .Q(\rf_reg[763] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[732]$_DFFE_PN0P_  (.D(_0702_),
    .Q(\rf_reg[764] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[733]$_DFFE_PN0P_  (.D(_0703_),
    .Q(\rf_reg[765] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[734]$_DFFE_PN0P_  (.D(_0704_),
    .Q(\rf_reg[766] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[735]$_DFFE_PN0P_  (.D(_0705_),
    .Q(\rf_reg[767] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[736]$_DFFE_PN0P_  (.D(_0706_),
    .Q(\rf_reg[768] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[737]$_DFFE_PN0P_  (.D(_0707_),
    .Q(\rf_reg[769] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[738]$_DFFE_PN0P_  (.D(_0708_),
    .Q(\rf_reg[770] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[739]$_DFFE_PN0P_  (.D(_0709_),
    .Q(\rf_reg[771] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[73]$_DFFE_PN0P_  (.D(_0710_),
    .Q(\rf_reg[105] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[740]$_DFFE_PN0P_  (.D(_0711_),
    .Q(\rf_reg[772] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[741]$_DFFE_PN0P_  (.D(_0712_),
    .Q(\rf_reg[773] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[742]$_DFFE_PN0P_  (.D(_0713_),
    .Q(\rf_reg[774] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[743]$_DFFE_PN0P_  (.D(_0714_),
    .Q(\rf_reg[775] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[744]$_DFFE_PN0P_  (.D(_0715_),
    .Q(\rf_reg[776] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[745]$_DFFE_PN0P_  (.D(_0716_),
    .Q(\rf_reg[777] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[746]$_DFFE_PN0P_  (.D(_0717_),
    .Q(\rf_reg[778] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[747]$_DFFE_PN0P_  (.D(_0718_),
    .Q(\rf_reg[779] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[748]$_DFFE_PN0P_  (.D(_0719_),
    .Q(\rf_reg[780] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[749]$_DFFE_PN0P_  (.D(_0720_),
    .Q(\rf_reg[781] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[74]$_DFFE_PN0P_  (.D(_0721_),
    .Q(\rf_reg[106] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[750]$_DFFE_PN0P_  (.D(_0722_),
    .Q(\rf_reg[782] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[751]$_DFFE_PN0P_  (.D(_0723_),
    .Q(\rf_reg[783] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[752]$_DFFE_PN0P_  (.D(_0724_),
    .Q(\rf_reg[784] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[753]$_DFFE_PN0P_  (.D(_0725_),
    .Q(\rf_reg[785] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[754]$_DFFE_PN0P_  (.D(_0726_),
    .Q(\rf_reg[786] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[755]$_DFFE_PN0P_  (.D(_0727_),
    .Q(\rf_reg[787] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[756]$_DFFE_PN0P_  (.D(_0728_),
    .Q(\rf_reg[788] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[757]$_DFFE_PN0P_  (.D(_0729_),
    .Q(\rf_reg[789] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[758]$_DFFE_PN0P_  (.D(_0730_),
    .Q(\rf_reg[790] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[759]$_DFFE_PN0P_  (.D(_0731_),
    .Q(\rf_reg[791] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[75]$_DFFE_PN0P_  (.D(_0732_),
    .Q(\rf_reg[107] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[760]$_DFFE_PN0P_  (.D(_0733_),
    .Q(\rf_reg[792] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[761]$_DFFE_PN0P_  (.D(_0734_),
    .Q(\rf_reg[793] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[762]$_DFFE_PN0P_  (.D(_0735_),
    .Q(\rf_reg[794] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[763]$_DFFE_PN0P_  (.D(_0736_),
    .Q(\rf_reg[795] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[764]$_DFFE_PN0P_  (.D(_0737_),
    .Q(\rf_reg[796] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[765]$_DFFE_PN0P_  (.D(_0738_),
    .Q(\rf_reg[797] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[766]$_DFFE_PN0P_  (.D(_0739_),
    .Q(\rf_reg[798] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[767]$_DFFE_PN0P_  (.D(_0740_),
    .Q(\rf_reg[799] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[768]$_DFFE_PN0P_  (.D(_0741_),
    .Q(\rf_reg[800] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[769]$_DFFE_PN0P_  (.D(_0742_),
    .Q(\rf_reg[801] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[76]$_DFFE_PN0P_  (.D(_0743_),
    .Q(\rf_reg[108] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[770]$_DFFE_PN0P_  (.D(_0744_),
    .Q(\rf_reg[802] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[771]$_DFFE_PN0P_  (.D(_0745_),
    .Q(\rf_reg[803] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[772]$_DFFE_PN0P_  (.D(_0746_),
    .Q(\rf_reg[804] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[773]$_DFFE_PN0P_  (.D(_0747_),
    .Q(\rf_reg[805] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[774]$_DFFE_PN0P_  (.D(_0748_),
    .Q(\rf_reg[806] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[775]$_DFFE_PN0P_  (.D(_0749_),
    .Q(\rf_reg[807] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[776]$_DFFE_PN0P_  (.D(_0750_),
    .Q(\rf_reg[808] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[777]$_DFFE_PN0P_  (.D(_0751_),
    .Q(\rf_reg[809] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[778]$_DFFE_PN0P_  (.D(_0752_),
    .Q(\rf_reg[810] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[779]$_DFFE_PN0P_  (.D(_0753_),
    .Q(\rf_reg[811] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[77]$_DFFE_PN0P_  (.D(_0754_),
    .Q(\rf_reg[109] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[780]$_DFFE_PN0P_  (.D(_0755_),
    .Q(\rf_reg[812] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[781]$_DFFE_PN0P_  (.D(_0756_),
    .Q(\rf_reg[813] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[782]$_DFFE_PN0P_  (.D(_0757_),
    .Q(\rf_reg[814] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[783]$_DFFE_PN0P_  (.D(_0758_),
    .Q(\rf_reg[815] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[784]$_DFFE_PN0P_  (.D(_0759_),
    .Q(\rf_reg[816] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[785]$_DFFE_PN0P_  (.D(_0760_),
    .Q(\rf_reg[817] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[786]$_DFFE_PN0P_  (.D(_0761_),
    .Q(\rf_reg[818] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[787]$_DFFE_PN0P_  (.D(_0762_),
    .Q(\rf_reg[819] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[788]$_DFFE_PN0P_  (.D(_0763_),
    .Q(\rf_reg[820] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[789]$_DFFE_PN0P_  (.D(_0764_),
    .Q(\rf_reg[821] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[78]$_DFFE_PN0P_  (.D(_0765_),
    .Q(\rf_reg[110] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[790]$_DFFE_PN0P_  (.D(_0766_),
    .Q(\rf_reg[822] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[791]$_DFFE_PN0P_  (.D(_0767_),
    .Q(\rf_reg[823] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[792]$_DFFE_PN0P_  (.D(_0768_),
    .Q(\rf_reg[824] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[793]$_DFFE_PN0P_  (.D(_0769_),
    .Q(\rf_reg[825] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[794]$_DFFE_PN0P_  (.D(_0770_),
    .Q(\rf_reg[826] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[795]$_DFFE_PN0P_  (.D(_0771_),
    .Q(\rf_reg[827] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[796]$_DFFE_PN0P_  (.D(_0772_),
    .Q(\rf_reg[828] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[797]$_DFFE_PN0P_  (.D(_0773_),
    .Q(\rf_reg[829] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[798]$_DFFE_PN0P_  (.D(_0774_),
    .Q(\rf_reg[830] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[799]$_DFFE_PN0P_  (.D(_0775_),
    .Q(\rf_reg[831] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[79]$_DFFE_PN0P_  (.D(_0776_),
    .Q(\rf_reg[111] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[7]$_DFFE_PN0P_  (.D(_0777_),
    .Q(\rf_reg[39] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[800]$_DFFE_PN0P_  (.D(_0778_),
    .Q(\rf_reg[832] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[801]$_DFFE_PN0P_  (.D(_0779_),
    .Q(\rf_reg[833] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[802]$_DFFE_PN0P_  (.D(_0780_),
    .Q(\rf_reg[834] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[803]$_DFFE_PN0P_  (.D(_0781_),
    .Q(\rf_reg[835] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[804]$_DFFE_PN0P_  (.D(_0782_),
    .Q(\rf_reg[836] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[805]$_DFFE_PN0P_  (.D(_0783_),
    .Q(\rf_reg[837] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[806]$_DFFE_PN0P_  (.D(_0784_),
    .Q(\rf_reg[838] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[807]$_DFFE_PN0P_  (.D(_0785_),
    .Q(\rf_reg[839] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[808]$_DFFE_PN0P_  (.D(_0786_),
    .Q(\rf_reg[840] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[809]$_DFFE_PN0P_  (.D(_0787_),
    .Q(\rf_reg[841] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[80]$_DFFE_PN0P_  (.D(_0788_),
    .Q(\rf_reg[112] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[810]$_DFFE_PN0P_  (.D(_0789_),
    .Q(\rf_reg[842] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[811]$_DFFE_PN0P_  (.D(_0790_),
    .Q(\rf_reg[843] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[812]$_DFFE_PN0P_  (.D(_0791_),
    .Q(\rf_reg[844] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[813]$_DFFE_PN0P_  (.D(_0792_),
    .Q(\rf_reg[845] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[814]$_DFFE_PN0P_  (.D(_0793_),
    .Q(\rf_reg[846] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[815]$_DFFE_PN0P_  (.D(_0794_),
    .Q(\rf_reg[847] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[816]$_DFFE_PN0P_  (.D(_0795_),
    .Q(\rf_reg[848] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[817]$_DFFE_PN0P_  (.D(_0796_),
    .Q(\rf_reg[849] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[818]$_DFFE_PN0P_  (.D(_0797_),
    .Q(\rf_reg[850] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[819]$_DFFE_PN0P_  (.D(_0798_),
    .Q(\rf_reg[851] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[81]$_DFFE_PN0P_  (.D(_0799_),
    .Q(\rf_reg[113] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[820]$_DFFE_PN0P_  (.D(_0800_),
    .Q(\rf_reg[852] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[821]$_DFFE_PN0P_  (.D(_0801_),
    .Q(\rf_reg[853] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[822]$_DFFE_PN0P_  (.D(_0802_),
    .Q(\rf_reg[854] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[823]$_DFFE_PN0P_  (.D(_0803_),
    .Q(\rf_reg[855] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[824]$_DFFE_PN0P_  (.D(_0804_),
    .Q(\rf_reg[856] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[825]$_DFFE_PN0P_  (.D(_0805_),
    .Q(\rf_reg[857] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[826]$_DFFE_PN0P_  (.D(_0806_),
    .Q(\rf_reg[858] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[827]$_DFFE_PN0P_  (.D(_0807_),
    .Q(\rf_reg[859] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[828]$_DFFE_PN0P_  (.D(_0808_),
    .Q(\rf_reg[860] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[829]$_DFFE_PN0P_  (.D(_0809_),
    .Q(\rf_reg[861] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[82]$_DFFE_PN0P_  (.D(_0810_),
    .Q(\rf_reg[114] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[830]$_DFFE_PN0P_  (.D(_0811_),
    .Q(\rf_reg[862] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[831]$_DFFE_PN0P_  (.D(_0812_),
    .Q(\rf_reg[863] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[832]$_DFFE_PN0P_  (.D(_0813_),
    .Q(\rf_reg[864] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[833]$_DFFE_PN0P_  (.D(_0814_),
    .Q(\rf_reg[865] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[834]$_DFFE_PN0P_  (.D(_0815_),
    .Q(\rf_reg[866] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[835]$_DFFE_PN0P_  (.D(_0816_),
    .Q(\rf_reg[867] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[836]$_DFFE_PN0P_  (.D(_0817_),
    .Q(\rf_reg[868] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[837]$_DFFE_PN0P_  (.D(_0818_),
    .Q(\rf_reg[869] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[838]$_DFFE_PN0P_  (.D(_0819_),
    .Q(\rf_reg[870] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[839]$_DFFE_PN0P_  (.D(_0820_),
    .Q(\rf_reg[871] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[83]$_DFFE_PN0P_  (.D(_0821_),
    .Q(\rf_reg[115] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[840]$_DFFE_PN0P_  (.D(_0822_),
    .Q(\rf_reg[872] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[841]$_DFFE_PN0P_  (.D(_0823_),
    .Q(\rf_reg[873] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[842]$_DFFE_PN0P_  (.D(_0824_),
    .Q(\rf_reg[874] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[843]$_DFFE_PN0P_  (.D(_0825_),
    .Q(\rf_reg[875] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[844]$_DFFE_PN0P_  (.D(_0826_),
    .Q(\rf_reg[876] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[845]$_DFFE_PN0P_  (.D(_0827_),
    .Q(\rf_reg[877] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[846]$_DFFE_PN0P_  (.D(_0828_),
    .Q(\rf_reg[878] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[847]$_DFFE_PN0P_  (.D(_0829_),
    .Q(\rf_reg[879] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[848]$_DFFE_PN0P_  (.D(_0830_),
    .Q(\rf_reg[880] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[849]$_DFFE_PN0P_  (.D(_0831_),
    .Q(\rf_reg[881] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[84]$_DFFE_PN0P_  (.D(_0832_),
    .Q(\rf_reg[116] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[850]$_DFFE_PN0P_  (.D(_0833_),
    .Q(\rf_reg[882] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[851]$_DFFE_PN0P_  (.D(_0834_),
    .Q(\rf_reg[883] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[852]$_DFFE_PN0P_  (.D(_0835_),
    .Q(\rf_reg[884] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[853]$_DFFE_PN0P_  (.D(_0836_),
    .Q(\rf_reg[885] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[854]$_DFFE_PN0P_  (.D(_0837_),
    .Q(\rf_reg[886] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[855]$_DFFE_PN0P_  (.D(_0838_),
    .Q(\rf_reg[887] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[856]$_DFFE_PN0P_  (.D(_0839_),
    .Q(\rf_reg[888] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[857]$_DFFE_PN0P_  (.D(_0840_),
    .Q(\rf_reg[889] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[858]$_DFFE_PN0P_  (.D(_0841_),
    .Q(\rf_reg[890] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[859]$_DFFE_PN0P_  (.D(_0842_),
    .Q(\rf_reg[891] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[85]$_DFFE_PN0P_  (.D(_0843_),
    .Q(\rf_reg[117] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[860]$_DFFE_PN0P_  (.D(_0844_),
    .Q(\rf_reg[892] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[861]$_DFFE_PN0P_  (.D(_0845_),
    .Q(\rf_reg[893] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[862]$_DFFE_PN0P_  (.D(_0846_),
    .Q(\rf_reg[894] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[863]$_DFFE_PN0P_  (.D(_0847_),
    .Q(\rf_reg[895] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[864]$_DFFE_PN0P_  (.D(_0848_),
    .Q(\rf_reg[896] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[865]$_DFFE_PN0P_  (.D(_0849_),
    .Q(\rf_reg[897] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[866]$_DFFE_PN0P_  (.D(_0850_),
    .Q(\rf_reg[898] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[867]$_DFFE_PN0P_  (.D(_0851_),
    .Q(\rf_reg[899] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[868]$_DFFE_PN0P_  (.D(_0852_),
    .Q(\rf_reg[900] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[869]$_DFFE_PN0P_  (.D(_0853_),
    .Q(\rf_reg[901] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[86]$_DFFE_PN0P_  (.D(_0854_),
    .Q(\rf_reg[118] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[870]$_DFFE_PN0P_  (.D(_0855_),
    .Q(\rf_reg[902] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[871]$_DFFE_PN0P_  (.D(_0856_),
    .Q(\rf_reg[903] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[872]$_DFFE_PN0P_  (.D(_0857_),
    .Q(\rf_reg[904] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[873]$_DFFE_PN0P_  (.D(_0858_),
    .Q(\rf_reg[905] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[874]$_DFFE_PN0P_  (.D(_0859_),
    .Q(\rf_reg[906] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[875]$_DFFE_PN0P_  (.D(_0860_),
    .Q(\rf_reg[907] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[876]$_DFFE_PN0P_  (.D(_0861_),
    .Q(\rf_reg[908] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[877]$_DFFE_PN0P_  (.D(_0862_),
    .Q(\rf_reg[909] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[878]$_DFFE_PN0P_  (.D(_0863_),
    .Q(\rf_reg[910] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[879]$_DFFE_PN0P_  (.D(_0864_),
    .Q(\rf_reg[911] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[87]$_DFFE_PN0P_  (.D(_0865_),
    .Q(\rf_reg[119] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[880]$_DFFE_PN0P_  (.D(_0866_),
    .Q(\rf_reg[912] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[881]$_DFFE_PN0P_  (.D(_0867_),
    .Q(\rf_reg[913] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[882]$_DFFE_PN0P_  (.D(_0868_),
    .Q(\rf_reg[914] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[883]$_DFFE_PN0P_  (.D(_0869_),
    .Q(\rf_reg[915] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[884]$_DFFE_PN0P_  (.D(_0870_),
    .Q(\rf_reg[916] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[885]$_DFFE_PN0P_  (.D(_0871_),
    .Q(\rf_reg[917] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[886]$_DFFE_PN0P_  (.D(_0872_),
    .Q(\rf_reg[918] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[887]$_DFFE_PN0P_  (.D(_0873_),
    .Q(\rf_reg[919] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[888]$_DFFE_PN0P_  (.D(_0874_),
    .Q(\rf_reg[920] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[889]$_DFFE_PN0P_  (.D(_0875_),
    .Q(\rf_reg[921] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[88]$_DFFE_PN0P_  (.D(_0876_),
    .Q(\rf_reg[120] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[890]$_DFFE_PN0P_  (.D(_0877_),
    .Q(\rf_reg[922] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[891]$_DFFE_PN0P_  (.D(_0878_),
    .Q(\rf_reg[923] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[892]$_DFFE_PN0P_  (.D(_0879_),
    .Q(\rf_reg[924] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[893]$_DFFE_PN0P_  (.D(_0880_),
    .Q(\rf_reg[925] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[894]$_DFFE_PN0P_  (.D(_0881_),
    .Q(\rf_reg[926] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[895]$_DFFE_PN0P_  (.D(_0882_),
    .Q(\rf_reg[927] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[896]$_DFFE_PN0P_  (.D(_0883_),
    .Q(\rf_reg[928] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[897]$_DFFE_PN0P_  (.D(_0884_),
    .Q(\rf_reg[929] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[898]$_DFFE_PN0P_  (.D(_0885_),
    .Q(\rf_reg[930] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[899]$_DFFE_PN0P_  (.D(_0886_),
    .Q(\rf_reg[931] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[89]$_DFFE_PN0P_  (.D(_0887_),
    .Q(\rf_reg[121] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[8]$_DFFE_PN0P_  (.D(_0888_),
    .Q(\rf_reg[40] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[900]$_DFFE_PN0P_  (.D(_0889_),
    .Q(\rf_reg[932] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[901]$_DFFE_PN0P_  (.D(_0890_),
    .Q(\rf_reg[933] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[902]$_DFFE_PN0P_  (.D(_0891_),
    .Q(\rf_reg[934] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[903]$_DFFE_PN0P_  (.D(_0892_),
    .Q(\rf_reg[935] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[904]$_DFFE_PN0P_  (.D(_0893_),
    .Q(\rf_reg[936] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[905]$_DFFE_PN0P_  (.D(_0894_),
    .Q(\rf_reg[937] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[906]$_DFFE_PN0P_  (.D(_0895_),
    .Q(\rf_reg[938] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[907]$_DFFE_PN0P_  (.D(_0896_),
    .Q(\rf_reg[939] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[908]$_DFFE_PN0P_  (.D(_0897_),
    .Q(\rf_reg[940] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[909]$_DFFE_PN0P_  (.D(_0898_),
    .Q(\rf_reg[941] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[90]$_DFFE_PN0P_  (.D(_0899_),
    .Q(\rf_reg[122] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[910]$_DFFE_PN0P_  (.D(_0900_),
    .Q(\rf_reg[942] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[911]$_DFFE_PN0P_  (.D(_0901_),
    .Q(\rf_reg[943] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[912]$_DFFE_PN0P_  (.D(_0902_),
    .Q(\rf_reg[944] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[913]$_DFFE_PN0P_  (.D(_0903_),
    .Q(\rf_reg[945] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[914]$_DFFE_PN0P_  (.D(_0904_),
    .Q(\rf_reg[946] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[915]$_DFFE_PN0P_  (.D(_0905_),
    .Q(\rf_reg[947] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[916]$_DFFE_PN0P_  (.D(_0906_),
    .Q(\rf_reg[948] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[917]$_DFFE_PN0P_  (.D(_0907_),
    .Q(\rf_reg[949] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[918]$_DFFE_PN0P_  (.D(_0908_),
    .Q(\rf_reg[950] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[919]$_DFFE_PN0P_  (.D(_0909_),
    .Q(\rf_reg[951] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[91]$_DFFE_PN0P_  (.D(_0910_),
    .Q(\rf_reg[123] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[920]$_DFFE_PN0P_  (.D(_0911_),
    .Q(\rf_reg[952] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[921]$_DFFE_PN0P_  (.D(_0912_),
    .Q(\rf_reg[953] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[922]$_DFFE_PN0P_  (.D(_0913_),
    .Q(\rf_reg[954] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[923]$_DFFE_PN0P_  (.D(_0914_),
    .Q(\rf_reg[955] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[924]$_DFFE_PN0P_  (.D(_0915_),
    .Q(\rf_reg[956] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[925]$_DFFE_PN0P_  (.D(_0916_),
    .Q(\rf_reg[957] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[926]$_DFFE_PN0P_  (.D(_0917_),
    .Q(\rf_reg[958] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[927]$_DFFE_PN0P_  (.D(_0918_),
    .Q(\rf_reg[959] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[928]$_DFFE_PN0P_  (.D(_0919_),
    .Q(\rf_reg[960] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[929]$_DFFE_PN0P_  (.D(_0920_),
    .Q(\rf_reg[961] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[92]$_DFFE_PN0P_  (.D(_0921_),
    .Q(\rf_reg[124] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[930]$_DFFE_PN0P_  (.D(_0922_),
    .Q(\rf_reg[962] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[931]$_DFFE_PN0P_  (.D(_0923_),
    .Q(\rf_reg[963] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[932]$_DFFE_PN0P_  (.D(_0924_),
    .Q(\rf_reg[964] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[933]$_DFFE_PN0P_  (.D(_0925_),
    .Q(\rf_reg[965] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[934]$_DFFE_PN0P_  (.D(_0926_),
    .Q(\rf_reg[966] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[935]$_DFFE_PN0P_  (.D(_0927_),
    .Q(\rf_reg[967] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[936]$_DFFE_PN0P_  (.D(_0928_),
    .Q(\rf_reg[968] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[937]$_DFFE_PN0P_  (.D(_0929_),
    .Q(\rf_reg[969] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[938]$_DFFE_PN0P_  (.D(_0930_),
    .Q(\rf_reg[970] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[939]$_DFFE_PN0P_  (.D(_0931_),
    .Q(\rf_reg[971] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[93]$_DFFE_PN0P_  (.D(_0932_),
    .Q(\rf_reg[125] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[940]$_DFFE_PN0P_  (.D(_0933_),
    .Q(\rf_reg[972] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[941]$_DFFE_PN0P_  (.D(_0934_),
    .Q(\rf_reg[973] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[942]$_DFFE_PN0P_  (.D(_0935_),
    .Q(\rf_reg[974] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[943]$_DFFE_PN0P_  (.D(_0936_),
    .Q(\rf_reg[975] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[944]$_DFFE_PN0P_  (.D(_0937_),
    .Q(\rf_reg[976] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[945]$_DFFE_PN0P_  (.D(_0938_),
    .Q(\rf_reg[977] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[946]$_DFFE_PN0P_  (.D(_0939_),
    .Q(\rf_reg[978] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[947]$_DFFE_PN0P_  (.D(_0940_),
    .Q(\rf_reg[979] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[948]$_DFFE_PN0P_  (.D(_0941_),
    .Q(\rf_reg[980] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[949]$_DFFE_PN0P_  (.D(_0942_),
    .Q(\rf_reg[981] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[94]$_DFFE_PN0P_  (.D(_0943_),
    .Q(\rf_reg[126] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[950]$_DFFE_PN0P_  (.D(_0944_),
    .Q(\rf_reg[982] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[951]$_DFFE_PN0P_  (.D(_0945_),
    .Q(\rf_reg[983] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[952]$_DFFE_PN0P_  (.D(_0946_),
    .Q(\rf_reg[984] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[953]$_DFFE_PN0P_  (.D(_0947_),
    .Q(\rf_reg[985] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[954]$_DFFE_PN0P_  (.D(_0948_),
    .Q(\rf_reg[986] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[955]$_DFFE_PN0P_  (.D(_0949_),
    .Q(\rf_reg[987] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[956]$_DFFE_PN0P_  (.D(_0950_),
    .Q(\rf_reg[988] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[957]$_DFFE_PN0P_  (.D(_0951_),
    .Q(\rf_reg[989] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[958]$_DFFE_PN0P_  (.D(_0952_),
    .Q(\rf_reg[990] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[959]$_DFFE_PN0P_  (.D(_0953_),
    .Q(\rf_reg[991] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[95]$_DFFE_PN0P_  (.D(_0954_),
    .Q(\rf_reg[127] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[960]$_DFFE_PN0P_  (.D(_0955_),
    .Q(\rf_reg[992] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[961]$_DFFE_PN0P_  (.D(_0956_),
    .Q(\rf_reg[993] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[962]$_DFFE_PN0P_  (.D(_0957_),
    .Q(\rf_reg[994] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[963]$_DFFE_PN0P_  (.D(_0958_),
    .Q(\rf_reg[995] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[964]$_DFFE_PN0P_  (.D(_0959_),
    .Q(\rf_reg[996] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[965]$_DFFE_PN0P_  (.D(_0960_),
    .Q(\rf_reg[997] ),
    .RESET_B(net10),
    .CLK(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[966]$_DFFE_PN0P_  (.D(_0961_),
    .Q(\rf_reg[998] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[967]$_DFFE_PN0P_  (.D(_0962_),
    .Q(\rf_reg[999] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[968]$_DFFE_PN0P_  (.D(_0963_),
    .Q(\rf_reg[1000] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[969]$_DFFE_PN0P_  (.D(_0964_),
    .Q(\rf_reg[1001] ),
    .RESET_B(net15),
    .CLK(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[96]$_DFFE_PN0P_  (.D(_0965_),
    .Q(\rf_reg[128] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[970]$_DFFE_PN0P_  (.D(_0966_),
    .Q(\rf_reg[1002] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[971]$_DFFE_PN0P_  (.D(_0967_),
    .Q(\rf_reg[1003] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[972]$_DFFE_PN0P_  (.D(_0968_),
    .Q(\rf_reg[1004] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[973]$_DFFE_PN0P_  (.D(_0969_),
    .Q(\rf_reg[1005] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[974]$_DFFE_PN0P_  (.D(_0970_),
    .Q(\rf_reg[1006] ),
    .RESET_B(net2),
    .CLK(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[975]$_DFFE_PN0P_  (.D(_0971_),
    .Q(\rf_reg[1007] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[976]$_DFFE_PN0P_  (.D(_0972_),
    .Q(\rf_reg[1008] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[977]$_DFFE_PN0P_  (.D(_0973_),
    .Q(\rf_reg[1009] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[978]$_DFFE_PN0P_  (.D(_0974_),
    .Q(\rf_reg[1010] ),
    .RESET_B(net14),
    .CLK(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[979]$_DFFE_PN0P_  (.D(_0975_),
    .Q(\rf_reg[1011] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[97]$_DFFE_PN0P_  (.D(_0976_),
    .Q(\rf_reg[129] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[980]$_DFFE_PN0P_  (.D(_0977_),
    .Q(\rf_reg[1012] ),
    .RESET_B(net12),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[981]$_DFFE_PN0P_  (.D(_0978_),
    .Q(\rf_reg[1013] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[982]$_DFFE_PN0P_  (.D(_0979_),
    .Q(\rf_reg[1014] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[983]$_DFFE_PN0P_  (.D(_0980_),
    .Q(\rf_reg[1015] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[984]$_DFFE_PN0P_  (.D(_0981_),
    .Q(\rf_reg[1016] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[985]$_DFFE_PN0P_  (.D(_0982_),
    .Q(\rf_reg[1017] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[986]$_DFFE_PN0P_  (.D(_0983_),
    .Q(\rf_reg[1018] ),
    .RESET_B(net11),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[987]$_DFFE_PN0P_  (.D(_0984_),
    .Q(\rf_reg[1019] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[988]$_DFFE_PN0P_  (.D(_0985_),
    .Q(\rf_reg[1020] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[989]$_DFFE_PN0P_  (.D(_0986_),
    .Q(\rf_reg[1021] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[98]$_DFFE_PN0P_  (.D(_0987_),
    .Q(\rf_reg[130] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[990]$_DFFE_PN0P_  (.D(_0988_),
    .Q(\rf_reg[1022] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[991]$_DFFE_PN0P_  (.D(_0989_),
    .Q(\rf_reg[1023] ),
    .RESET_B(net8),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[99]$_DFFE_PN0P_  (.D(_0990_),
    .Q(\rf_reg[131] ),
    .RESET_B(net9),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \rf_reg_q[9]$_DFFE_PN0P_  (.D(_0991_),
    .Q(\rf_reg[41] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2324 ();
 sky130_fd_sc_hd__clkbuf_16 load_slew8 (.A(net9),
    .X(net8));
 sky130_fd_sc_hd__buf_16 load_slew9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 load_slew10 (.A(net13),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 load_slew11 (.A(net12),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 load_slew12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_16 max_length13 (.A(net15),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_16 load_slew14 (.A(net2),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_16 load_slew15 (.A(net2),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input1 (.A(raddr_b_i[3]),
    .X(net1));
 sky130_fd_sc_hd__buf_16 input2 (.A(rst_ni),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(waddr_a_i[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(waddr_a_i[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(waddr_a_i[4]),
    .X(net5));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input6 (.A(wdata_a_i[0]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(wdata_a_i[10]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(wdata_a_i[11]),
    .X(net16));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input9 (.A(wdata_a_i[12]),
    .X(net17));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input10 (.A(wdata_a_i[13]),
    .X(net18));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input11 (.A(wdata_a_i[14]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input12 (.A(wdata_a_i[15]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input13 (.A(wdata_a_i[16]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input14 (.A(wdata_a_i[17]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input15 (.A(wdata_a_i[18]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input16 (.A(wdata_a_i[19]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input17 (.A(wdata_a_i[1]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input18 (.A(wdata_a_i[20]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input19 (.A(wdata_a_i[21]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input20 (.A(wdata_a_i[22]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input21 (.A(wdata_a_i[23]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input22 (.A(wdata_a_i[24]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input23 (.A(wdata_a_i[25]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input24 (.A(wdata_a_i[26]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input25 (.A(wdata_a_i[27]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input26 (.A(wdata_a_i[28]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input27 (.A(wdata_a_i[29]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input28 (.A(wdata_a_i[2]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input29 (.A(wdata_a_i[30]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input30 (.A(wdata_a_i[31]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input31 (.A(wdata_a_i[3]),
    .X(net39));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input32 (.A(wdata_a_i[4]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input33 (.A(wdata_a_i[5]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input34 (.A(wdata_a_i[6]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input35 (.A(wdata_a_i[7]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input36 (.A(wdata_a_i[8]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input37 (.A(wdata_a_i[9]),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input38 (.A(we_a_i),
    .X(net46));
 sky130_fd_sc_hd__buf_1 output39 (.A(net47),
    .X(rdata_a_o[0]));
 sky130_fd_sc_hd__buf_1 output40 (.A(net48),
    .X(rdata_a_o[10]));
 sky130_fd_sc_hd__buf_1 output41 (.A(net49),
    .X(rdata_a_o[11]));
 sky130_fd_sc_hd__buf_1 output42 (.A(net50),
    .X(rdata_a_o[12]));
 sky130_fd_sc_hd__buf_1 output43 (.A(net51),
    .X(rdata_a_o[13]));
 sky130_fd_sc_hd__buf_1 output44 (.A(net52),
    .X(rdata_a_o[14]));
 sky130_fd_sc_hd__buf_1 output45 (.A(net53),
    .X(rdata_a_o[15]));
 sky130_fd_sc_hd__buf_1 output46 (.A(net54),
    .X(rdata_a_o[16]));
 sky130_fd_sc_hd__buf_1 output47 (.A(net55),
    .X(rdata_a_o[17]));
 sky130_fd_sc_hd__buf_1 output48 (.A(net56),
    .X(rdata_a_o[18]));
 sky130_fd_sc_hd__buf_1 output49 (.A(net57),
    .X(rdata_a_o[19]));
 sky130_fd_sc_hd__buf_1 output50 (.A(net58),
    .X(rdata_a_o[1]));
 sky130_fd_sc_hd__buf_1 output51 (.A(net59),
    .X(rdata_a_o[20]));
 sky130_fd_sc_hd__buf_1 output52 (.A(net60),
    .X(rdata_a_o[21]));
 sky130_fd_sc_hd__buf_1 output53 (.A(net61),
    .X(rdata_a_o[22]));
 sky130_fd_sc_hd__buf_1 output54 (.A(net62),
    .X(rdata_a_o[23]));
 sky130_fd_sc_hd__buf_1 output55 (.A(net63),
    .X(rdata_a_o[24]));
 sky130_fd_sc_hd__buf_1 output56 (.A(net64),
    .X(rdata_a_o[25]));
 sky130_fd_sc_hd__buf_1 output57 (.A(net65),
    .X(rdata_a_o[26]));
 sky130_fd_sc_hd__buf_1 output58 (.A(net66),
    .X(rdata_a_o[27]));
 sky130_fd_sc_hd__buf_1 output59 (.A(net67),
    .X(rdata_a_o[28]));
 sky130_fd_sc_hd__buf_1 output60 (.A(net68),
    .X(rdata_a_o[29]));
 sky130_fd_sc_hd__buf_1 output61 (.A(net69),
    .X(rdata_a_o[2]));
 sky130_fd_sc_hd__buf_1 output62 (.A(net70),
    .X(rdata_a_o[30]));
 sky130_fd_sc_hd__buf_1 output63 (.A(net71),
    .X(rdata_a_o[31]));
 sky130_fd_sc_hd__buf_1 output64 (.A(net72),
    .X(rdata_a_o[3]));
 sky130_fd_sc_hd__buf_1 output65 (.A(net73),
    .X(rdata_a_o[4]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net74),
    .X(rdata_a_o[5]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net75),
    .X(rdata_a_o[6]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net76),
    .X(rdata_a_o[7]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net77),
    .X(rdata_a_o[8]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net78),
    .X(rdata_a_o[9]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net79),
    .X(rdata_b_o[0]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net80),
    .X(rdata_b_o[10]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net81),
    .X(rdata_b_o[11]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net82),
    .X(rdata_b_o[12]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net83),
    .X(rdata_b_o[13]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net84),
    .X(rdata_b_o[14]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net85),
    .X(rdata_b_o[15]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net86),
    .X(rdata_b_o[16]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net87),
    .X(rdata_b_o[17]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net88),
    .X(rdata_b_o[18]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net89),
    .X(rdata_b_o[19]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net90),
    .X(rdata_b_o[1]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net91),
    .X(rdata_b_o[20]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net92),
    .X(rdata_b_o[21]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net93),
    .X(rdata_b_o[22]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net94),
    .X(rdata_b_o[23]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net95),
    .X(rdata_b_o[24]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net96),
    .X(rdata_b_o[25]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net97),
    .X(rdata_b_o[26]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net98),
    .X(rdata_b_o[27]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net99),
    .X(rdata_b_o[28]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net100),
    .X(rdata_b_o[29]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net101),
    .X(rdata_b_o[2]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net102),
    .X(rdata_b_o[30]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net103),
    .X(rdata_b_o[31]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net104),
    .X(rdata_b_o[3]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net105),
    .X(rdata_b_o[4]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net106),
    .X(rdata_b_o[5]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net107),
    .X(rdata_b_o[6]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net108),
    .X(rdata_b_o[7]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net109),
    .X(rdata_b_o[8]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net110),
    .X(rdata_b_o[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i (.A(clknet_3_2__leaf_clk_i),
    .X(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_i (.A(clknet_3_3__leaf_clk_i),
    .X(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_i (.A(clknet_3_7__leaf_clk_i),
    .X(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_i (.A(clknet_3_6__leaf_clk_i),
    .X(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_i (.A(clknet_3_5__leaf_clk_i),
    .X(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_i (.A(clknet_3_4__leaf_clk_i),
    .X(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk_i (.A(clknet_3_1__leaf_clk_i),
    .X(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk_i (.A(clknet_3_0__leaf_clk_i),
    .X(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkload0 (.A(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkload1 (.A(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__clkinv_16 clkload3 (.A(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkload4 (.A(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload6 (.A(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload7 (.A(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload8 (.A(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload9 (.A(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload10 (.A(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload11 (.A(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload13 (.A(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload14 (.A(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload15 (.A(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__inv_6 clkload16 (.A(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload17 (.A(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload18 (.A(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload19 (.A(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload20 (.A(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload21 (.A(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload22 (.A(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload23 (.A(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload24 (.A(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload25 (.A(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload26 (.A(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload27 (.A(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload28 (.A(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload29 (.A(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload30 (.A(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload31 (.A(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload32 (.A(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload33 (.A(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload34 (.A(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload35 (.A(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload36 (.A(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload37 (.A(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload38 (.A(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload39 (.A(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload40 (.A(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload41 (.A(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload43 (.A(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload45 (.A(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload46 (.A(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload47 (.A(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload48 (.A(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload49 (.A(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload50 (.A(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload51 (.A(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload52 (.A(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload53 (.A(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload54 (.A(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__clkinvlp_4 clkload55 (.A(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload56 (.A(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload57 (.A(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload58 (.A(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload59 (.A(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload60 (.A(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload61 (.A(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload63 (.A(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__inv_6 clkload64 (.A(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload65 (.A(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload66 (.A(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload67 (.A(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload68 (.A(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload69 (.A(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload70 (.A(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload71 (.A(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload72 (.A(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload73 (.A(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload74 (.A(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload75 (.A(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload76 (.A(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload77 (.A(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload78 (.A(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload79 (.A(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload80 (.A(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload81 (.A(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload82 (.A(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload83 (.A(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload84 (.A(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload85 (.A(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload86 (.A(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload87 (.A(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload88 (.A(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload89 (.A(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload90 (.A(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload91 (.A(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload92 (.A(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_654 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_774 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_632 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_844 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_850 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_902 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_803 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_911 ();
endmodule
