VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA ibex_register_file_ff_via2_3_1600_480_1_5_320_320
  VIARULE M1M2_PR ;
  CUTSIZE 0.15 0.15 ;
  LAYERS met1 via met2 ;
  CUTSPACING 0.17 0.17 ;
  ENCLOSURE 0.085 0.165 0.055 0.085 ;
  ROWCOL 1 5 ;
END ibex_register_file_ff_via2_3_1600_480_1_5_320_320

VIA ibex_register_file_ff_via3_4_1600_480_1_4_400_400
  VIARULE M2M3_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met2 via2 met3 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.04 0.085 0.065 0.065 ;
  ROWCOL 1 4 ;
END ibex_register_file_ff_via3_4_1600_480_1_4_400_400

VIA ibex_register_file_ff_via4_5_1600_480_1_4_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.06 0.1 0.065 ;
  ROWCOL 1 4 ;
END ibex_register_file_ff_via4_5_1600_480_1_4_400_400

VIA ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600
  VIARULE M4M5_PR ;
  CUTSIZE 0.8 0.8 ;
  LAYERS met4 via4 met5 ;
  CUTSPACING 0.8 0.8 ;
  ENCLOSURE 0.4 0.19 0.31 0.4 ;
END ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600

MACRO ibex_register_file_ff
  FOREIGN ibex_register_file_ff 0 0 ;
  CLASS BLOCK ;
  SIZE 421.97 BY 421.97 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  27.72 409.92 409.28 411.52 ;
        RECT  27.72 382.72 409.28 384.32 ;
        RECT  27.72 355.52 409.28 357.12 ;
        RECT  27.72 328.32 409.28 329.92 ;
        RECT  27.72 301.12 409.28 302.72 ;
        RECT  27.72 273.92 409.28 275.52 ;
        RECT  27.72 246.72 409.28 248.32 ;
        RECT  27.72 219.52 409.28 221.12 ;
        RECT  27.72 192.32 409.28 193.92 ;
        RECT  27.72 165.12 409.28 166.72 ;
        RECT  27.72 137.92 409.28 139.52 ;
        RECT  27.72 110.72 409.28 112.32 ;
        RECT  27.72 83.52 409.28 85.12 ;
        RECT  27.72 56.32 409.28 57.92 ;
        RECT  27.72 29.12 409.28 30.72 ;
      LAYER met4 ;
        RECT  407.68 5.2 409.28 419.12 ;
        RECT  380.54 5.2 382.14 419.12 ;
        RECT  353.4 5.2 355 419.12 ;
        RECT  326.26 5.2 327.86 419.12 ;
        RECT  299.12 5.2 300.72 419.12 ;
        RECT  271.98 5.2 273.58 419.12 ;
        RECT  244.84 5.2 246.44 419.12 ;
        RECT  217.7 5.2 219.3 419.12 ;
        RECT  190.56 5.2 192.16 419.12 ;
        RECT  163.42 5.2 165.02 419.12 ;
        RECT  136.28 5.2 137.88 419.12 ;
        RECT  109.14 5.2 110.74 419.12 ;
        RECT  82 5.2 83.6 419.12 ;
        RECT  54.86 5.2 56.46 419.12 ;
        RECT  27.72 5.2 29.32 419.12 ;
      LAYER met1 ;
        RECT  1.38 418.64 420.9 419.12 ;
        RECT  1.38 413.2 420.9 413.68 ;
        RECT  1.38 407.76 420.9 408.24 ;
        RECT  1.38 402.32 420.9 402.8 ;
        RECT  1.38 396.88 420.9 397.36 ;
        RECT  1.38 391.44 420.9 391.92 ;
        RECT  1.38 386 420.9 386.48 ;
        RECT  1.38 380.56 420.9 381.04 ;
        RECT  1.38 375.12 420.9 375.6 ;
        RECT  1.38 369.68 420.9 370.16 ;
        RECT  1.38 364.24 420.9 364.72 ;
        RECT  1.38 358.8 420.9 359.28 ;
        RECT  1.38 353.36 420.9 353.84 ;
        RECT  1.38 347.92 420.9 348.4 ;
        RECT  1.38 342.48 420.9 342.96 ;
        RECT  1.38 337.04 420.9 337.52 ;
        RECT  1.38 331.6 420.9 332.08 ;
        RECT  1.38 326.16 420.9 326.64 ;
        RECT  1.38 320.72 420.9 321.2 ;
        RECT  1.38 315.28 420.9 315.76 ;
        RECT  1.38 309.84 420.9 310.32 ;
        RECT  1.38 304.4 420.9 304.88 ;
        RECT  1.38 298.96 420.9 299.44 ;
        RECT  1.38 293.52 420.9 294 ;
        RECT  1.38 288.08 420.9 288.56 ;
        RECT  1.38 282.64 420.9 283.12 ;
        RECT  1.38 277.2 420.9 277.68 ;
        RECT  1.38 271.76 420.9 272.24 ;
        RECT  1.38 266.32 420.9 266.8 ;
        RECT  1.38 260.88 420.9 261.36 ;
        RECT  1.38 255.44 420.9 255.92 ;
        RECT  1.38 250 420.9 250.48 ;
        RECT  1.38 244.56 420.9 245.04 ;
        RECT  1.38 239.12 420.9 239.6 ;
        RECT  1.38 233.68 420.9 234.16 ;
        RECT  1.38 228.24 420.9 228.72 ;
        RECT  1.38 222.8 420.9 223.28 ;
        RECT  1.38 217.36 420.9 217.84 ;
        RECT  1.38 211.92 420.9 212.4 ;
        RECT  1.38 206.48 420.9 206.96 ;
        RECT  1.38 201.04 420.9 201.52 ;
        RECT  1.38 195.6 420.9 196.08 ;
        RECT  1.38 190.16 420.9 190.64 ;
        RECT  1.38 184.72 420.9 185.2 ;
        RECT  1.38 179.28 420.9 179.76 ;
        RECT  1.38 173.84 420.9 174.32 ;
        RECT  1.38 168.4 420.9 168.88 ;
        RECT  1.38 162.96 420.9 163.44 ;
        RECT  1.38 157.52 420.9 158 ;
        RECT  1.38 152.08 420.9 152.56 ;
        RECT  1.38 146.64 420.9 147.12 ;
        RECT  1.38 141.2 420.9 141.68 ;
        RECT  1.38 135.76 420.9 136.24 ;
        RECT  1.38 130.32 420.9 130.8 ;
        RECT  1.38 124.88 420.9 125.36 ;
        RECT  1.38 119.44 420.9 119.92 ;
        RECT  1.38 114 420.9 114.48 ;
        RECT  1.38 108.56 420.9 109.04 ;
        RECT  1.38 103.12 420.9 103.6 ;
        RECT  1.38 97.68 420.9 98.16 ;
        RECT  1.38 92.24 420.9 92.72 ;
        RECT  1.38 86.8 420.9 87.28 ;
        RECT  1.38 81.36 420.9 81.84 ;
        RECT  1.38 75.92 420.9 76.4 ;
        RECT  1.38 70.48 420.9 70.96 ;
        RECT  1.38 65.04 420.9 65.52 ;
        RECT  1.38 59.6 420.9 60.08 ;
        RECT  1.38 54.16 420.9 54.64 ;
        RECT  1.38 48.72 420.9 49.2 ;
        RECT  1.38 43.28 420.9 43.76 ;
        RECT  1.38 37.84 420.9 38.32 ;
        RECT  1.38 32.4 420.9 32.88 ;
        RECT  1.38 26.96 420.9 27.44 ;
        RECT  1.38 21.52 420.9 22 ;
        RECT  1.38 16.08 420.9 16.56 ;
        RECT  1.38 10.64 420.9 11.12 ;
        RECT  1.38 5.2 420.9 5.68 ;
      VIA 408.48 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 408.48 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 381.34 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 354.2 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 327.06 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 299.92 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 410.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 383.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 356.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 329.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 301.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 274.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 247.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 220.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 193.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 165.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 138.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 111.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 84.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 57.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 29.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  407.69 418.715 409.27 419.045 ;
      VIA 408.48 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 418.695 409.25 419.065 ;
      VIA 408.48 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 413.275 409.27 413.605 ;
      VIA 408.48 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 413.255 409.25 413.625 ;
      VIA 408.48 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 407.835 409.27 408.165 ;
      VIA 408.48 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 407.815 409.25 408.185 ;
      VIA 408.48 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 402.395 409.27 402.725 ;
      VIA 408.48 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 402.375 409.25 402.745 ;
      VIA 408.48 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 396.955 409.27 397.285 ;
      VIA 408.48 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 396.935 409.25 397.305 ;
      VIA 408.48 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 391.515 409.27 391.845 ;
      VIA 408.48 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 391.495 409.25 391.865 ;
      VIA 408.48 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 386.075 409.27 386.405 ;
      VIA 408.48 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 386.055 409.25 386.425 ;
      VIA 408.48 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 380.635 409.27 380.965 ;
      VIA 408.48 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 380.615 409.25 380.985 ;
      VIA 408.48 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 375.195 409.27 375.525 ;
      VIA 408.48 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 375.175 409.25 375.545 ;
      VIA 408.48 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 369.755 409.27 370.085 ;
      VIA 408.48 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 369.735 409.25 370.105 ;
      VIA 408.48 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 364.315 409.27 364.645 ;
      VIA 408.48 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 364.295 409.25 364.665 ;
      VIA 408.48 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 358.875 409.27 359.205 ;
      VIA 408.48 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 358.855 409.25 359.225 ;
      VIA 408.48 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 353.435 409.27 353.765 ;
      VIA 408.48 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 353.415 409.25 353.785 ;
      VIA 408.48 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 347.995 409.27 348.325 ;
      VIA 408.48 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 347.975 409.25 348.345 ;
      VIA 408.48 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 342.555 409.27 342.885 ;
      VIA 408.48 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 342.535 409.25 342.905 ;
      VIA 408.48 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 337.115 409.27 337.445 ;
      VIA 408.48 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 337.095 409.25 337.465 ;
      VIA 408.48 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 331.675 409.27 332.005 ;
      VIA 408.48 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 331.655 409.25 332.025 ;
      VIA 408.48 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 326.235 409.27 326.565 ;
      VIA 408.48 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 326.215 409.25 326.585 ;
      VIA 408.48 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 320.795 409.27 321.125 ;
      VIA 408.48 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 320.775 409.25 321.145 ;
      VIA 408.48 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 315.355 409.27 315.685 ;
      VIA 408.48 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 315.335 409.25 315.705 ;
      VIA 408.48 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 309.915 409.27 310.245 ;
      VIA 408.48 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 309.895 409.25 310.265 ;
      VIA 408.48 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 304.475 409.27 304.805 ;
      VIA 408.48 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 304.455 409.25 304.825 ;
      VIA 408.48 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 299.035 409.27 299.365 ;
      VIA 408.48 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 299.015 409.25 299.385 ;
      VIA 408.48 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 293.595 409.27 293.925 ;
      VIA 408.48 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 293.575 409.25 293.945 ;
      VIA 408.48 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 288.155 409.27 288.485 ;
      VIA 408.48 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 288.135 409.25 288.505 ;
      VIA 408.48 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 282.715 409.27 283.045 ;
      VIA 408.48 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 282.695 409.25 283.065 ;
      VIA 408.48 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 277.275 409.27 277.605 ;
      VIA 408.48 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 277.255 409.25 277.625 ;
      VIA 408.48 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 271.835 409.27 272.165 ;
      VIA 408.48 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 271.815 409.25 272.185 ;
      VIA 408.48 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 266.395 409.27 266.725 ;
      VIA 408.48 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 266.375 409.25 266.745 ;
      VIA 408.48 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 260.955 409.27 261.285 ;
      VIA 408.48 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 260.935 409.25 261.305 ;
      VIA 408.48 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 255.515 409.27 255.845 ;
      VIA 408.48 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 255.495 409.25 255.865 ;
      VIA 408.48 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 250.075 409.27 250.405 ;
      VIA 408.48 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 250.055 409.25 250.425 ;
      VIA 408.48 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 244.635 409.27 244.965 ;
      VIA 408.48 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 244.615 409.25 244.985 ;
      VIA 408.48 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 239.195 409.27 239.525 ;
      VIA 408.48 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 239.175 409.25 239.545 ;
      VIA 408.48 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 233.755 409.27 234.085 ;
      VIA 408.48 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 233.735 409.25 234.105 ;
      VIA 408.48 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 228.315 409.27 228.645 ;
      VIA 408.48 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 228.295 409.25 228.665 ;
      VIA 408.48 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 222.875 409.27 223.205 ;
      VIA 408.48 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 222.855 409.25 223.225 ;
      VIA 408.48 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 217.435 409.27 217.765 ;
      VIA 408.48 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 217.415 409.25 217.785 ;
      VIA 408.48 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 211.995 409.27 212.325 ;
      VIA 408.48 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 211.975 409.25 212.345 ;
      VIA 408.48 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 206.555 409.27 206.885 ;
      VIA 408.48 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 206.535 409.25 206.905 ;
      VIA 408.48 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 201.115 409.27 201.445 ;
      VIA 408.48 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 201.095 409.25 201.465 ;
      VIA 408.48 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 195.675 409.27 196.005 ;
      VIA 408.48 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 195.655 409.25 196.025 ;
      VIA 408.48 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 190.235 409.27 190.565 ;
      VIA 408.48 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 190.215 409.25 190.585 ;
      VIA 408.48 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 184.795 409.27 185.125 ;
      VIA 408.48 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 184.775 409.25 185.145 ;
      VIA 408.48 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 179.355 409.27 179.685 ;
      VIA 408.48 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 179.335 409.25 179.705 ;
      VIA 408.48 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 173.915 409.27 174.245 ;
      VIA 408.48 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 173.895 409.25 174.265 ;
      VIA 408.48 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 168.475 409.27 168.805 ;
      VIA 408.48 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 168.455 409.25 168.825 ;
      VIA 408.48 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 163.035 409.27 163.365 ;
      VIA 408.48 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 163.015 409.25 163.385 ;
      VIA 408.48 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 157.595 409.27 157.925 ;
      VIA 408.48 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 157.575 409.25 157.945 ;
      VIA 408.48 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 152.155 409.27 152.485 ;
      VIA 408.48 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 152.135 409.25 152.505 ;
      VIA 408.48 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 146.715 409.27 147.045 ;
      VIA 408.48 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 146.695 409.25 147.065 ;
      VIA 408.48 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 141.275 409.27 141.605 ;
      VIA 408.48 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 141.255 409.25 141.625 ;
      VIA 408.48 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 135.835 409.27 136.165 ;
      VIA 408.48 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 135.815 409.25 136.185 ;
      VIA 408.48 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 130.395 409.27 130.725 ;
      VIA 408.48 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 130.375 409.25 130.745 ;
      VIA 408.48 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 124.955 409.27 125.285 ;
      VIA 408.48 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 124.935 409.25 125.305 ;
      VIA 408.48 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 119.515 409.27 119.845 ;
      VIA 408.48 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 119.495 409.25 119.865 ;
      VIA 408.48 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 114.075 409.27 114.405 ;
      VIA 408.48 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 114.055 409.25 114.425 ;
      VIA 408.48 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 108.635 409.27 108.965 ;
      VIA 408.48 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 108.615 409.25 108.985 ;
      VIA 408.48 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 103.195 409.27 103.525 ;
      VIA 408.48 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 103.175 409.25 103.545 ;
      VIA 408.48 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 97.755 409.27 98.085 ;
      VIA 408.48 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 97.735 409.25 98.105 ;
      VIA 408.48 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 92.315 409.27 92.645 ;
      VIA 408.48 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 92.295 409.25 92.665 ;
      VIA 408.48 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 86.875 409.27 87.205 ;
      VIA 408.48 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 86.855 409.25 87.225 ;
      VIA 408.48 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 81.435 409.27 81.765 ;
      VIA 408.48 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 81.415 409.25 81.785 ;
      VIA 408.48 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 75.995 409.27 76.325 ;
      VIA 408.48 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 75.975 409.25 76.345 ;
      VIA 408.48 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 70.555 409.27 70.885 ;
      VIA 408.48 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 70.535 409.25 70.905 ;
      VIA 408.48 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 65.115 409.27 65.445 ;
      VIA 408.48 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 65.095 409.25 65.465 ;
      VIA 408.48 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 59.675 409.27 60.005 ;
      VIA 408.48 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 59.655 409.25 60.025 ;
      VIA 408.48 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 54.235 409.27 54.565 ;
      VIA 408.48 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 54.215 409.25 54.585 ;
      VIA 408.48 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 48.795 409.27 49.125 ;
      VIA 408.48 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 48.775 409.25 49.145 ;
      VIA 408.48 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 43.355 409.27 43.685 ;
      VIA 408.48 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 43.335 409.25 43.705 ;
      VIA 408.48 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 37.915 409.27 38.245 ;
      VIA 408.48 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 37.895 409.25 38.265 ;
      VIA 408.48 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 32.475 409.27 32.805 ;
      VIA 408.48 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 32.455 409.25 32.825 ;
      VIA 408.48 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 27.035 409.27 27.365 ;
      VIA 408.48 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 27.015 409.25 27.385 ;
      VIA 408.48 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 21.595 409.27 21.925 ;
      VIA 408.48 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 21.575 409.25 21.945 ;
      VIA 408.48 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 16.155 409.27 16.485 ;
      VIA 408.48 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 16.135 409.25 16.505 ;
      VIA 408.48 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 10.715 409.27 11.045 ;
      VIA 408.48 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 10.695 409.25 11.065 ;
      VIA 408.48 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  407.69 5.275 409.27 5.605 ;
      VIA 408.48 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  407.71 5.255 409.25 5.625 ;
      VIA 408.48 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 408.48 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 418.715 382.13 419.045 ;
      VIA 381.34 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 418.695 382.11 419.065 ;
      VIA 381.34 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 413.275 382.13 413.605 ;
      VIA 381.34 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 413.255 382.11 413.625 ;
      VIA 381.34 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 407.835 382.13 408.165 ;
      VIA 381.34 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 407.815 382.11 408.185 ;
      VIA 381.34 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 402.395 382.13 402.725 ;
      VIA 381.34 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 402.375 382.11 402.745 ;
      VIA 381.34 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 396.955 382.13 397.285 ;
      VIA 381.34 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 396.935 382.11 397.305 ;
      VIA 381.34 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 391.515 382.13 391.845 ;
      VIA 381.34 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 391.495 382.11 391.865 ;
      VIA 381.34 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 386.075 382.13 386.405 ;
      VIA 381.34 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 386.055 382.11 386.425 ;
      VIA 381.34 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 380.635 382.13 380.965 ;
      VIA 381.34 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 380.615 382.11 380.985 ;
      VIA 381.34 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 375.195 382.13 375.525 ;
      VIA 381.34 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 375.175 382.11 375.545 ;
      VIA 381.34 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 369.755 382.13 370.085 ;
      VIA 381.34 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 369.735 382.11 370.105 ;
      VIA 381.34 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 364.315 382.13 364.645 ;
      VIA 381.34 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 364.295 382.11 364.665 ;
      VIA 381.34 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 358.875 382.13 359.205 ;
      VIA 381.34 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 358.855 382.11 359.225 ;
      VIA 381.34 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 353.435 382.13 353.765 ;
      VIA 381.34 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 353.415 382.11 353.785 ;
      VIA 381.34 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 347.995 382.13 348.325 ;
      VIA 381.34 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 347.975 382.11 348.345 ;
      VIA 381.34 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 342.555 382.13 342.885 ;
      VIA 381.34 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 342.535 382.11 342.905 ;
      VIA 381.34 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 337.115 382.13 337.445 ;
      VIA 381.34 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 337.095 382.11 337.465 ;
      VIA 381.34 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 331.675 382.13 332.005 ;
      VIA 381.34 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 331.655 382.11 332.025 ;
      VIA 381.34 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 326.235 382.13 326.565 ;
      VIA 381.34 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 326.215 382.11 326.585 ;
      VIA 381.34 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 320.795 382.13 321.125 ;
      VIA 381.34 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 320.775 382.11 321.145 ;
      VIA 381.34 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 315.355 382.13 315.685 ;
      VIA 381.34 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 315.335 382.11 315.705 ;
      VIA 381.34 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 309.915 382.13 310.245 ;
      VIA 381.34 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 309.895 382.11 310.265 ;
      VIA 381.34 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 304.475 382.13 304.805 ;
      VIA 381.34 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 304.455 382.11 304.825 ;
      VIA 381.34 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 299.035 382.13 299.365 ;
      VIA 381.34 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 299.015 382.11 299.385 ;
      VIA 381.34 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 293.595 382.13 293.925 ;
      VIA 381.34 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 293.575 382.11 293.945 ;
      VIA 381.34 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 288.155 382.13 288.485 ;
      VIA 381.34 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 288.135 382.11 288.505 ;
      VIA 381.34 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 282.715 382.13 283.045 ;
      VIA 381.34 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 282.695 382.11 283.065 ;
      VIA 381.34 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 277.275 382.13 277.605 ;
      VIA 381.34 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 277.255 382.11 277.625 ;
      VIA 381.34 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 271.835 382.13 272.165 ;
      VIA 381.34 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 271.815 382.11 272.185 ;
      VIA 381.34 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 266.395 382.13 266.725 ;
      VIA 381.34 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 266.375 382.11 266.745 ;
      VIA 381.34 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 260.955 382.13 261.285 ;
      VIA 381.34 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 260.935 382.11 261.305 ;
      VIA 381.34 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 255.515 382.13 255.845 ;
      VIA 381.34 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 255.495 382.11 255.865 ;
      VIA 381.34 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 250.075 382.13 250.405 ;
      VIA 381.34 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 250.055 382.11 250.425 ;
      VIA 381.34 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 244.635 382.13 244.965 ;
      VIA 381.34 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 244.615 382.11 244.985 ;
      VIA 381.34 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 239.195 382.13 239.525 ;
      VIA 381.34 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 239.175 382.11 239.545 ;
      VIA 381.34 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 233.755 382.13 234.085 ;
      VIA 381.34 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 233.735 382.11 234.105 ;
      VIA 381.34 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 228.315 382.13 228.645 ;
      VIA 381.34 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 228.295 382.11 228.665 ;
      VIA 381.34 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 222.875 382.13 223.205 ;
      VIA 381.34 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 222.855 382.11 223.225 ;
      VIA 381.34 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 217.435 382.13 217.765 ;
      VIA 381.34 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 217.415 382.11 217.785 ;
      VIA 381.34 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 211.995 382.13 212.325 ;
      VIA 381.34 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 211.975 382.11 212.345 ;
      VIA 381.34 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 206.555 382.13 206.885 ;
      VIA 381.34 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 206.535 382.11 206.905 ;
      VIA 381.34 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 201.115 382.13 201.445 ;
      VIA 381.34 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 201.095 382.11 201.465 ;
      VIA 381.34 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 195.675 382.13 196.005 ;
      VIA 381.34 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 195.655 382.11 196.025 ;
      VIA 381.34 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 190.235 382.13 190.565 ;
      VIA 381.34 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 190.215 382.11 190.585 ;
      VIA 381.34 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 184.795 382.13 185.125 ;
      VIA 381.34 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 184.775 382.11 185.145 ;
      VIA 381.34 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 179.355 382.13 179.685 ;
      VIA 381.34 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 179.335 382.11 179.705 ;
      VIA 381.34 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 173.915 382.13 174.245 ;
      VIA 381.34 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 173.895 382.11 174.265 ;
      VIA 381.34 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 168.475 382.13 168.805 ;
      VIA 381.34 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 168.455 382.11 168.825 ;
      VIA 381.34 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 163.035 382.13 163.365 ;
      VIA 381.34 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 163.015 382.11 163.385 ;
      VIA 381.34 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 157.595 382.13 157.925 ;
      VIA 381.34 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 157.575 382.11 157.945 ;
      VIA 381.34 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 152.155 382.13 152.485 ;
      VIA 381.34 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 152.135 382.11 152.505 ;
      VIA 381.34 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 146.715 382.13 147.045 ;
      VIA 381.34 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 146.695 382.11 147.065 ;
      VIA 381.34 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 141.275 382.13 141.605 ;
      VIA 381.34 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 141.255 382.11 141.625 ;
      VIA 381.34 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 135.835 382.13 136.165 ;
      VIA 381.34 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 135.815 382.11 136.185 ;
      VIA 381.34 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 130.395 382.13 130.725 ;
      VIA 381.34 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 130.375 382.11 130.745 ;
      VIA 381.34 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 124.955 382.13 125.285 ;
      VIA 381.34 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 124.935 382.11 125.305 ;
      VIA 381.34 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 119.515 382.13 119.845 ;
      VIA 381.34 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 119.495 382.11 119.865 ;
      VIA 381.34 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 114.075 382.13 114.405 ;
      VIA 381.34 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 114.055 382.11 114.425 ;
      VIA 381.34 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 108.635 382.13 108.965 ;
      VIA 381.34 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 108.615 382.11 108.985 ;
      VIA 381.34 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 103.195 382.13 103.525 ;
      VIA 381.34 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 103.175 382.11 103.545 ;
      VIA 381.34 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 97.755 382.13 98.085 ;
      VIA 381.34 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 97.735 382.11 98.105 ;
      VIA 381.34 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 92.315 382.13 92.645 ;
      VIA 381.34 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 92.295 382.11 92.665 ;
      VIA 381.34 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 86.875 382.13 87.205 ;
      VIA 381.34 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 86.855 382.11 87.225 ;
      VIA 381.34 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 81.435 382.13 81.765 ;
      VIA 381.34 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 81.415 382.11 81.785 ;
      VIA 381.34 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 75.995 382.13 76.325 ;
      VIA 381.34 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 75.975 382.11 76.345 ;
      VIA 381.34 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 70.555 382.13 70.885 ;
      VIA 381.34 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 70.535 382.11 70.905 ;
      VIA 381.34 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 65.115 382.13 65.445 ;
      VIA 381.34 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 65.095 382.11 65.465 ;
      VIA 381.34 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 59.675 382.13 60.005 ;
      VIA 381.34 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 59.655 382.11 60.025 ;
      VIA 381.34 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 54.235 382.13 54.565 ;
      VIA 381.34 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 54.215 382.11 54.585 ;
      VIA 381.34 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 48.795 382.13 49.125 ;
      VIA 381.34 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 48.775 382.11 49.145 ;
      VIA 381.34 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 43.355 382.13 43.685 ;
      VIA 381.34 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 43.335 382.11 43.705 ;
      VIA 381.34 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 37.915 382.13 38.245 ;
      VIA 381.34 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 37.895 382.11 38.265 ;
      VIA 381.34 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 32.475 382.13 32.805 ;
      VIA 381.34 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 32.455 382.11 32.825 ;
      VIA 381.34 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 27.035 382.13 27.365 ;
      VIA 381.34 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 27.015 382.11 27.385 ;
      VIA 381.34 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 21.595 382.13 21.925 ;
      VIA 381.34 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 21.575 382.11 21.945 ;
      VIA 381.34 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 16.155 382.13 16.485 ;
      VIA 381.34 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 16.135 382.11 16.505 ;
      VIA 381.34 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 10.715 382.13 11.045 ;
      VIA 381.34 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 10.695 382.11 11.065 ;
      VIA 381.34 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  380.55 5.275 382.13 5.605 ;
      VIA 381.34 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  380.57 5.255 382.11 5.625 ;
      VIA 381.34 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 381.34 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 418.715 354.99 419.045 ;
      VIA 354.2 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 418.695 354.97 419.065 ;
      VIA 354.2 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 413.275 354.99 413.605 ;
      VIA 354.2 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 413.255 354.97 413.625 ;
      VIA 354.2 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 407.835 354.99 408.165 ;
      VIA 354.2 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 407.815 354.97 408.185 ;
      VIA 354.2 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 402.395 354.99 402.725 ;
      VIA 354.2 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 402.375 354.97 402.745 ;
      VIA 354.2 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 396.955 354.99 397.285 ;
      VIA 354.2 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 396.935 354.97 397.305 ;
      VIA 354.2 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 391.515 354.99 391.845 ;
      VIA 354.2 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 391.495 354.97 391.865 ;
      VIA 354.2 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 386.075 354.99 386.405 ;
      VIA 354.2 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 386.055 354.97 386.425 ;
      VIA 354.2 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 380.635 354.99 380.965 ;
      VIA 354.2 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 380.615 354.97 380.985 ;
      VIA 354.2 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 375.195 354.99 375.525 ;
      VIA 354.2 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 375.175 354.97 375.545 ;
      VIA 354.2 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 369.755 354.99 370.085 ;
      VIA 354.2 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 369.735 354.97 370.105 ;
      VIA 354.2 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 364.315 354.99 364.645 ;
      VIA 354.2 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 364.295 354.97 364.665 ;
      VIA 354.2 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 358.875 354.99 359.205 ;
      VIA 354.2 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 358.855 354.97 359.225 ;
      VIA 354.2 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 353.435 354.99 353.765 ;
      VIA 354.2 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 353.415 354.97 353.785 ;
      VIA 354.2 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 347.995 354.99 348.325 ;
      VIA 354.2 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 347.975 354.97 348.345 ;
      VIA 354.2 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 342.555 354.99 342.885 ;
      VIA 354.2 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 342.535 354.97 342.905 ;
      VIA 354.2 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 337.115 354.99 337.445 ;
      VIA 354.2 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 337.095 354.97 337.465 ;
      VIA 354.2 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 331.675 354.99 332.005 ;
      VIA 354.2 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 331.655 354.97 332.025 ;
      VIA 354.2 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 326.235 354.99 326.565 ;
      VIA 354.2 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 326.215 354.97 326.585 ;
      VIA 354.2 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 320.795 354.99 321.125 ;
      VIA 354.2 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 320.775 354.97 321.145 ;
      VIA 354.2 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 315.355 354.99 315.685 ;
      VIA 354.2 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 315.335 354.97 315.705 ;
      VIA 354.2 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 309.915 354.99 310.245 ;
      VIA 354.2 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 309.895 354.97 310.265 ;
      VIA 354.2 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 304.475 354.99 304.805 ;
      VIA 354.2 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 304.455 354.97 304.825 ;
      VIA 354.2 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 299.035 354.99 299.365 ;
      VIA 354.2 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 299.015 354.97 299.385 ;
      VIA 354.2 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 293.595 354.99 293.925 ;
      VIA 354.2 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 293.575 354.97 293.945 ;
      VIA 354.2 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 288.155 354.99 288.485 ;
      VIA 354.2 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 288.135 354.97 288.505 ;
      VIA 354.2 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 282.715 354.99 283.045 ;
      VIA 354.2 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 282.695 354.97 283.065 ;
      VIA 354.2 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 277.275 354.99 277.605 ;
      VIA 354.2 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 277.255 354.97 277.625 ;
      VIA 354.2 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 271.835 354.99 272.165 ;
      VIA 354.2 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 271.815 354.97 272.185 ;
      VIA 354.2 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 266.395 354.99 266.725 ;
      VIA 354.2 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 266.375 354.97 266.745 ;
      VIA 354.2 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 260.955 354.99 261.285 ;
      VIA 354.2 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 260.935 354.97 261.305 ;
      VIA 354.2 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 255.515 354.99 255.845 ;
      VIA 354.2 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 255.495 354.97 255.865 ;
      VIA 354.2 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 250.075 354.99 250.405 ;
      VIA 354.2 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 250.055 354.97 250.425 ;
      VIA 354.2 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 244.635 354.99 244.965 ;
      VIA 354.2 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 244.615 354.97 244.985 ;
      VIA 354.2 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 239.195 354.99 239.525 ;
      VIA 354.2 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 239.175 354.97 239.545 ;
      VIA 354.2 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 233.755 354.99 234.085 ;
      VIA 354.2 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 233.735 354.97 234.105 ;
      VIA 354.2 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 228.315 354.99 228.645 ;
      VIA 354.2 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 228.295 354.97 228.665 ;
      VIA 354.2 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 222.875 354.99 223.205 ;
      VIA 354.2 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 222.855 354.97 223.225 ;
      VIA 354.2 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 217.435 354.99 217.765 ;
      VIA 354.2 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 217.415 354.97 217.785 ;
      VIA 354.2 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 211.995 354.99 212.325 ;
      VIA 354.2 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 211.975 354.97 212.345 ;
      VIA 354.2 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 206.555 354.99 206.885 ;
      VIA 354.2 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 206.535 354.97 206.905 ;
      VIA 354.2 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 201.115 354.99 201.445 ;
      VIA 354.2 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 201.095 354.97 201.465 ;
      VIA 354.2 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 195.675 354.99 196.005 ;
      VIA 354.2 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 195.655 354.97 196.025 ;
      VIA 354.2 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 190.235 354.99 190.565 ;
      VIA 354.2 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 190.215 354.97 190.585 ;
      VIA 354.2 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 184.795 354.99 185.125 ;
      VIA 354.2 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 184.775 354.97 185.145 ;
      VIA 354.2 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 179.355 354.99 179.685 ;
      VIA 354.2 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 179.335 354.97 179.705 ;
      VIA 354.2 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 173.915 354.99 174.245 ;
      VIA 354.2 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 173.895 354.97 174.265 ;
      VIA 354.2 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 168.475 354.99 168.805 ;
      VIA 354.2 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 168.455 354.97 168.825 ;
      VIA 354.2 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 163.035 354.99 163.365 ;
      VIA 354.2 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 163.015 354.97 163.385 ;
      VIA 354.2 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 157.595 354.99 157.925 ;
      VIA 354.2 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 157.575 354.97 157.945 ;
      VIA 354.2 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 152.155 354.99 152.485 ;
      VIA 354.2 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 152.135 354.97 152.505 ;
      VIA 354.2 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 146.715 354.99 147.045 ;
      VIA 354.2 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 146.695 354.97 147.065 ;
      VIA 354.2 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 141.275 354.99 141.605 ;
      VIA 354.2 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 141.255 354.97 141.625 ;
      VIA 354.2 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 135.835 354.99 136.165 ;
      VIA 354.2 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 135.815 354.97 136.185 ;
      VIA 354.2 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 130.395 354.99 130.725 ;
      VIA 354.2 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 130.375 354.97 130.745 ;
      VIA 354.2 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 124.955 354.99 125.285 ;
      VIA 354.2 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 124.935 354.97 125.305 ;
      VIA 354.2 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 119.515 354.99 119.845 ;
      VIA 354.2 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 119.495 354.97 119.865 ;
      VIA 354.2 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 114.075 354.99 114.405 ;
      VIA 354.2 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 114.055 354.97 114.425 ;
      VIA 354.2 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 108.635 354.99 108.965 ;
      VIA 354.2 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 108.615 354.97 108.985 ;
      VIA 354.2 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 103.195 354.99 103.525 ;
      VIA 354.2 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 103.175 354.97 103.545 ;
      VIA 354.2 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 97.755 354.99 98.085 ;
      VIA 354.2 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 97.735 354.97 98.105 ;
      VIA 354.2 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 92.315 354.99 92.645 ;
      VIA 354.2 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 92.295 354.97 92.665 ;
      VIA 354.2 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 86.875 354.99 87.205 ;
      VIA 354.2 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 86.855 354.97 87.225 ;
      VIA 354.2 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 81.435 354.99 81.765 ;
      VIA 354.2 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 81.415 354.97 81.785 ;
      VIA 354.2 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 75.995 354.99 76.325 ;
      VIA 354.2 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 75.975 354.97 76.345 ;
      VIA 354.2 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 70.555 354.99 70.885 ;
      VIA 354.2 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 70.535 354.97 70.905 ;
      VIA 354.2 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 65.115 354.99 65.445 ;
      VIA 354.2 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 65.095 354.97 65.465 ;
      VIA 354.2 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 59.675 354.99 60.005 ;
      VIA 354.2 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 59.655 354.97 60.025 ;
      VIA 354.2 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 54.235 354.99 54.565 ;
      VIA 354.2 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 54.215 354.97 54.585 ;
      VIA 354.2 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 48.795 354.99 49.125 ;
      VIA 354.2 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 48.775 354.97 49.145 ;
      VIA 354.2 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 43.355 354.99 43.685 ;
      VIA 354.2 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 43.335 354.97 43.705 ;
      VIA 354.2 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 37.915 354.99 38.245 ;
      VIA 354.2 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 37.895 354.97 38.265 ;
      VIA 354.2 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 32.475 354.99 32.805 ;
      VIA 354.2 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 32.455 354.97 32.825 ;
      VIA 354.2 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 27.035 354.99 27.365 ;
      VIA 354.2 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 27.015 354.97 27.385 ;
      VIA 354.2 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 21.595 354.99 21.925 ;
      VIA 354.2 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 21.575 354.97 21.945 ;
      VIA 354.2 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 16.155 354.99 16.485 ;
      VIA 354.2 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 16.135 354.97 16.505 ;
      VIA 354.2 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 10.715 354.99 11.045 ;
      VIA 354.2 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 10.695 354.97 11.065 ;
      VIA 354.2 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  353.41 5.275 354.99 5.605 ;
      VIA 354.2 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  353.43 5.255 354.97 5.625 ;
      VIA 354.2 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 354.2 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 418.715 327.85 419.045 ;
      VIA 327.06 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 418.695 327.83 419.065 ;
      VIA 327.06 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 413.275 327.85 413.605 ;
      VIA 327.06 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 413.255 327.83 413.625 ;
      VIA 327.06 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 407.835 327.85 408.165 ;
      VIA 327.06 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 407.815 327.83 408.185 ;
      VIA 327.06 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 402.395 327.85 402.725 ;
      VIA 327.06 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 402.375 327.83 402.745 ;
      VIA 327.06 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 396.955 327.85 397.285 ;
      VIA 327.06 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 396.935 327.83 397.305 ;
      VIA 327.06 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 391.515 327.85 391.845 ;
      VIA 327.06 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 391.495 327.83 391.865 ;
      VIA 327.06 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 386.075 327.85 386.405 ;
      VIA 327.06 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 386.055 327.83 386.425 ;
      VIA 327.06 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 380.635 327.85 380.965 ;
      VIA 327.06 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 380.615 327.83 380.985 ;
      VIA 327.06 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 375.195 327.85 375.525 ;
      VIA 327.06 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 375.175 327.83 375.545 ;
      VIA 327.06 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 369.755 327.85 370.085 ;
      VIA 327.06 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 369.735 327.83 370.105 ;
      VIA 327.06 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 364.315 327.85 364.645 ;
      VIA 327.06 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 364.295 327.83 364.665 ;
      VIA 327.06 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 358.875 327.85 359.205 ;
      VIA 327.06 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 358.855 327.83 359.225 ;
      VIA 327.06 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 353.435 327.85 353.765 ;
      VIA 327.06 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 353.415 327.83 353.785 ;
      VIA 327.06 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 347.995 327.85 348.325 ;
      VIA 327.06 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 347.975 327.83 348.345 ;
      VIA 327.06 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 342.555 327.85 342.885 ;
      VIA 327.06 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 342.535 327.83 342.905 ;
      VIA 327.06 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 337.115 327.85 337.445 ;
      VIA 327.06 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 337.095 327.83 337.465 ;
      VIA 327.06 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 331.675 327.85 332.005 ;
      VIA 327.06 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 331.655 327.83 332.025 ;
      VIA 327.06 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 326.235 327.85 326.565 ;
      VIA 327.06 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 326.215 327.83 326.585 ;
      VIA 327.06 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 320.795 327.85 321.125 ;
      VIA 327.06 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 320.775 327.83 321.145 ;
      VIA 327.06 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 315.355 327.85 315.685 ;
      VIA 327.06 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 315.335 327.83 315.705 ;
      VIA 327.06 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 309.915 327.85 310.245 ;
      VIA 327.06 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 309.895 327.83 310.265 ;
      VIA 327.06 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 304.475 327.85 304.805 ;
      VIA 327.06 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 304.455 327.83 304.825 ;
      VIA 327.06 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 299.035 327.85 299.365 ;
      VIA 327.06 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 299.015 327.83 299.385 ;
      VIA 327.06 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 293.595 327.85 293.925 ;
      VIA 327.06 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 293.575 327.83 293.945 ;
      VIA 327.06 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 288.155 327.85 288.485 ;
      VIA 327.06 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 288.135 327.83 288.505 ;
      VIA 327.06 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 282.715 327.85 283.045 ;
      VIA 327.06 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 282.695 327.83 283.065 ;
      VIA 327.06 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 277.275 327.85 277.605 ;
      VIA 327.06 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 277.255 327.83 277.625 ;
      VIA 327.06 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 271.835 327.85 272.165 ;
      VIA 327.06 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 271.815 327.83 272.185 ;
      VIA 327.06 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 266.395 327.85 266.725 ;
      VIA 327.06 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 266.375 327.83 266.745 ;
      VIA 327.06 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 260.955 327.85 261.285 ;
      VIA 327.06 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 260.935 327.83 261.305 ;
      VIA 327.06 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 255.515 327.85 255.845 ;
      VIA 327.06 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 255.495 327.83 255.865 ;
      VIA 327.06 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 250.075 327.85 250.405 ;
      VIA 327.06 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 250.055 327.83 250.425 ;
      VIA 327.06 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 244.635 327.85 244.965 ;
      VIA 327.06 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 244.615 327.83 244.985 ;
      VIA 327.06 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 239.195 327.85 239.525 ;
      VIA 327.06 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 239.175 327.83 239.545 ;
      VIA 327.06 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 233.755 327.85 234.085 ;
      VIA 327.06 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 233.735 327.83 234.105 ;
      VIA 327.06 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 228.315 327.85 228.645 ;
      VIA 327.06 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 228.295 327.83 228.665 ;
      VIA 327.06 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 222.875 327.85 223.205 ;
      VIA 327.06 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 222.855 327.83 223.225 ;
      VIA 327.06 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 217.435 327.85 217.765 ;
      VIA 327.06 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 217.415 327.83 217.785 ;
      VIA 327.06 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 211.995 327.85 212.325 ;
      VIA 327.06 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 211.975 327.83 212.345 ;
      VIA 327.06 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 206.555 327.85 206.885 ;
      VIA 327.06 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 206.535 327.83 206.905 ;
      VIA 327.06 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 201.115 327.85 201.445 ;
      VIA 327.06 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 201.095 327.83 201.465 ;
      VIA 327.06 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 195.675 327.85 196.005 ;
      VIA 327.06 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 195.655 327.83 196.025 ;
      VIA 327.06 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 190.235 327.85 190.565 ;
      VIA 327.06 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 190.215 327.83 190.585 ;
      VIA 327.06 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 184.795 327.85 185.125 ;
      VIA 327.06 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 184.775 327.83 185.145 ;
      VIA 327.06 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 179.355 327.85 179.685 ;
      VIA 327.06 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 179.335 327.83 179.705 ;
      VIA 327.06 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 173.915 327.85 174.245 ;
      VIA 327.06 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 173.895 327.83 174.265 ;
      VIA 327.06 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 168.475 327.85 168.805 ;
      VIA 327.06 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 168.455 327.83 168.825 ;
      VIA 327.06 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 163.035 327.85 163.365 ;
      VIA 327.06 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 163.015 327.83 163.385 ;
      VIA 327.06 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 157.595 327.85 157.925 ;
      VIA 327.06 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 157.575 327.83 157.945 ;
      VIA 327.06 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 152.155 327.85 152.485 ;
      VIA 327.06 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 152.135 327.83 152.505 ;
      VIA 327.06 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 146.715 327.85 147.045 ;
      VIA 327.06 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 146.695 327.83 147.065 ;
      VIA 327.06 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 141.275 327.85 141.605 ;
      VIA 327.06 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 141.255 327.83 141.625 ;
      VIA 327.06 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 135.835 327.85 136.165 ;
      VIA 327.06 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 135.815 327.83 136.185 ;
      VIA 327.06 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 130.395 327.85 130.725 ;
      VIA 327.06 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 130.375 327.83 130.745 ;
      VIA 327.06 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 124.955 327.85 125.285 ;
      VIA 327.06 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 124.935 327.83 125.305 ;
      VIA 327.06 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 119.515 327.85 119.845 ;
      VIA 327.06 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 119.495 327.83 119.865 ;
      VIA 327.06 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 114.075 327.85 114.405 ;
      VIA 327.06 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 114.055 327.83 114.425 ;
      VIA 327.06 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 108.635 327.85 108.965 ;
      VIA 327.06 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 108.615 327.83 108.985 ;
      VIA 327.06 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 103.195 327.85 103.525 ;
      VIA 327.06 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 103.175 327.83 103.545 ;
      VIA 327.06 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 97.755 327.85 98.085 ;
      VIA 327.06 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 97.735 327.83 98.105 ;
      VIA 327.06 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 92.315 327.85 92.645 ;
      VIA 327.06 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 92.295 327.83 92.665 ;
      VIA 327.06 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 86.875 327.85 87.205 ;
      VIA 327.06 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 86.855 327.83 87.225 ;
      VIA 327.06 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 81.435 327.85 81.765 ;
      VIA 327.06 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 81.415 327.83 81.785 ;
      VIA 327.06 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 75.995 327.85 76.325 ;
      VIA 327.06 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 75.975 327.83 76.345 ;
      VIA 327.06 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 70.555 327.85 70.885 ;
      VIA 327.06 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 70.535 327.83 70.905 ;
      VIA 327.06 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 65.115 327.85 65.445 ;
      VIA 327.06 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 65.095 327.83 65.465 ;
      VIA 327.06 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 59.675 327.85 60.005 ;
      VIA 327.06 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 59.655 327.83 60.025 ;
      VIA 327.06 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 54.235 327.85 54.565 ;
      VIA 327.06 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 54.215 327.83 54.585 ;
      VIA 327.06 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 48.795 327.85 49.125 ;
      VIA 327.06 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 48.775 327.83 49.145 ;
      VIA 327.06 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 43.355 327.85 43.685 ;
      VIA 327.06 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 43.335 327.83 43.705 ;
      VIA 327.06 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 37.915 327.85 38.245 ;
      VIA 327.06 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 37.895 327.83 38.265 ;
      VIA 327.06 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 32.475 327.85 32.805 ;
      VIA 327.06 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 32.455 327.83 32.825 ;
      VIA 327.06 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 27.035 327.85 27.365 ;
      VIA 327.06 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 27.015 327.83 27.385 ;
      VIA 327.06 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 21.595 327.85 21.925 ;
      VIA 327.06 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 21.575 327.83 21.945 ;
      VIA 327.06 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 16.155 327.85 16.485 ;
      VIA 327.06 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 16.135 327.83 16.505 ;
      VIA 327.06 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 10.715 327.85 11.045 ;
      VIA 327.06 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 10.695 327.83 11.065 ;
      VIA 327.06 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  326.27 5.275 327.85 5.605 ;
      VIA 327.06 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  326.29 5.255 327.83 5.625 ;
      VIA 327.06 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 327.06 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 418.715 300.71 419.045 ;
      VIA 299.92 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 418.695 300.69 419.065 ;
      VIA 299.92 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 413.275 300.71 413.605 ;
      VIA 299.92 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 413.255 300.69 413.625 ;
      VIA 299.92 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 407.835 300.71 408.165 ;
      VIA 299.92 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 407.815 300.69 408.185 ;
      VIA 299.92 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 402.395 300.71 402.725 ;
      VIA 299.92 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 402.375 300.69 402.745 ;
      VIA 299.92 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 396.955 300.71 397.285 ;
      VIA 299.92 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 396.935 300.69 397.305 ;
      VIA 299.92 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 391.515 300.71 391.845 ;
      VIA 299.92 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 391.495 300.69 391.865 ;
      VIA 299.92 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 386.075 300.71 386.405 ;
      VIA 299.92 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 386.055 300.69 386.425 ;
      VIA 299.92 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 380.635 300.71 380.965 ;
      VIA 299.92 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 380.615 300.69 380.985 ;
      VIA 299.92 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 375.195 300.71 375.525 ;
      VIA 299.92 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 375.175 300.69 375.545 ;
      VIA 299.92 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 369.755 300.71 370.085 ;
      VIA 299.92 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 369.735 300.69 370.105 ;
      VIA 299.92 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 364.315 300.71 364.645 ;
      VIA 299.92 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 364.295 300.69 364.665 ;
      VIA 299.92 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 358.875 300.71 359.205 ;
      VIA 299.92 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 358.855 300.69 359.225 ;
      VIA 299.92 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 353.435 300.71 353.765 ;
      VIA 299.92 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 353.415 300.69 353.785 ;
      VIA 299.92 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 347.995 300.71 348.325 ;
      VIA 299.92 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 347.975 300.69 348.345 ;
      VIA 299.92 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 342.555 300.71 342.885 ;
      VIA 299.92 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 342.535 300.69 342.905 ;
      VIA 299.92 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 337.115 300.71 337.445 ;
      VIA 299.92 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 337.095 300.69 337.465 ;
      VIA 299.92 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 331.675 300.71 332.005 ;
      VIA 299.92 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 331.655 300.69 332.025 ;
      VIA 299.92 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 326.235 300.71 326.565 ;
      VIA 299.92 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 326.215 300.69 326.585 ;
      VIA 299.92 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 320.795 300.71 321.125 ;
      VIA 299.92 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 320.775 300.69 321.145 ;
      VIA 299.92 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 315.355 300.71 315.685 ;
      VIA 299.92 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 315.335 300.69 315.705 ;
      VIA 299.92 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 309.915 300.71 310.245 ;
      VIA 299.92 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 309.895 300.69 310.265 ;
      VIA 299.92 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 304.475 300.71 304.805 ;
      VIA 299.92 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 304.455 300.69 304.825 ;
      VIA 299.92 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 299.035 300.71 299.365 ;
      VIA 299.92 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 299.015 300.69 299.385 ;
      VIA 299.92 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 293.595 300.71 293.925 ;
      VIA 299.92 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 293.575 300.69 293.945 ;
      VIA 299.92 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 288.155 300.71 288.485 ;
      VIA 299.92 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 288.135 300.69 288.505 ;
      VIA 299.92 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 282.715 300.71 283.045 ;
      VIA 299.92 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 282.695 300.69 283.065 ;
      VIA 299.92 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 277.275 300.71 277.605 ;
      VIA 299.92 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 277.255 300.69 277.625 ;
      VIA 299.92 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 271.835 300.71 272.165 ;
      VIA 299.92 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 271.815 300.69 272.185 ;
      VIA 299.92 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 266.395 300.71 266.725 ;
      VIA 299.92 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 266.375 300.69 266.745 ;
      VIA 299.92 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 260.955 300.71 261.285 ;
      VIA 299.92 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 260.935 300.69 261.305 ;
      VIA 299.92 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 255.515 300.71 255.845 ;
      VIA 299.92 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 255.495 300.69 255.865 ;
      VIA 299.92 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 250.075 300.71 250.405 ;
      VIA 299.92 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 250.055 300.69 250.425 ;
      VIA 299.92 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 244.635 300.71 244.965 ;
      VIA 299.92 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 244.615 300.69 244.985 ;
      VIA 299.92 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 239.195 300.71 239.525 ;
      VIA 299.92 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 239.175 300.69 239.545 ;
      VIA 299.92 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 233.755 300.71 234.085 ;
      VIA 299.92 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 233.735 300.69 234.105 ;
      VIA 299.92 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 228.315 300.71 228.645 ;
      VIA 299.92 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 228.295 300.69 228.665 ;
      VIA 299.92 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 222.875 300.71 223.205 ;
      VIA 299.92 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 222.855 300.69 223.225 ;
      VIA 299.92 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 217.435 300.71 217.765 ;
      VIA 299.92 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 217.415 300.69 217.785 ;
      VIA 299.92 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 211.995 300.71 212.325 ;
      VIA 299.92 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 211.975 300.69 212.345 ;
      VIA 299.92 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 206.555 300.71 206.885 ;
      VIA 299.92 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 206.535 300.69 206.905 ;
      VIA 299.92 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 201.115 300.71 201.445 ;
      VIA 299.92 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 201.095 300.69 201.465 ;
      VIA 299.92 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 195.675 300.71 196.005 ;
      VIA 299.92 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 195.655 300.69 196.025 ;
      VIA 299.92 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 190.235 300.71 190.565 ;
      VIA 299.92 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 190.215 300.69 190.585 ;
      VIA 299.92 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 184.795 300.71 185.125 ;
      VIA 299.92 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 184.775 300.69 185.145 ;
      VIA 299.92 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 179.355 300.71 179.685 ;
      VIA 299.92 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 179.335 300.69 179.705 ;
      VIA 299.92 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 173.915 300.71 174.245 ;
      VIA 299.92 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 173.895 300.69 174.265 ;
      VIA 299.92 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 168.475 300.71 168.805 ;
      VIA 299.92 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 168.455 300.69 168.825 ;
      VIA 299.92 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 163.035 300.71 163.365 ;
      VIA 299.92 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 163.015 300.69 163.385 ;
      VIA 299.92 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 157.595 300.71 157.925 ;
      VIA 299.92 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 157.575 300.69 157.945 ;
      VIA 299.92 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 152.155 300.71 152.485 ;
      VIA 299.92 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 152.135 300.69 152.505 ;
      VIA 299.92 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 146.715 300.71 147.045 ;
      VIA 299.92 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 146.695 300.69 147.065 ;
      VIA 299.92 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 141.275 300.71 141.605 ;
      VIA 299.92 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 141.255 300.69 141.625 ;
      VIA 299.92 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 135.835 300.71 136.165 ;
      VIA 299.92 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 135.815 300.69 136.185 ;
      VIA 299.92 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 130.395 300.71 130.725 ;
      VIA 299.92 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 130.375 300.69 130.745 ;
      VIA 299.92 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 124.955 300.71 125.285 ;
      VIA 299.92 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 124.935 300.69 125.305 ;
      VIA 299.92 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 119.515 300.71 119.845 ;
      VIA 299.92 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 119.495 300.69 119.865 ;
      VIA 299.92 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 114.075 300.71 114.405 ;
      VIA 299.92 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 114.055 300.69 114.425 ;
      VIA 299.92 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 108.635 300.71 108.965 ;
      VIA 299.92 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 108.615 300.69 108.985 ;
      VIA 299.92 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 103.195 300.71 103.525 ;
      VIA 299.92 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 103.175 300.69 103.545 ;
      VIA 299.92 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 97.755 300.71 98.085 ;
      VIA 299.92 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 97.735 300.69 98.105 ;
      VIA 299.92 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 92.315 300.71 92.645 ;
      VIA 299.92 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 92.295 300.69 92.665 ;
      VIA 299.92 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 86.875 300.71 87.205 ;
      VIA 299.92 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 86.855 300.69 87.225 ;
      VIA 299.92 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 81.435 300.71 81.765 ;
      VIA 299.92 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 81.415 300.69 81.785 ;
      VIA 299.92 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 75.995 300.71 76.325 ;
      VIA 299.92 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 75.975 300.69 76.345 ;
      VIA 299.92 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 70.555 300.71 70.885 ;
      VIA 299.92 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 70.535 300.69 70.905 ;
      VIA 299.92 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 65.115 300.71 65.445 ;
      VIA 299.92 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 65.095 300.69 65.465 ;
      VIA 299.92 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 59.675 300.71 60.005 ;
      VIA 299.92 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 59.655 300.69 60.025 ;
      VIA 299.92 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 54.235 300.71 54.565 ;
      VIA 299.92 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 54.215 300.69 54.585 ;
      VIA 299.92 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 48.795 300.71 49.125 ;
      VIA 299.92 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 48.775 300.69 49.145 ;
      VIA 299.92 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 43.355 300.71 43.685 ;
      VIA 299.92 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 43.335 300.69 43.705 ;
      VIA 299.92 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 37.915 300.71 38.245 ;
      VIA 299.92 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 37.895 300.69 38.265 ;
      VIA 299.92 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 32.475 300.71 32.805 ;
      VIA 299.92 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 32.455 300.69 32.825 ;
      VIA 299.92 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 27.035 300.71 27.365 ;
      VIA 299.92 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 27.015 300.69 27.385 ;
      VIA 299.92 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 21.595 300.71 21.925 ;
      VIA 299.92 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 21.575 300.69 21.945 ;
      VIA 299.92 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 16.155 300.71 16.485 ;
      VIA 299.92 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 16.135 300.69 16.505 ;
      VIA 299.92 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 10.715 300.71 11.045 ;
      VIA 299.92 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 10.695 300.69 11.065 ;
      VIA 299.92 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  299.13 5.275 300.71 5.605 ;
      VIA 299.92 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  299.15 5.255 300.69 5.625 ;
      VIA 299.92 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 299.92 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 418.715 273.57 419.045 ;
      VIA 272.78 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 418.695 273.55 419.065 ;
      VIA 272.78 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 413.275 273.57 413.605 ;
      VIA 272.78 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 413.255 273.55 413.625 ;
      VIA 272.78 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 407.835 273.57 408.165 ;
      VIA 272.78 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 407.815 273.55 408.185 ;
      VIA 272.78 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 402.395 273.57 402.725 ;
      VIA 272.78 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 402.375 273.55 402.745 ;
      VIA 272.78 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 396.955 273.57 397.285 ;
      VIA 272.78 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 396.935 273.55 397.305 ;
      VIA 272.78 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 391.515 273.57 391.845 ;
      VIA 272.78 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 391.495 273.55 391.865 ;
      VIA 272.78 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 386.075 273.57 386.405 ;
      VIA 272.78 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 386.055 273.55 386.425 ;
      VIA 272.78 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 380.635 273.57 380.965 ;
      VIA 272.78 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 380.615 273.55 380.985 ;
      VIA 272.78 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 375.195 273.57 375.525 ;
      VIA 272.78 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 375.175 273.55 375.545 ;
      VIA 272.78 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 369.755 273.57 370.085 ;
      VIA 272.78 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 369.735 273.55 370.105 ;
      VIA 272.78 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 364.315 273.57 364.645 ;
      VIA 272.78 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 364.295 273.55 364.665 ;
      VIA 272.78 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 358.875 273.57 359.205 ;
      VIA 272.78 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 358.855 273.55 359.225 ;
      VIA 272.78 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 353.435 273.57 353.765 ;
      VIA 272.78 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 353.415 273.55 353.785 ;
      VIA 272.78 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 347.995 273.57 348.325 ;
      VIA 272.78 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 347.975 273.55 348.345 ;
      VIA 272.78 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 342.555 273.57 342.885 ;
      VIA 272.78 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 342.535 273.55 342.905 ;
      VIA 272.78 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 337.115 273.57 337.445 ;
      VIA 272.78 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 337.095 273.55 337.465 ;
      VIA 272.78 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 331.675 273.57 332.005 ;
      VIA 272.78 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 331.655 273.55 332.025 ;
      VIA 272.78 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 326.235 273.57 326.565 ;
      VIA 272.78 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 326.215 273.55 326.585 ;
      VIA 272.78 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 320.795 273.57 321.125 ;
      VIA 272.78 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 320.775 273.55 321.145 ;
      VIA 272.78 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 315.355 273.57 315.685 ;
      VIA 272.78 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 315.335 273.55 315.705 ;
      VIA 272.78 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 309.915 273.57 310.245 ;
      VIA 272.78 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 309.895 273.55 310.265 ;
      VIA 272.78 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 304.475 273.57 304.805 ;
      VIA 272.78 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 304.455 273.55 304.825 ;
      VIA 272.78 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 299.035 273.57 299.365 ;
      VIA 272.78 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 299.015 273.55 299.385 ;
      VIA 272.78 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 293.595 273.57 293.925 ;
      VIA 272.78 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 293.575 273.55 293.945 ;
      VIA 272.78 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 288.155 273.57 288.485 ;
      VIA 272.78 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 288.135 273.55 288.505 ;
      VIA 272.78 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 282.715 273.57 283.045 ;
      VIA 272.78 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 282.695 273.55 283.065 ;
      VIA 272.78 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 277.275 273.57 277.605 ;
      VIA 272.78 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 277.255 273.55 277.625 ;
      VIA 272.78 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 271.835 273.57 272.165 ;
      VIA 272.78 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 271.815 273.55 272.185 ;
      VIA 272.78 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 266.395 273.57 266.725 ;
      VIA 272.78 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 266.375 273.55 266.745 ;
      VIA 272.78 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 260.955 273.57 261.285 ;
      VIA 272.78 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 260.935 273.55 261.305 ;
      VIA 272.78 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 255.515 273.57 255.845 ;
      VIA 272.78 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 255.495 273.55 255.865 ;
      VIA 272.78 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 250.075 273.57 250.405 ;
      VIA 272.78 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 250.055 273.55 250.425 ;
      VIA 272.78 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 244.635 273.57 244.965 ;
      VIA 272.78 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 244.615 273.55 244.985 ;
      VIA 272.78 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 239.195 273.57 239.525 ;
      VIA 272.78 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 239.175 273.55 239.545 ;
      VIA 272.78 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 233.755 273.57 234.085 ;
      VIA 272.78 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 233.735 273.55 234.105 ;
      VIA 272.78 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 228.315 273.57 228.645 ;
      VIA 272.78 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 228.295 273.55 228.665 ;
      VIA 272.78 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 222.875 273.57 223.205 ;
      VIA 272.78 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 222.855 273.55 223.225 ;
      VIA 272.78 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 217.435 273.57 217.765 ;
      VIA 272.78 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 217.415 273.55 217.785 ;
      VIA 272.78 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 211.995 273.57 212.325 ;
      VIA 272.78 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 211.975 273.55 212.345 ;
      VIA 272.78 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 206.555 273.57 206.885 ;
      VIA 272.78 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 206.535 273.55 206.905 ;
      VIA 272.78 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 201.115 273.57 201.445 ;
      VIA 272.78 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 201.095 273.55 201.465 ;
      VIA 272.78 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 195.675 273.57 196.005 ;
      VIA 272.78 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 195.655 273.55 196.025 ;
      VIA 272.78 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 190.235 273.57 190.565 ;
      VIA 272.78 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 190.215 273.55 190.585 ;
      VIA 272.78 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 184.795 273.57 185.125 ;
      VIA 272.78 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 184.775 273.55 185.145 ;
      VIA 272.78 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 179.355 273.57 179.685 ;
      VIA 272.78 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 179.335 273.55 179.705 ;
      VIA 272.78 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 173.915 273.57 174.245 ;
      VIA 272.78 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 173.895 273.55 174.265 ;
      VIA 272.78 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 168.475 273.57 168.805 ;
      VIA 272.78 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 168.455 273.55 168.825 ;
      VIA 272.78 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 163.035 273.57 163.365 ;
      VIA 272.78 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 163.015 273.55 163.385 ;
      VIA 272.78 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 157.595 273.57 157.925 ;
      VIA 272.78 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 157.575 273.55 157.945 ;
      VIA 272.78 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 152.155 273.57 152.485 ;
      VIA 272.78 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 152.135 273.55 152.505 ;
      VIA 272.78 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 146.715 273.57 147.045 ;
      VIA 272.78 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 146.695 273.55 147.065 ;
      VIA 272.78 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 141.275 273.57 141.605 ;
      VIA 272.78 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 141.255 273.55 141.625 ;
      VIA 272.78 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 135.835 273.57 136.165 ;
      VIA 272.78 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 135.815 273.55 136.185 ;
      VIA 272.78 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 130.395 273.57 130.725 ;
      VIA 272.78 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 130.375 273.55 130.745 ;
      VIA 272.78 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 124.955 273.57 125.285 ;
      VIA 272.78 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 124.935 273.55 125.305 ;
      VIA 272.78 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 119.515 273.57 119.845 ;
      VIA 272.78 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 119.495 273.55 119.865 ;
      VIA 272.78 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 114.075 273.57 114.405 ;
      VIA 272.78 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 114.055 273.55 114.425 ;
      VIA 272.78 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 108.635 273.57 108.965 ;
      VIA 272.78 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 108.615 273.55 108.985 ;
      VIA 272.78 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 103.195 273.57 103.525 ;
      VIA 272.78 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 103.175 273.55 103.545 ;
      VIA 272.78 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 97.755 273.57 98.085 ;
      VIA 272.78 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 97.735 273.55 98.105 ;
      VIA 272.78 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 92.315 273.57 92.645 ;
      VIA 272.78 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 92.295 273.55 92.665 ;
      VIA 272.78 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 86.875 273.57 87.205 ;
      VIA 272.78 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 86.855 273.55 87.225 ;
      VIA 272.78 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 81.435 273.57 81.765 ;
      VIA 272.78 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 81.415 273.55 81.785 ;
      VIA 272.78 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 75.995 273.57 76.325 ;
      VIA 272.78 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 75.975 273.55 76.345 ;
      VIA 272.78 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 70.555 273.57 70.885 ;
      VIA 272.78 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 70.535 273.55 70.905 ;
      VIA 272.78 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 65.115 273.57 65.445 ;
      VIA 272.78 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 65.095 273.55 65.465 ;
      VIA 272.78 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 59.675 273.57 60.005 ;
      VIA 272.78 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 59.655 273.55 60.025 ;
      VIA 272.78 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 54.235 273.57 54.565 ;
      VIA 272.78 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 54.215 273.55 54.585 ;
      VIA 272.78 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 48.795 273.57 49.125 ;
      VIA 272.78 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 48.775 273.55 49.145 ;
      VIA 272.78 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 43.355 273.57 43.685 ;
      VIA 272.78 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 43.335 273.55 43.705 ;
      VIA 272.78 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 37.915 273.57 38.245 ;
      VIA 272.78 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 37.895 273.55 38.265 ;
      VIA 272.78 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 32.475 273.57 32.805 ;
      VIA 272.78 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 32.455 273.55 32.825 ;
      VIA 272.78 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 27.035 273.57 27.365 ;
      VIA 272.78 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 27.015 273.55 27.385 ;
      VIA 272.78 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 21.595 273.57 21.925 ;
      VIA 272.78 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 21.575 273.55 21.945 ;
      VIA 272.78 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 16.155 273.57 16.485 ;
      VIA 272.78 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 16.135 273.55 16.505 ;
      VIA 272.78 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 10.715 273.57 11.045 ;
      VIA 272.78 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 10.695 273.55 11.065 ;
      VIA 272.78 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 5.275 273.57 5.605 ;
      VIA 272.78 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 5.255 273.55 5.625 ;
      VIA 272.78 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 418.715 246.43 419.045 ;
      VIA 245.64 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 418.695 246.41 419.065 ;
      VIA 245.64 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 413.275 246.43 413.605 ;
      VIA 245.64 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 413.255 246.41 413.625 ;
      VIA 245.64 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 407.835 246.43 408.165 ;
      VIA 245.64 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 407.815 246.41 408.185 ;
      VIA 245.64 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 402.395 246.43 402.725 ;
      VIA 245.64 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 402.375 246.41 402.745 ;
      VIA 245.64 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 396.955 246.43 397.285 ;
      VIA 245.64 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 396.935 246.41 397.305 ;
      VIA 245.64 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 391.515 246.43 391.845 ;
      VIA 245.64 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 391.495 246.41 391.865 ;
      VIA 245.64 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 386.075 246.43 386.405 ;
      VIA 245.64 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 386.055 246.41 386.425 ;
      VIA 245.64 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 380.635 246.43 380.965 ;
      VIA 245.64 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 380.615 246.41 380.985 ;
      VIA 245.64 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 375.195 246.43 375.525 ;
      VIA 245.64 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 375.175 246.41 375.545 ;
      VIA 245.64 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 369.755 246.43 370.085 ;
      VIA 245.64 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 369.735 246.41 370.105 ;
      VIA 245.64 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 364.315 246.43 364.645 ;
      VIA 245.64 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 364.295 246.41 364.665 ;
      VIA 245.64 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 358.875 246.43 359.205 ;
      VIA 245.64 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 358.855 246.41 359.225 ;
      VIA 245.64 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 353.435 246.43 353.765 ;
      VIA 245.64 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 353.415 246.41 353.785 ;
      VIA 245.64 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 347.995 246.43 348.325 ;
      VIA 245.64 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 347.975 246.41 348.345 ;
      VIA 245.64 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 342.555 246.43 342.885 ;
      VIA 245.64 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 342.535 246.41 342.905 ;
      VIA 245.64 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 337.115 246.43 337.445 ;
      VIA 245.64 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 337.095 246.41 337.465 ;
      VIA 245.64 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 331.675 246.43 332.005 ;
      VIA 245.64 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 331.655 246.41 332.025 ;
      VIA 245.64 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 326.235 246.43 326.565 ;
      VIA 245.64 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 326.215 246.41 326.585 ;
      VIA 245.64 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 320.795 246.43 321.125 ;
      VIA 245.64 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 320.775 246.41 321.145 ;
      VIA 245.64 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 315.355 246.43 315.685 ;
      VIA 245.64 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 315.335 246.41 315.705 ;
      VIA 245.64 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 309.915 246.43 310.245 ;
      VIA 245.64 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 309.895 246.41 310.265 ;
      VIA 245.64 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 304.475 246.43 304.805 ;
      VIA 245.64 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 304.455 246.41 304.825 ;
      VIA 245.64 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 299.035 246.43 299.365 ;
      VIA 245.64 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 299.015 246.41 299.385 ;
      VIA 245.64 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 293.595 246.43 293.925 ;
      VIA 245.64 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 293.575 246.41 293.945 ;
      VIA 245.64 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 288.155 246.43 288.485 ;
      VIA 245.64 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 288.135 246.41 288.505 ;
      VIA 245.64 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 282.715 246.43 283.045 ;
      VIA 245.64 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 282.695 246.41 283.065 ;
      VIA 245.64 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 277.275 246.43 277.605 ;
      VIA 245.64 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 277.255 246.41 277.625 ;
      VIA 245.64 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 271.835 246.43 272.165 ;
      VIA 245.64 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 271.815 246.41 272.185 ;
      VIA 245.64 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 266.395 246.43 266.725 ;
      VIA 245.64 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 266.375 246.41 266.745 ;
      VIA 245.64 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 260.955 246.43 261.285 ;
      VIA 245.64 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 260.935 246.41 261.305 ;
      VIA 245.64 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 255.515 246.43 255.845 ;
      VIA 245.64 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 255.495 246.41 255.865 ;
      VIA 245.64 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 250.075 246.43 250.405 ;
      VIA 245.64 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 250.055 246.41 250.425 ;
      VIA 245.64 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 244.635 246.43 244.965 ;
      VIA 245.64 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 244.615 246.41 244.985 ;
      VIA 245.64 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 239.195 246.43 239.525 ;
      VIA 245.64 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 239.175 246.41 239.545 ;
      VIA 245.64 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 233.755 246.43 234.085 ;
      VIA 245.64 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 233.735 246.41 234.105 ;
      VIA 245.64 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 228.315 246.43 228.645 ;
      VIA 245.64 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 228.295 246.41 228.665 ;
      VIA 245.64 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 222.875 246.43 223.205 ;
      VIA 245.64 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 222.855 246.41 223.225 ;
      VIA 245.64 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 217.435 246.43 217.765 ;
      VIA 245.64 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 217.415 246.41 217.785 ;
      VIA 245.64 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 211.995 246.43 212.325 ;
      VIA 245.64 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 211.975 246.41 212.345 ;
      VIA 245.64 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 206.555 246.43 206.885 ;
      VIA 245.64 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 206.535 246.41 206.905 ;
      VIA 245.64 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 201.115 246.43 201.445 ;
      VIA 245.64 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 201.095 246.41 201.465 ;
      VIA 245.64 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 195.675 246.43 196.005 ;
      VIA 245.64 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 195.655 246.41 196.025 ;
      VIA 245.64 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 190.235 246.43 190.565 ;
      VIA 245.64 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 190.215 246.41 190.585 ;
      VIA 245.64 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 184.795 246.43 185.125 ;
      VIA 245.64 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 184.775 246.41 185.145 ;
      VIA 245.64 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 179.355 246.43 179.685 ;
      VIA 245.64 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 179.335 246.41 179.705 ;
      VIA 245.64 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 173.915 246.43 174.245 ;
      VIA 245.64 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 173.895 246.41 174.265 ;
      VIA 245.64 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 168.475 246.43 168.805 ;
      VIA 245.64 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 168.455 246.41 168.825 ;
      VIA 245.64 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 163.035 246.43 163.365 ;
      VIA 245.64 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 163.015 246.41 163.385 ;
      VIA 245.64 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 157.595 246.43 157.925 ;
      VIA 245.64 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 157.575 246.41 157.945 ;
      VIA 245.64 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 152.155 246.43 152.485 ;
      VIA 245.64 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 152.135 246.41 152.505 ;
      VIA 245.64 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 146.715 246.43 147.045 ;
      VIA 245.64 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 146.695 246.41 147.065 ;
      VIA 245.64 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 141.275 246.43 141.605 ;
      VIA 245.64 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 141.255 246.41 141.625 ;
      VIA 245.64 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 135.835 246.43 136.165 ;
      VIA 245.64 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 135.815 246.41 136.185 ;
      VIA 245.64 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 130.395 246.43 130.725 ;
      VIA 245.64 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 130.375 246.41 130.745 ;
      VIA 245.64 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 124.955 246.43 125.285 ;
      VIA 245.64 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 124.935 246.41 125.305 ;
      VIA 245.64 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 119.515 246.43 119.845 ;
      VIA 245.64 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 119.495 246.41 119.865 ;
      VIA 245.64 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 114.075 246.43 114.405 ;
      VIA 245.64 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 114.055 246.41 114.425 ;
      VIA 245.64 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 108.635 246.43 108.965 ;
      VIA 245.64 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 108.615 246.41 108.985 ;
      VIA 245.64 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 103.195 246.43 103.525 ;
      VIA 245.64 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 103.175 246.41 103.545 ;
      VIA 245.64 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 97.755 246.43 98.085 ;
      VIA 245.64 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 97.735 246.41 98.105 ;
      VIA 245.64 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 92.315 246.43 92.645 ;
      VIA 245.64 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 92.295 246.41 92.665 ;
      VIA 245.64 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 86.875 246.43 87.205 ;
      VIA 245.64 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 86.855 246.41 87.225 ;
      VIA 245.64 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 81.435 246.43 81.765 ;
      VIA 245.64 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 81.415 246.41 81.785 ;
      VIA 245.64 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 75.995 246.43 76.325 ;
      VIA 245.64 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 75.975 246.41 76.345 ;
      VIA 245.64 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 70.555 246.43 70.885 ;
      VIA 245.64 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 70.535 246.41 70.905 ;
      VIA 245.64 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 65.115 246.43 65.445 ;
      VIA 245.64 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 65.095 246.41 65.465 ;
      VIA 245.64 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 59.675 246.43 60.005 ;
      VIA 245.64 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 59.655 246.41 60.025 ;
      VIA 245.64 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 54.235 246.43 54.565 ;
      VIA 245.64 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 54.215 246.41 54.585 ;
      VIA 245.64 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 48.795 246.43 49.125 ;
      VIA 245.64 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 48.775 246.41 49.145 ;
      VIA 245.64 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 43.355 246.43 43.685 ;
      VIA 245.64 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 43.335 246.41 43.705 ;
      VIA 245.64 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 37.915 246.43 38.245 ;
      VIA 245.64 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 37.895 246.41 38.265 ;
      VIA 245.64 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 32.475 246.43 32.805 ;
      VIA 245.64 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 32.455 246.41 32.825 ;
      VIA 245.64 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 27.035 246.43 27.365 ;
      VIA 245.64 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 27.015 246.41 27.385 ;
      VIA 245.64 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 21.595 246.43 21.925 ;
      VIA 245.64 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 21.575 246.41 21.945 ;
      VIA 245.64 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 16.155 246.43 16.485 ;
      VIA 245.64 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 16.135 246.41 16.505 ;
      VIA 245.64 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 10.715 246.43 11.045 ;
      VIA 245.64 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 10.695 246.41 11.065 ;
      VIA 245.64 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 5.275 246.43 5.605 ;
      VIA 245.64 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 5.255 246.41 5.625 ;
      VIA 245.64 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 418.715 219.29 419.045 ;
      VIA 218.5 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 418.695 219.27 419.065 ;
      VIA 218.5 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 413.275 219.29 413.605 ;
      VIA 218.5 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 413.255 219.27 413.625 ;
      VIA 218.5 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 407.835 219.29 408.165 ;
      VIA 218.5 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 407.815 219.27 408.185 ;
      VIA 218.5 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 402.395 219.29 402.725 ;
      VIA 218.5 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 402.375 219.27 402.745 ;
      VIA 218.5 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 396.955 219.29 397.285 ;
      VIA 218.5 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 396.935 219.27 397.305 ;
      VIA 218.5 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 391.515 219.29 391.845 ;
      VIA 218.5 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 391.495 219.27 391.865 ;
      VIA 218.5 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 386.075 219.29 386.405 ;
      VIA 218.5 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 386.055 219.27 386.425 ;
      VIA 218.5 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 380.635 219.29 380.965 ;
      VIA 218.5 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 380.615 219.27 380.985 ;
      VIA 218.5 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 375.195 219.29 375.525 ;
      VIA 218.5 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 375.175 219.27 375.545 ;
      VIA 218.5 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 369.755 219.29 370.085 ;
      VIA 218.5 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 369.735 219.27 370.105 ;
      VIA 218.5 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 364.315 219.29 364.645 ;
      VIA 218.5 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 364.295 219.27 364.665 ;
      VIA 218.5 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 358.875 219.29 359.205 ;
      VIA 218.5 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 358.855 219.27 359.225 ;
      VIA 218.5 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 353.435 219.29 353.765 ;
      VIA 218.5 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 353.415 219.27 353.785 ;
      VIA 218.5 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 347.995 219.29 348.325 ;
      VIA 218.5 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 347.975 219.27 348.345 ;
      VIA 218.5 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 342.555 219.29 342.885 ;
      VIA 218.5 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 342.535 219.27 342.905 ;
      VIA 218.5 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 337.115 219.29 337.445 ;
      VIA 218.5 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 337.095 219.27 337.465 ;
      VIA 218.5 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 331.675 219.29 332.005 ;
      VIA 218.5 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 331.655 219.27 332.025 ;
      VIA 218.5 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 326.235 219.29 326.565 ;
      VIA 218.5 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 326.215 219.27 326.585 ;
      VIA 218.5 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 320.795 219.29 321.125 ;
      VIA 218.5 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 320.775 219.27 321.145 ;
      VIA 218.5 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 315.355 219.29 315.685 ;
      VIA 218.5 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 315.335 219.27 315.705 ;
      VIA 218.5 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 309.915 219.29 310.245 ;
      VIA 218.5 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 309.895 219.27 310.265 ;
      VIA 218.5 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 304.475 219.29 304.805 ;
      VIA 218.5 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 304.455 219.27 304.825 ;
      VIA 218.5 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 299.035 219.29 299.365 ;
      VIA 218.5 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 299.015 219.27 299.385 ;
      VIA 218.5 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 293.595 219.29 293.925 ;
      VIA 218.5 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 293.575 219.27 293.945 ;
      VIA 218.5 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 288.155 219.29 288.485 ;
      VIA 218.5 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 288.135 219.27 288.505 ;
      VIA 218.5 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 282.715 219.29 283.045 ;
      VIA 218.5 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 282.695 219.27 283.065 ;
      VIA 218.5 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 277.275 219.29 277.605 ;
      VIA 218.5 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 277.255 219.27 277.625 ;
      VIA 218.5 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 271.835 219.29 272.165 ;
      VIA 218.5 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 271.815 219.27 272.185 ;
      VIA 218.5 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 266.395 219.29 266.725 ;
      VIA 218.5 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 266.375 219.27 266.745 ;
      VIA 218.5 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 260.955 219.29 261.285 ;
      VIA 218.5 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 260.935 219.27 261.305 ;
      VIA 218.5 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 255.515 219.29 255.845 ;
      VIA 218.5 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 255.495 219.27 255.865 ;
      VIA 218.5 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 250.075 219.29 250.405 ;
      VIA 218.5 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 250.055 219.27 250.425 ;
      VIA 218.5 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 244.635 219.29 244.965 ;
      VIA 218.5 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 244.615 219.27 244.985 ;
      VIA 218.5 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 239.195 219.29 239.525 ;
      VIA 218.5 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 239.175 219.27 239.545 ;
      VIA 218.5 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 233.755 219.29 234.085 ;
      VIA 218.5 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 233.735 219.27 234.105 ;
      VIA 218.5 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 228.315 219.29 228.645 ;
      VIA 218.5 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 228.295 219.27 228.665 ;
      VIA 218.5 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 222.875 219.29 223.205 ;
      VIA 218.5 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 222.855 219.27 223.225 ;
      VIA 218.5 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 217.435 219.29 217.765 ;
      VIA 218.5 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 217.415 219.27 217.785 ;
      VIA 218.5 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 211.995 219.29 212.325 ;
      VIA 218.5 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 211.975 219.27 212.345 ;
      VIA 218.5 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 206.555 219.29 206.885 ;
      VIA 218.5 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 206.535 219.27 206.905 ;
      VIA 218.5 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 201.115 219.29 201.445 ;
      VIA 218.5 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 201.095 219.27 201.465 ;
      VIA 218.5 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 195.675 219.29 196.005 ;
      VIA 218.5 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 195.655 219.27 196.025 ;
      VIA 218.5 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 190.235 219.29 190.565 ;
      VIA 218.5 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 190.215 219.27 190.585 ;
      VIA 218.5 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 184.795 219.29 185.125 ;
      VIA 218.5 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 184.775 219.27 185.145 ;
      VIA 218.5 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 179.355 219.29 179.685 ;
      VIA 218.5 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 179.335 219.27 179.705 ;
      VIA 218.5 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 173.915 219.29 174.245 ;
      VIA 218.5 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 173.895 219.27 174.265 ;
      VIA 218.5 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 168.475 219.29 168.805 ;
      VIA 218.5 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 168.455 219.27 168.825 ;
      VIA 218.5 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 163.035 219.29 163.365 ;
      VIA 218.5 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 163.015 219.27 163.385 ;
      VIA 218.5 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 157.595 219.29 157.925 ;
      VIA 218.5 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 157.575 219.27 157.945 ;
      VIA 218.5 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 152.155 219.29 152.485 ;
      VIA 218.5 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 152.135 219.27 152.505 ;
      VIA 218.5 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 146.715 219.29 147.045 ;
      VIA 218.5 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 146.695 219.27 147.065 ;
      VIA 218.5 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 141.275 219.29 141.605 ;
      VIA 218.5 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 141.255 219.27 141.625 ;
      VIA 218.5 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 135.835 219.29 136.165 ;
      VIA 218.5 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 135.815 219.27 136.185 ;
      VIA 218.5 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 130.395 219.29 130.725 ;
      VIA 218.5 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 130.375 219.27 130.745 ;
      VIA 218.5 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 124.955 219.29 125.285 ;
      VIA 218.5 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 124.935 219.27 125.305 ;
      VIA 218.5 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 119.515 219.29 119.845 ;
      VIA 218.5 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 119.495 219.27 119.865 ;
      VIA 218.5 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 114.075 219.29 114.405 ;
      VIA 218.5 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 114.055 219.27 114.425 ;
      VIA 218.5 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 108.635 219.29 108.965 ;
      VIA 218.5 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 108.615 219.27 108.985 ;
      VIA 218.5 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 103.195 219.29 103.525 ;
      VIA 218.5 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 103.175 219.27 103.545 ;
      VIA 218.5 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 97.755 219.29 98.085 ;
      VIA 218.5 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 97.735 219.27 98.105 ;
      VIA 218.5 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 92.315 219.29 92.645 ;
      VIA 218.5 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 92.295 219.27 92.665 ;
      VIA 218.5 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 86.875 219.29 87.205 ;
      VIA 218.5 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 86.855 219.27 87.225 ;
      VIA 218.5 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 81.435 219.29 81.765 ;
      VIA 218.5 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 81.415 219.27 81.785 ;
      VIA 218.5 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 75.995 219.29 76.325 ;
      VIA 218.5 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 75.975 219.27 76.345 ;
      VIA 218.5 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 70.555 219.29 70.885 ;
      VIA 218.5 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 70.535 219.27 70.905 ;
      VIA 218.5 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 65.115 219.29 65.445 ;
      VIA 218.5 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 65.095 219.27 65.465 ;
      VIA 218.5 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 59.675 219.29 60.005 ;
      VIA 218.5 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 59.655 219.27 60.025 ;
      VIA 218.5 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 54.235 219.29 54.565 ;
      VIA 218.5 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 54.215 219.27 54.585 ;
      VIA 218.5 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 48.795 219.29 49.125 ;
      VIA 218.5 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 48.775 219.27 49.145 ;
      VIA 218.5 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 43.355 219.29 43.685 ;
      VIA 218.5 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 43.335 219.27 43.705 ;
      VIA 218.5 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 37.915 219.29 38.245 ;
      VIA 218.5 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 37.895 219.27 38.265 ;
      VIA 218.5 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 32.475 219.29 32.805 ;
      VIA 218.5 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 32.455 219.27 32.825 ;
      VIA 218.5 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 27.035 219.29 27.365 ;
      VIA 218.5 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 27.015 219.27 27.385 ;
      VIA 218.5 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 21.595 219.29 21.925 ;
      VIA 218.5 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 21.575 219.27 21.945 ;
      VIA 218.5 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 16.155 219.29 16.485 ;
      VIA 218.5 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 16.135 219.27 16.505 ;
      VIA 218.5 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 10.715 219.29 11.045 ;
      VIA 218.5 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 10.695 219.27 11.065 ;
      VIA 218.5 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 5.275 219.29 5.605 ;
      VIA 218.5 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 5.255 219.27 5.625 ;
      VIA 218.5 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 418.715 192.15 419.045 ;
      VIA 191.36 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 418.695 192.13 419.065 ;
      VIA 191.36 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 413.275 192.15 413.605 ;
      VIA 191.36 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 413.255 192.13 413.625 ;
      VIA 191.36 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 407.835 192.15 408.165 ;
      VIA 191.36 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 407.815 192.13 408.185 ;
      VIA 191.36 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 402.395 192.15 402.725 ;
      VIA 191.36 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 402.375 192.13 402.745 ;
      VIA 191.36 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 396.955 192.15 397.285 ;
      VIA 191.36 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 396.935 192.13 397.305 ;
      VIA 191.36 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 391.515 192.15 391.845 ;
      VIA 191.36 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 391.495 192.13 391.865 ;
      VIA 191.36 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 386.075 192.15 386.405 ;
      VIA 191.36 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 386.055 192.13 386.425 ;
      VIA 191.36 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 380.635 192.15 380.965 ;
      VIA 191.36 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 380.615 192.13 380.985 ;
      VIA 191.36 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 375.195 192.15 375.525 ;
      VIA 191.36 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 375.175 192.13 375.545 ;
      VIA 191.36 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 369.755 192.15 370.085 ;
      VIA 191.36 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 369.735 192.13 370.105 ;
      VIA 191.36 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 364.315 192.15 364.645 ;
      VIA 191.36 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 364.295 192.13 364.665 ;
      VIA 191.36 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 358.875 192.15 359.205 ;
      VIA 191.36 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 358.855 192.13 359.225 ;
      VIA 191.36 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 353.435 192.15 353.765 ;
      VIA 191.36 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 353.415 192.13 353.785 ;
      VIA 191.36 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 347.995 192.15 348.325 ;
      VIA 191.36 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 347.975 192.13 348.345 ;
      VIA 191.36 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 342.555 192.15 342.885 ;
      VIA 191.36 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 342.535 192.13 342.905 ;
      VIA 191.36 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 337.115 192.15 337.445 ;
      VIA 191.36 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 337.095 192.13 337.465 ;
      VIA 191.36 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 331.675 192.15 332.005 ;
      VIA 191.36 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 331.655 192.13 332.025 ;
      VIA 191.36 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 326.235 192.15 326.565 ;
      VIA 191.36 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 326.215 192.13 326.585 ;
      VIA 191.36 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 320.795 192.15 321.125 ;
      VIA 191.36 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 320.775 192.13 321.145 ;
      VIA 191.36 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 315.355 192.15 315.685 ;
      VIA 191.36 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 315.335 192.13 315.705 ;
      VIA 191.36 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 309.915 192.15 310.245 ;
      VIA 191.36 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 309.895 192.13 310.265 ;
      VIA 191.36 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 304.475 192.15 304.805 ;
      VIA 191.36 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 304.455 192.13 304.825 ;
      VIA 191.36 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 299.035 192.15 299.365 ;
      VIA 191.36 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 299.015 192.13 299.385 ;
      VIA 191.36 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 293.595 192.15 293.925 ;
      VIA 191.36 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 293.575 192.13 293.945 ;
      VIA 191.36 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 288.155 192.15 288.485 ;
      VIA 191.36 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 288.135 192.13 288.505 ;
      VIA 191.36 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 282.715 192.15 283.045 ;
      VIA 191.36 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 282.695 192.13 283.065 ;
      VIA 191.36 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 277.275 192.15 277.605 ;
      VIA 191.36 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 277.255 192.13 277.625 ;
      VIA 191.36 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 271.835 192.15 272.165 ;
      VIA 191.36 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 271.815 192.13 272.185 ;
      VIA 191.36 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 266.395 192.15 266.725 ;
      VIA 191.36 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 266.375 192.13 266.745 ;
      VIA 191.36 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 260.955 192.15 261.285 ;
      VIA 191.36 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 260.935 192.13 261.305 ;
      VIA 191.36 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 255.515 192.15 255.845 ;
      VIA 191.36 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 255.495 192.13 255.865 ;
      VIA 191.36 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 250.075 192.15 250.405 ;
      VIA 191.36 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 250.055 192.13 250.425 ;
      VIA 191.36 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 244.635 192.15 244.965 ;
      VIA 191.36 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 244.615 192.13 244.985 ;
      VIA 191.36 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 239.195 192.15 239.525 ;
      VIA 191.36 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 239.175 192.13 239.545 ;
      VIA 191.36 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 233.755 192.15 234.085 ;
      VIA 191.36 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 233.735 192.13 234.105 ;
      VIA 191.36 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 228.315 192.15 228.645 ;
      VIA 191.36 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 228.295 192.13 228.665 ;
      VIA 191.36 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 222.875 192.15 223.205 ;
      VIA 191.36 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 222.855 192.13 223.225 ;
      VIA 191.36 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 217.435 192.15 217.765 ;
      VIA 191.36 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 217.415 192.13 217.785 ;
      VIA 191.36 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 211.995 192.15 212.325 ;
      VIA 191.36 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 211.975 192.13 212.345 ;
      VIA 191.36 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 206.555 192.15 206.885 ;
      VIA 191.36 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 206.535 192.13 206.905 ;
      VIA 191.36 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 201.115 192.15 201.445 ;
      VIA 191.36 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 201.095 192.13 201.465 ;
      VIA 191.36 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 195.675 192.15 196.005 ;
      VIA 191.36 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 195.655 192.13 196.025 ;
      VIA 191.36 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 190.235 192.15 190.565 ;
      VIA 191.36 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 190.215 192.13 190.585 ;
      VIA 191.36 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 184.795 192.15 185.125 ;
      VIA 191.36 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 184.775 192.13 185.145 ;
      VIA 191.36 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 179.355 192.15 179.685 ;
      VIA 191.36 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 179.335 192.13 179.705 ;
      VIA 191.36 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 173.915 192.15 174.245 ;
      VIA 191.36 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 173.895 192.13 174.265 ;
      VIA 191.36 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 168.475 192.15 168.805 ;
      VIA 191.36 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 168.455 192.13 168.825 ;
      VIA 191.36 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 163.035 192.15 163.365 ;
      VIA 191.36 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 163.015 192.13 163.385 ;
      VIA 191.36 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 157.595 192.15 157.925 ;
      VIA 191.36 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 157.575 192.13 157.945 ;
      VIA 191.36 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 152.155 192.15 152.485 ;
      VIA 191.36 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 152.135 192.13 152.505 ;
      VIA 191.36 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 146.715 192.15 147.045 ;
      VIA 191.36 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 146.695 192.13 147.065 ;
      VIA 191.36 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 141.275 192.15 141.605 ;
      VIA 191.36 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 141.255 192.13 141.625 ;
      VIA 191.36 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 135.835 192.15 136.165 ;
      VIA 191.36 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 135.815 192.13 136.185 ;
      VIA 191.36 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 130.395 192.15 130.725 ;
      VIA 191.36 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 130.375 192.13 130.745 ;
      VIA 191.36 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 124.955 192.15 125.285 ;
      VIA 191.36 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 124.935 192.13 125.305 ;
      VIA 191.36 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 119.515 192.15 119.845 ;
      VIA 191.36 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 119.495 192.13 119.865 ;
      VIA 191.36 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 114.075 192.15 114.405 ;
      VIA 191.36 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 114.055 192.13 114.425 ;
      VIA 191.36 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 108.635 192.15 108.965 ;
      VIA 191.36 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 108.615 192.13 108.985 ;
      VIA 191.36 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 103.195 192.15 103.525 ;
      VIA 191.36 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 103.175 192.13 103.545 ;
      VIA 191.36 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 97.755 192.15 98.085 ;
      VIA 191.36 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 97.735 192.13 98.105 ;
      VIA 191.36 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 92.315 192.15 92.645 ;
      VIA 191.36 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 92.295 192.13 92.665 ;
      VIA 191.36 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 86.875 192.15 87.205 ;
      VIA 191.36 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 86.855 192.13 87.225 ;
      VIA 191.36 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 81.435 192.15 81.765 ;
      VIA 191.36 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 81.415 192.13 81.785 ;
      VIA 191.36 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 75.995 192.15 76.325 ;
      VIA 191.36 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 75.975 192.13 76.345 ;
      VIA 191.36 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 70.555 192.15 70.885 ;
      VIA 191.36 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 70.535 192.13 70.905 ;
      VIA 191.36 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 65.115 192.15 65.445 ;
      VIA 191.36 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 65.095 192.13 65.465 ;
      VIA 191.36 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 59.675 192.15 60.005 ;
      VIA 191.36 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 59.655 192.13 60.025 ;
      VIA 191.36 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 54.235 192.15 54.565 ;
      VIA 191.36 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 54.215 192.13 54.585 ;
      VIA 191.36 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 48.795 192.15 49.125 ;
      VIA 191.36 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 48.775 192.13 49.145 ;
      VIA 191.36 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 43.355 192.15 43.685 ;
      VIA 191.36 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 43.335 192.13 43.705 ;
      VIA 191.36 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 37.915 192.15 38.245 ;
      VIA 191.36 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 37.895 192.13 38.265 ;
      VIA 191.36 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 32.475 192.15 32.805 ;
      VIA 191.36 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 32.455 192.13 32.825 ;
      VIA 191.36 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 27.035 192.15 27.365 ;
      VIA 191.36 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 27.015 192.13 27.385 ;
      VIA 191.36 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 21.595 192.15 21.925 ;
      VIA 191.36 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 21.575 192.13 21.945 ;
      VIA 191.36 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 16.155 192.15 16.485 ;
      VIA 191.36 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 16.135 192.13 16.505 ;
      VIA 191.36 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 10.715 192.15 11.045 ;
      VIA 191.36 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 10.695 192.13 11.065 ;
      VIA 191.36 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 5.275 192.15 5.605 ;
      VIA 191.36 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 5.255 192.13 5.625 ;
      VIA 191.36 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 418.715 165.01 419.045 ;
      VIA 164.22 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 418.695 164.99 419.065 ;
      VIA 164.22 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 413.275 165.01 413.605 ;
      VIA 164.22 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 413.255 164.99 413.625 ;
      VIA 164.22 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 407.835 165.01 408.165 ;
      VIA 164.22 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 407.815 164.99 408.185 ;
      VIA 164.22 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 402.395 165.01 402.725 ;
      VIA 164.22 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 402.375 164.99 402.745 ;
      VIA 164.22 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 396.955 165.01 397.285 ;
      VIA 164.22 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 396.935 164.99 397.305 ;
      VIA 164.22 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 391.515 165.01 391.845 ;
      VIA 164.22 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 391.495 164.99 391.865 ;
      VIA 164.22 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 386.075 165.01 386.405 ;
      VIA 164.22 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 386.055 164.99 386.425 ;
      VIA 164.22 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 380.635 165.01 380.965 ;
      VIA 164.22 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 380.615 164.99 380.985 ;
      VIA 164.22 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 375.195 165.01 375.525 ;
      VIA 164.22 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 375.175 164.99 375.545 ;
      VIA 164.22 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 369.755 165.01 370.085 ;
      VIA 164.22 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 369.735 164.99 370.105 ;
      VIA 164.22 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 364.315 165.01 364.645 ;
      VIA 164.22 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 364.295 164.99 364.665 ;
      VIA 164.22 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 358.875 165.01 359.205 ;
      VIA 164.22 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 358.855 164.99 359.225 ;
      VIA 164.22 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 353.435 165.01 353.765 ;
      VIA 164.22 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 353.415 164.99 353.785 ;
      VIA 164.22 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 347.995 165.01 348.325 ;
      VIA 164.22 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 347.975 164.99 348.345 ;
      VIA 164.22 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 342.555 165.01 342.885 ;
      VIA 164.22 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 342.535 164.99 342.905 ;
      VIA 164.22 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 337.115 165.01 337.445 ;
      VIA 164.22 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 337.095 164.99 337.465 ;
      VIA 164.22 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 331.675 165.01 332.005 ;
      VIA 164.22 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 331.655 164.99 332.025 ;
      VIA 164.22 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 326.235 165.01 326.565 ;
      VIA 164.22 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 326.215 164.99 326.585 ;
      VIA 164.22 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 320.795 165.01 321.125 ;
      VIA 164.22 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 320.775 164.99 321.145 ;
      VIA 164.22 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 315.355 165.01 315.685 ;
      VIA 164.22 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 315.335 164.99 315.705 ;
      VIA 164.22 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 309.915 165.01 310.245 ;
      VIA 164.22 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 309.895 164.99 310.265 ;
      VIA 164.22 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 304.475 165.01 304.805 ;
      VIA 164.22 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 304.455 164.99 304.825 ;
      VIA 164.22 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 299.035 165.01 299.365 ;
      VIA 164.22 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 299.015 164.99 299.385 ;
      VIA 164.22 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 293.595 165.01 293.925 ;
      VIA 164.22 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 293.575 164.99 293.945 ;
      VIA 164.22 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 288.155 165.01 288.485 ;
      VIA 164.22 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 288.135 164.99 288.505 ;
      VIA 164.22 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 282.715 165.01 283.045 ;
      VIA 164.22 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 282.695 164.99 283.065 ;
      VIA 164.22 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 277.275 165.01 277.605 ;
      VIA 164.22 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 277.255 164.99 277.625 ;
      VIA 164.22 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 271.835 165.01 272.165 ;
      VIA 164.22 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 271.815 164.99 272.185 ;
      VIA 164.22 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 266.395 165.01 266.725 ;
      VIA 164.22 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 266.375 164.99 266.745 ;
      VIA 164.22 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 260.955 165.01 261.285 ;
      VIA 164.22 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 260.935 164.99 261.305 ;
      VIA 164.22 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 255.515 165.01 255.845 ;
      VIA 164.22 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 255.495 164.99 255.865 ;
      VIA 164.22 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 250.075 165.01 250.405 ;
      VIA 164.22 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 250.055 164.99 250.425 ;
      VIA 164.22 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 244.635 165.01 244.965 ;
      VIA 164.22 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 244.615 164.99 244.985 ;
      VIA 164.22 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 239.195 165.01 239.525 ;
      VIA 164.22 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 239.175 164.99 239.545 ;
      VIA 164.22 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 233.755 165.01 234.085 ;
      VIA 164.22 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 233.735 164.99 234.105 ;
      VIA 164.22 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 228.315 165.01 228.645 ;
      VIA 164.22 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 228.295 164.99 228.665 ;
      VIA 164.22 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 222.875 165.01 223.205 ;
      VIA 164.22 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 222.855 164.99 223.225 ;
      VIA 164.22 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 217.435 165.01 217.765 ;
      VIA 164.22 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 217.415 164.99 217.785 ;
      VIA 164.22 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 211.995 165.01 212.325 ;
      VIA 164.22 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 211.975 164.99 212.345 ;
      VIA 164.22 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 206.555 165.01 206.885 ;
      VIA 164.22 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 206.535 164.99 206.905 ;
      VIA 164.22 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 201.115 165.01 201.445 ;
      VIA 164.22 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 201.095 164.99 201.465 ;
      VIA 164.22 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 195.675 165.01 196.005 ;
      VIA 164.22 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 195.655 164.99 196.025 ;
      VIA 164.22 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 190.235 165.01 190.565 ;
      VIA 164.22 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 190.215 164.99 190.585 ;
      VIA 164.22 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 184.795 165.01 185.125 ;
      VIA 164.22 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 184.775 164.99 185.145 ;
      VIA 164.22 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 179.355 165.01 179.685 ;
      VIA 164.22 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 179.335 164.99 179.705 ;
      VIA 164.22 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 173.915 165.01 174.245 ;
      VIA 164.22 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 173.895 164.99 174.265 ;
      VIA 164.22 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 168.475 165.01 168.805 ;
      VIA 164.22 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 168.455 164.99 168.825 ;
      VIA 164.22 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 163.035 165.01 163.365 ;
      VIA 164.22 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 163.015 164.99 163.385 ;
      VIA 164.22 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 157.595 165.01 157.925 ;
      VIA 164.22 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 157.575 164.99 157.945 ;
      VIA 164.22 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 152.155 165.01 152.485 ;
      VIA 164.22 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 152.135 164.99 152.505 ;
      VIA 164.22 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 146.715 165.01 147.045 ;
      VIA 164.22 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 146.695 164.99 147.065 ;
      VIA 164.22 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 141.275 165.01 141.605 ;
      VIA 164.22 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 141.255 164.99 141.625 ;
      VIA 164.22 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 135.835 165.01 136.165 ;
      VIA 164.22 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 135.815 164.99 136.185 ;
      VIA 164.22 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 130.395 165.01 130.725 ;
      VIA 164.22 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 130.375 164.99 130.745 ;
      VIA 164.22 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 124.955 165.01 125.285 ;
      VIA 164.22 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 124.935 164.99 125.305 ;
      VIA 164.22 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 119.515 165.01 119.845 ;
      VIA 164.22 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 119.495 164.99 119.865 ;
      VIA 164.22 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 114.075 165.01 114.405 ;
      VIA 164.22 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 114.055 164.99 114.425 ;
      VIA 164.22 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 108.635 165.01 108.965 ;
      VIA 164.22 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 108.615 164.99 108.985 ;
      VIA 164.22 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 103.195 165.01 103.525 ;
      VIA 164.22 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 103.175 164.99 103.545 ;
      VIA 164.22 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 97.755 165.01 98.085 ;
      VIA 164.22 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 97.735 164.99 98.105 ;
      VIA 164.22 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 92.315 165.01 92.645 ;
      VIA 164.22 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 92.295 164.99 92.665 ;
      VIA 164.22 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 86.875 165.01 87.205 ;
      VIA 164.22 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 86.855 164.99 87.225 ;
      VIA 164.22 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 81.435 165.01 81.765 ;
      VIA 164.22 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 81.415 164.99 81.785 ;
      VIA 164.22 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 75.995 165.01 76.325 ;
      VIA 164.22 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 75.975 164.99 76.345 ;
      VIA 164.22 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 70.555 165.01 70.885 ;
      VIA 164.22 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 70.535 164.99 70.905 ;
      VIA 164.22 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 65.115 165.01 65.445 ;
      VIA 164.22 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 65.095 164.99 65.465 ;
      VIA 164.22 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 59.675 165.01 60.005 ;
      VIA 164.22 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 59.655 164.99 60.025 ;
      VIA 164.22 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 54.235 165.01 54.565 ;
      VIA 164.22 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 54.215 164.99 54.585 ;
      VIA 164.22 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 48.795 165.01 49.125 ;
      VIA 164.22 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 48.775 164.99 49.145 ;
      VIA 164.22 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 43.355 165.01 43.685 ;
      VIA 164.22 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 43.335 164.99 43.705 ;
      VIA 164.22 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 37.915 165.01 38.245 ;
      VIA 164.22 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 37.895 164.99 38.265 ;
      VIA 164.22 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 32.475 165.01 32.805 ;
      VIA 164.22 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 32.455 164.99 32.825 ;
      VIA 164.22 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 27.035 165.01 27.365 ;
      VIA 164.22 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 27.015 164.99 27.385 ;
      VIA 164.22 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 21.595 165.01 21.925 ;
      VIA 164.22 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 21.575 164.99 21.945 ;
      VIA 164.22 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 16.155 165.01 16.485 ;
      VIA 164.22 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 16.135 164.99 16.505 ;
      VIA 164.22 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 10.715 165.01 11.045 ;
      VIA 164.22 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 10.695 164.99 11.065 ;
      VIA 164.22 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 5.275 165.01 5.605 ;
      VIA 164.22 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 5.255 164.99 5.625 ;
      VIA 164.22 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 418.715 137.87 419.045 ;
      VIA 137.08 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 418.695 137.85 419.065 ;
      VIA 137.08 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 413.275 137.87 413.605 ;
      VIA 137.08 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 413.255 137.85 413.625 ;
      VIA 137.08 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 407.835 137.87 408.165 ;
      VIA 137.08 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 407.815 137.85 408.185 ;
      VIA 137.08 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 402.395 137.87 402.725 ;
      VIA 137.08 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 402.375 137.85 402.745 ;
      VIA 137.08 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 396.955 137.87 397.285 ;
      VIA 137.08 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 396.935 137.85 397.305 ;
      VIA 137.08 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 391.515 137.87 391.845 ;
      VIA 137.08 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 391.495 137.85 391.865 ;
      VIA 137.08 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 386.075 137.87 386.405 ;
      VIA 137.08 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 386.055 137.85 386.425 ;
      VIA 137.08 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 380.635 137.87 380.965 ;
      VIA 137.08 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 380.615 137.85 380.985 ;
      VIA 137.08 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 375.195 137.87 375.525 ;
      VIA 137.08 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 375.175 137.85 375.545 ;
      VIA 137.08 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 369.755 137.87 370.085 ;
      VIA 137.08 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 369.735 137.85 370.105 ;
      VIA 137.08 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 364.315 137.87 364.645 ;
      VIA 137.08 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 364.295 137.85 364.665 ;
      VIA 137.08 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 358.875 137.87 359.205 ;
      VIA 137.08 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 358.855 137.85 359.225 ;
      VIA 137.08 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 353.435 137.87 353.765 ;
      VIA 137.08 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 353.415 137.85 353.785 ;
      VIA 137.08 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 347.995 137.87 348.325 ;
      VIA 137.08 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 347.975 137.85 348.345 ;
      VIA 137.08 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 342.555 137.87 342.885 ;
      VIA 137.08 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 342.535 137.85 342.905 ;
      VIA 137.08 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 337.115 137.87 337.445 ;
      VIA 137.08 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 337.095 137.85 337.465 ;
      VIA 137.08 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 331.675 137.87 332.005 ;
      VIA 137.08 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 331.655 137.85 332.025 ;
      VIA 137.08 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 326.235 137.87 326.565 ;
      VIA 137.08 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 326.215 137.85 326.585 ;
      VIA 137.08 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 320.795 137.87 321.125 ;
      VIA 137.08 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 320.775 137.85 321.145 ;
      VIA 137.08 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 315.355 137.87 315.685 ;
      VIA 137.08 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 315.335 137.85 315.705 ;
      VIA 137.08 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 309.915 137.87 310.245 ;
      VIA 137.08 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 309.895 137.85 310.265 ;
      VIA 137.08 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 304.475 137.87 304.805 ;
      VIA 137.08 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 304.455 137.85 304.825 ;
      VIA 137.08 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 299.035 137.87 299.365 ;
      VIA 137.08 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 299.015 137.85 299.385 ;
      VIA 137.08 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 293.595 137.87 293.925 ;
      VIA 137.08 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 293.575 137.85 293.945 ;
      VIA 137.08 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 288.155 137.87 288.485 ;
      VIA 137.08 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 288.135 137.85 288.505 ;
      VIA 137.08 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 282.715 137.87 283.045 ;
      VIA 137.08 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 282.695 137.85 283.065 ;
      VIA 137.08 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 277.275 137.87 277.605 ;
      VIA 137.08 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 277.255 137.85 277.625 ;
      VIA 137.08 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 271.835 137.87 272.165 ;
      VIA 137.08 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 271.815 137.85 272.185 ;
      VIA 137.08 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 266.395 137.87 266.725 ;
      VIA 137.08 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 266.375 137.85 266.745 ;
      VIA 137.08 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 260.955 137.87 261.285 ;
      VIA 137.08 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 260.935 137.85 261.305 ;
      VIA 137.08 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 255.515 137.87 255.845 ;
      VIA 137.08 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 255.495 137.85 255.865 ;
      VIA 137.08 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 250.075 137.87 250.405 ;
      VIA 137.08 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 250.055 137.85 250.425 ;
      VIA 137.08 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 244.635 137.87 244.965 ;
      VIA 137.08 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 244.615 137.85 244.985 ;
      VIA 137.08 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 239.195 137.87 239.525 ;
      VIA 137.08 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 239.175 137.85 239.545 ;
      VIA 137.08 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 233.755 137.87 234.085 ;
      VIA 137.08 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 233.735 137.85 234.105 ;
      VIA 137.08 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 228.315 137.87 228.645 ;
      VIA 137.08 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 228.295 137.85 228.665 ;
      VIA 137.08 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 222.875 137.87 223.205 ;
      VIA 137.08 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 222.855 137.85 223.225 ;
      VIA 137.08 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 217.435 137.87 217.765 ;
      VIA 137.08 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 217.415 137.85 217.785 ;
      VIA 137.08 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 211.995 137.87 212.325 ;
      VIA 137.08 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 211.975 137.85 212.345 ;
      VIA 137.08 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 206.555 137.87 206.885 ;
      VIA 137.08 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 206.535 137.85 206.905 ;
      VIA 137.08 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 201.115 137.87 201.445 ;
      VIA 137.08 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 201.095 137.85 201.465 ;
      VIA 137.08 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 195.675 137.87 196.005 ;
      VIA 137.08 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 195.655 137.85 196.025 ;
      VIA 137.08 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 190.235 137.87 190.565 ;
      VIA 137.08 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 190.215 137.85 190.585 ;
      VIA 137.08 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 184.795 137.87 185.125 ;
      VIA 137.08 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 184.775 137.85 185.145 ;
      VIA 137.08 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 179.355 137.87 179.685 ;
      VIA 137.08 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 179.335 137.85 179.705 ;
      VIA 137.08 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 173.915 137.87 174.245 ;
      VIA 137.08 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 173.895 137.85 174.265 ;
      VIA 137.08 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 168.475 137.87 168.805 ;
      VIA 137.08 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 168.455 137.85 168.825 ;
      VIA 137.08 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 163.035 137.87 163.365 ;
      VIA 137.08 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 163.015 137.85 163.385 ;
      VIA 137.08 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 157.595 137.87 157.925 ;
      VIA 137.08 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 157.575 137.85 157.945 ;
      VIA 137.08 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 152.155 137.87 152.485 ;
      VIA 137.08 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 152.135 137.85 152.505 ;
      VIA 137.08 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 146.715 137.87 147.045 ;
      VIA 137.08 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 146.695 137.85 147.065 ;
      VIA 137.08 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 141.275 137.87 141.605 ;
      VIA 137.08 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 141.255 137.85 141.625 ;
      VIA 137.08 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 135.835 137.87 136.165 ;
      VIA 137.08 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 135.815 137.85 136.185 ;
      VIA 137.08 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 130.395 137.87 130.725 ;
      VIA 137.08 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 130.375 137.85 130.745 ;
      VIA 137.08 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 124.955 137.87 125.285 ;
      VIA 137.08 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 124.935 137.85 125.305 ;
      VIA 137.08 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 119.515 137.87 119.845 ;
      VIA 137.08 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 119.495 137.85 119.865 ;
      VIA 137.08 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 114.075 137.87 114.405 ;
      VIA 137.08 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 114.055 137.85 114.425 ;
      VIA 137.08 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 108.635 137.87 108.965 ;
      VIA 137.08 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 108.615 137.85 108.985 ;
      VIA 137.08 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 103.195 137.87 103.525 ;
      VIA 137.08 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 103.175 137.85 103.545 ;
      VIA 137.08 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 97.755 137.87 98.085 ;
      VIA 137.08 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 97.735 137.85 98.105 ;
      VIA 137.08 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 92.315 137.87 92.645 ;
      VIA 137.08 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 92.295 137.85 92.665 ;
      VIA 137.08 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 86.875 137.87 87.205 ;
      VIA 137.08 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 86.855 137.85 87.225 ;
      VIA 137.08 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 81.435 137.87 81.765 ;
      VIA 137.08 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 81.415 137.85 81.785 ;
      VIA 137.08 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 75.995 137.87 76.325 ;
      VIA 137.08 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 75.975 137.85 76.345 ;
      VIA 137.08 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 70.555 137.87 70.885 ;
      VIA 137.08 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 70.535 137.85 70.905 ;
      VIA 137.08 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 65.115 137.87 65.445 ;
      VIA 137.08 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 65.095 137.85 65.465 ;
      VIA 137.08 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 59.675 137.87 60.005 ;
      VIA 137.08 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 59.655 137.85 60.025 ;
      VIA 137.08 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 54.235 137.87 54.565 ;
      VIA 137.08 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 54.215 137.85 54.585 ;
      VIA 137.08 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 48.795 137.87 49.125 ;
      VIA 137.08 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 48.775 137.85 49.145 ;
      VIA 137.08 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 43.355 137.87 43.685 ;
      VIA 137.08 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 43.335 137.85 43.705 ;
      VIA 137.08 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 37.915 137.87 38.245 ;
      VIA 137.08 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 37.895 137.85 38.265 ;
      VIA 137.08 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 32.475 137.87 32.805 ;
      VIA 137.08 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 32.455 137.85 32.825 ;
      VIA 137.08 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 27.035 137.87 27.365 ;
      VIA 137.08 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 27.015 137.85 27.385 ;
      VIA 137.08 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 21.595 137.87 21.925 ;
      VIA 137.08 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 21.575 137.85 21.945 ;
      VIA 137.08 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 16.155 137.87 16.485 ;
      VIA 137.08 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 16.135 137.85 16.505 ;
      VIA 137.08 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 10.715 137.87 11.045 ;
      VIA 137.08 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 10.695 137.85 11.065 ;
      VIA 137.08 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 5.275 137.87 5.605 ;
      VIA 137.08 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 5.255 137.85 5.625 ;
      VIA 137.08 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 418.715 110.73 419.045 ;
      VIA 109.94 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 418.695 110.71 419.065 ;
      VIA 109.94 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 413.275 110.73 413.605 ;
      VIA 109.94 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 413.255 110.71 413.625 ;
      VIA 109.94 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 407.835 110.73 408.165 ;
      VIA 109.94 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 407.815 110.71 408.185 ;
      VIA 109.94 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 402.395 110.73 402.725 ;
      VIA 109.94 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 402.375 110.71 402.745 ;
      VIA 109.94 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 396.955 110.73 397.285 ;
      VIA 109.94 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 396.935 110.71 397.305 ;
      VIA 109.94 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 391.515 110.73 391.845 ;
      VIA 109.94 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 391.495 110.71 391.865 ;
      VIA 109.94 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 386.075 110.73 386.405 ;
      VIA 109.94 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 386.055 110.71 386.425 ;
      VIA 109.94 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 380.635 110.73 380.965 ;
      VIA 109.94 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 380.615 110.71 380.985 ;
      VIA 109.94 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 375.195 110.73 375.525 ;
      VIA 109.94 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 375.175 110.71 375.545 ;
      VIA 109.94 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 369.755 110.73 370.085 ;
      VIA 109.94 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 369.735 110.71 370.105 ;
      VIA 109.94 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 364.315 110.73 364.645 ;
      VIA 109.94 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 364.295 110.71 364.665 ;
      VIA 109.94 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 358.875 110.73 359.205 ;
      VIA 109.94 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 358.855 110.71 359.225 ;
      VIA 109.94 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 353.435 110.73 353.765 ;
      VIA 109.94 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 353.415 110.71 353.785 ;
      VIA 109.94 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 347.995 110.73 348.325 ;
      VIA 109.94 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 347.975 110.71 348.345 ;
      VIA 109.94 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 342.555 110.73 342.885 ;
      VIA 109.94 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 342.535 110.71 342.905 ;
      VIA 109.94 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 337.115 110.73 337.445 ;
      VIA 109.94 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 337.095 110.71 337.465 ;
      VIA 109.94 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 331.675 110.73 332.005 ;
      VIA 109.94 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 331.655 110.71 332.025 ;
      VIA 109.94 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 326.235 110.73 326.565 ;
      VIA 109.94 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 326.215 110.71 326.585 ;
      VIA 109.94 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 320.795 110.73 321.125 ;
      VIA 109.94 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 320.775 110.71 321.145 ;
      VIA 109.94 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 315.355 110.73 315.685 ;
      VIA 109.94 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 315.335 110.71 315.705 ;
      VIA 109.94 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 309.915 110.73 310.245 ;
      VIA 109.94 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 309.895 110.71 310.265 ;
      VIA 109.94 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 304.475 110.73 304.805 ;
      VIA 109.94 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 304.455 110.71 304.825 ;
      VIA 109.94 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 299.035 110.73 299.365 ;
      VIA 109.94 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 299.015 110.71 299.385 ;
      VIA 109.94 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 293.595 110.73 293.925 ;
      VIA 109.94 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 293.575 110.71 293.945 ;
      VIA 109.94 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 288.155 110.73 288.485 ;
      VIA 109.94 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 288.135 110.71 288.505 ;
      VIA 109.94 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 282.715 110.73 283.045 ;
      VIA 109.94 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 282.695 110.71 283.065 ;
      VIA 109.94 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 277.275 110.73 277.605 ;
      VIA 109.94 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 277.255 110.71 277.625 ;
      VIA 109.94 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 271.835 110.73 272.165 ;
      VIA 109.94 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 271.815 110.71 272.185 ;
      VIA 109.94 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 266.395 110.73 266.725 ;
      VIA 109.94 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 266.375 110.71 266.745 ;
      VIA 109.94 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 260.955 110.73 261.285 ;
      VIA 109.94 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 260.935 110.71 261.305 ;
      VIA 109.94 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 255.515 110.73 255.845 ;
      VIA 109.94 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 255.495 110.71 255.865 ;
      VIA 109.94 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 250.075 110.73 250.405 ;
      VIA 109.94 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 250.055 110.71 250.425 ;
      VIA 109.94 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 244.635 110.73 244.965 ;
      VIA 109.94 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 244.615 110.71 244.985 ;
      VIA 109.94 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 239.195 110.73 239.525 ;
      VIA 109.94 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 239.175 110.71 239.545 ;
      VIA 109.94 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 233.755 110.73 234.085 ;
      VIA 109.94 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 233.735 110.71 234.105 ;
      VIA 109.94 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 228.315 110.73 228.645 ;
      VIA 109.94 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 228.295 110.71 228.665 ;
      VIA 109.94 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 222.875 110.73 223.205 ;
      VIA 109.94 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 222.855 110.71 223.225 ;
      VIA 109.94 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 217.435 110.73 217.765 ;
      VIA 109.94 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 217.415 110.71 217.785 ;
      VIA 109.94 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 211.995 110.73 212.325 ;
      VIA 109.94 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 211.975 110.71 212.345 ;
      VIA 109.94 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 206.555 110.73 206.885 ;
      VIA 109.94 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 206.535 110.71 206.905 ;
      VIA 109.94 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 201.115 110.73 201.445 ;
      VIA 109.94 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 201.095 110.71 201.465 ;
      VIA 109.94 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 195.675 110.73 196.005 ;
      VIA 109.94 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 195.655 110.71 196.025 ;
      VIA 109.94 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 190.235 110.73 190.565 ;
      VIA 109.94 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 190.215 110.71 190.585 ;
      VIA 109.94 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 184.795 110.73 185.125 ;
      VIA 109.94 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 184.775 110.71 185.145 ;
      VIA 109.94 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 179.355 110.73 179.685 ;
      VIA 109.94 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 179.335 110.71 179.705 ;
      VIA 109.94 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 173.915 110.73 174.245 ;
      VIA 109.94 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 173.895 110.71 174.265 ;
      VIA 109.94 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 168.475 110.73 168.805 ;
      VIA 109.94 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 168.455 110.71 168.825 ;
      VIA 109.94 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 163.035 110.73 163.365 ;
      VIA 109.94 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 163.015 110.71 163.385 ;
      VIA 109.94 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 157.595 110.73 157.925 ;
      VIA 109.94 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 157.575 110.71 157.945 ;
      VIA 109.94 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 152.155 110.73 152.485 ;
      VIA 109.94 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 152.135 110.71 152.505 ;
      VIA 109.94 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 146.715 110.73 147.045 ;
      VIA 109.94 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 146.695 110.71 147.065 ;
      VIA 109.94 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 141.275 110.73 141.605 ;
      VIA 109.94 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 141.255 110.71 141.625 ;
      VIA 109.94 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 135.835 110.73 136.165 ;
      VIA 109.94 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 135.815 110.71 136.185 ;
      VIA 109.94 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 130.395 110.73 130.725 ;
      VIA 109.94 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 130.375 110.71 130.745 ;
      VIA 109.94 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 124.955 110.73 125.285 ;
      VIA 109.94 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 124.935 110.71 125.305 ;
      VIA 109.94 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 119.515 110.73 119.845 ;
      VIA 109.94 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 119.495 110.71 119.865 ;
      VIA 109.94 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 114.075 110.73 114.405 ;
      VIA 109.94 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 114.055 110.71 114.425 ;
      VIA 109.94 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 108.635 110.73 108.965 ;
      VIA 109.94 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 108.615 110.71 108.985 ;
      VIA 109.94 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 103.195 110.73 103.525 ;
      VIA 109.94 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 103.175 110.71 103.545 ;
      VIA 109.94 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 97.755 110.73 98.085 ;
      VIA 109.94 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 97.735 110.71 98.105 ;
      VIA 109.94 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 92.315 110.73 92.645 ;
      VIA 109.94 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 92.295 110.71 92.665 ;
      VIA 109.94 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 86.875 110.73 87.205 ;
      VIA 109.94 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 86.855 110.71 87.225 ;
      VIA 109.94 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 81.435 110.73 81.765 ;
      VIA 109.94 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 81.415 110.71 81.785 ;
      VIA 109.94 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 75.995 110.73 76.325 ;
      VIA 109.94 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 75.975 110.71 76.345 ;
      VIA 109.94 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 70.555 110.73 70.885 ;
      VIA 109.94 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 70.535 110.71 70.905 ;
      VIA 109.94 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 65.115 110.73 65.445 ;
      VIA 109.94 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 65.095 110.71 65.465 ;
      VIA 109.94 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 59.675 110.73 60.005 ;
      VIA 109.94 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 59.655 110.71 60.025 ;
      VIA 109.94 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 54.235 110.73 54.565 ;
      VIA 109.94 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 54.215 110.71 54.585 ;
      VIA 109.94 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 48.795 110.73 49.125 ;
      VIA 109.94 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 48.775 110.71 49.145 ;
      VIA 109.94 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 43.355 110.73 43.685 ;
      VIA 109.94 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 43.335 110.71 43.705 ;
      VIA 109.94 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 37.915 110.73 38.245 ;
      VIA 109.94 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 37.895 110.71 38.265 ;
      VIA 109.94 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 32.475 110.73 32.805 ;
      VIA 109.94 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 32.455 110.71 32.825 ;
      VIA 109.94 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 27.035 110.73 27.365 ;
      VIA 109.94 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 27.015 110.71 27.385 ;
      VIA 109.94 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 21.595 110.73 21.925 ;
      VIA 109.94 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 21.575 110.71 21.945 ;
      VIA 109.94 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 16.155 110.73 16.485 ;
      VIA 109.94 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 16.135 110.71 16.505 ;
      VIA 109.94 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 10.715 110.73 11.045 ;
      VIA 109.94 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 10.695 110.71 11.065 ;
      VIA 109.94 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 5.275 110.73 5.605 ;
      VIA 109.94 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 5.255 110.71 5.625 ;
      VIA 109.94 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 418.715 83.59 419.045 ;
      VIA 82.8 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 418.695 83.57 419.065 ;
      VIA 82.8 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 413.275 83.59 413.605 ;
      VIA 82.8 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 413.255 83.57 413.625 ;
      VIA 82.8 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 407.835 83.59 408.165 ;
      VIA 82.8 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 407.815 83.57 408.185 ;
      VIA 82.8 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 402.395 83.59 402.725 ;
      VIA 82.8 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 402.375 83.57 402.745 ;
      VIA 82.8 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 396.955 83.59 397.285 ;
      VIA 82.8 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 396.935 83.57 397.305 ;
      VIA 82.8 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 391.515 83.59 391.845 ;
      VIA 82.8 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 391.495 83.57 391.865 ;
      VIA 82.8 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 386.075 83.59 386.405 ;
      VIA 82.8 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 386.055 83.57 386.425 ;
      VIA 82.8 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 380.635 83.59 380.965 ;
      VIA 82.8 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 380.615 83.57 380.985 ;
      VIA 82.8 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 375.195 83.59 375.525 ;
      VIA 82.8 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 375.175 83.57 375.545 ;
      VIA 82.8 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 369.755 83.59 370.085 ;
      VIA 82.8 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 369.735 83.57 370.105 ;
      VIA 82.8 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 364.315 83.59 364.645 ;
      VIA 82.8 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 364.295 83.57 364.665 ;
      VIA 82.8 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 358.875 83.59 359.205 ;
      VIA 82.8 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 358.855 83.57 359.225 ;
      VIA 82.8 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 353.435 83.59 353.765 ;
      VIA 82.8 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 353.415 83.57 353.785 ;
      VIA 82.8 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 347.995 83.59 348.325 ;
      VIA 82.8 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 347.975 83.57 348.345 ;
      VIA 82.8 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 342.555 83.59 342.885 ;
      VIA 82.8 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 342.535 83.57 342.905 ;
      VIA 82.8 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 337.115 83.59 337.445 ;
      VIA 82.8 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 337.095 83.57 337.465 ;
      VIA 82.8 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 331.675 83.59 332.005 ;
      VIA 82.8 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 331.655 83.57 332.025 ;
      VIA 82.8 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 326.235 83.59 326.565 ;
      VIA 82.8 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 326.215 83.57 326.585 ;
      VIA 82.8 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 320.795 83.59 321.125 ;
      VIA 82.8 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 320.775 83.57 321.145 ;
      VIA 82.8 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 315.355 83.59 315.685 ;
      VIA 82.8 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 315.335 83.57 315.705 ;
      VIA 82.8 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 309.915 83.59 310.245 ;
      VIA 82.8 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 309.895 83.57 310.265 ;
      VIA 82.8 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 304.475 83.59 304.805 ;
      VIA 82.8 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 304.455 83.57 304.825 ;
      VIA 82.8 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 299.035 83.59 299.365 ;
      VIA 82.8 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 299.015 83.57 299.385 ;
      VIA 82.8 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 293.595 83.59 293.925 ;
      VIA 82.8 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 293.575 83.57 293.945 ;
      VIA 82.8 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 288.155 83.59 288.485 ;
      VIA 82.8 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 288.135 83.57 288.505 ;
      VIA 82.8 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 282.715 83.59 283.045 ;
      VIA 82.8 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 282.695 83.57 283.065 ;
      VIA 82.8 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 277.275 83.59 277.605 ;
      VIA 82.8 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 277.255 83.57 277.625 ;
      VIA 82.8 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 271.835 83.59 272.165 ;
      VIA 82.8 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 271.815 83.57 272.185 ;
      VIA 82.8 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 266.395 83.59 266.725 ;
      VIA 82.8 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 266.375 83.57 266.745 ;
      VIA 82.8 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 260.955 83.59 261.285 ;
      VIA 82.8 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 260.935 83.57 261.305 ;
      VIA 82.8 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 255.515 83.59 255.845 ;
      VIA 82.8 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 255.495 83.57 255.865 ;
      VIA 82.8 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 250.075 83.59 250.405 ;
      VIA 82.8 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 250.055 83.57 250.425 ;
      VIA 82.8 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 244.635 83.59 244.965 ;
      VIA 82.8 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 244.615 83.57 244.985 ;
      VIA 82.8 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 239.195 83.59 239.525 ;
      VIA 82.8 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 239.175 83.57 239.545 ;
      VIA 82.8 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 233.755 83.59 234.085 ;
      VIA 82.8 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 233.735 83.57 234.105 ;
      VIA 82.8 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 228.315 83.59 228.645 ;
      VIA 82.8 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 228.295 83.57 228.665 ;
      VIA 82.8 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 222.875 83.59 223.205 ;
      VIA 82.8 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 222.855 83.57 223.225 ;
      VIA 82.8 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 217.435 83.59 217.765 ;
      VIA 82.8 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 217.415 83.57 217.785 ;
      VIA 82.8 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 211.995 83.59 212.325 ;
      VIA 82.8 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 211.975 83.57 212.345 ;
      VIA 82.8 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 206.555 83.59 206.885 ;
      VIA 82.8 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 206.535 83.57 206.905 ;
      VIA 82.8 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 201.115 83.59 201.445 ;
      VIA 82.8 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 201.095 83.57 201.465 ;
      VIA 82.8 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 195.675 83.59 196.005 ;
      VIA 82.8 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 195.655 83.57 196.025 ;
      VIA 82.8 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 190.235 83.59 190.565 ;
      VIA 82.8 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 190.215 83.57 190.585 ;
      VIA 82.8 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 184.795 83.59 185.125 ;
      VIA 82.8 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 184.775 83.57 185.145 ;
      VIA 82.8 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 179.355 83.59 179.685 ;
      VIA 82.8 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 179.335 83.57 179.705 ;
      VIA 82.8 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 173.915 83.59 174.245 ;
      VIA 82.8 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 173.895 83.57 174.265 ;
      VIA 82.8 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 168.475 83.59 168.805 ;
      VIA 82.8 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 168.455 83.57 168.825 ;
      VIA 82.8 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 163.035 83.59 163.365 ;
      VIA 82.8 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 163.015 83.57 163.385 ;
      VIA 82.8 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 157.595 83.59 157.925 ;
      VIA 82.8 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 157.575 83.57 157.945 ;
      VIA 82.8 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 152.155 83.59 152.485 ;
      VIA 82.8 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 152.135 83.57 152.505 ;
      VIA 82.8 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 146.715 83.59 147.045 ;
      VIA 82.8 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 146.695 83.57 147.065 ;
      VIA 82.8 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 141.275 83.59 141.605 ;
      VIA 82.8 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 141.255 83.57 141.625 ;
      VIA 82.8 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 135.835 83.59 136.165 ;
      VIA 82.8 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 135.815 83.57 136.185 ;
      VIA 82.8 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 130.395 83.59 130.725 ;
      VIA 82.8 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 130.375 83.57 130.745 ;
      VIA 82.8 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 124.955 83.59 125.285 ;
      VIA 82.8 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 124.935 83.57 125.305 ;
      VIA 82.8 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 119.515 83.59 119.845 ;
      VIA 82.8 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 119.495 83.57 119.865 ;
      VIA 82.8 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 114.075 83.59 114.405 ;
      VIA 82.8 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 114.055 83.57 114.425 ;
      VIA 82.8 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 108.635 83.59 108.965 ;
      VIA 82.8 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 108.615 83.57 108.985 ;
      VIA 82.8 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 103.195 83.59 103.525 ;
      VIA 82.8 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 103.175 83.57 103.545 ;
      VIA 82.8 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 97.755 83.59 98.085 ;
      VIA 82.8 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 97.735 83.57 98.105 ;
      VIA 82.8 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 92.315 83.59 92.645 ;
      VIA 82.8 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 92.295 83.57 92.665 ;
      VIA 82.8 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 86.875 83.59 87.205 ;
      VIA 82.8 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 86.855 83.57 87.225 ;
      VIA 82.8 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 81.435 83.59 81.765 ;
      VIA 82.8 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 81.415 83.57 81.785 ;
      VIA 82.8 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 75.995 83.59 76.325 ;
      VIA 82.8 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 75.975 83.57 76.345 ;
      VIA 82.8 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 70.555 83.59 70.885 ;
      VIA 82.8 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 70.535 83.57 70.905 ;
      VIA 82.8 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 65.115 83.59 65.445 ;
      VIA 82.8 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 65.095 83.57 65.465 ;
      VIA 82.8 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 59.675 83.59 60.005 ;
      VIA 82.8 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 59.655 83.57 60.025 ;
      VIA 82.8 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 54.235 83.59 54.565 ;
      VIA 82.8 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 54.215 83.57 54.585 ;
      VIA 82.8 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 48.795 83.59 49.125 ;
      VIA 82.8 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 48.775 83.57 49.145 ;
      VIA 82.8 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 43.355 83.59 43.685 ;
      VIA 82.8 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 43.335 83.57 43.705 ;
      VIA 82.8 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 37.915 83.59 38.245 ;
      VIA 82.8 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 37.895 83.57 38.265 ;
      VIA 82.8 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 32.475 83.59 32.805 ;
      VIA 82.8 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 32.455 83.57 32.825 ;
      VIA 82.8 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 27.035 83.59 27.365 ;
      VIA 82.8 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 27.015 83.57 27.385 ;
      VIA 82.8 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 21.595 83.59 21.925 ;
      VIA 82.8 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 21.575 83.57 21.945 ;
      VIA 82.8 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 16.155 83.59 16.485 ;
      VIA 82.8 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 16.135 83.57 16.505 ;
      VIA 82.8 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 10.715 83.59 11.045 ;
      VIA 82.8 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 10.695 83.57 11.065 ;
      VIA 82.8 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 5.275 83.59 5.605 ;
      VIA 82.8 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 5.255 83.57 5.625 ;
      VIA 82.8 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 418.715 56.45 419.045 ;
      VIA 55.66 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 418.695 56.43 419.065 ;
      VIA 55.66 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 413.275 56.45 413.605 ;
      VIA 55.66 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 413.255 56.43 413.625 ;
      VIA 55.66 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 407.835 56.45 408.165 ;
      VIA 55.66 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 407.815 56.43 408.185 ;
      VIA 55.66 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 402.395 56.45 402.725 ;
      VIA 55.66 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 402.375 56.43 402.745 ;
      VIA 55.66 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 396.955 56.45 397.285 ;
      VIA 55.66 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 396.935 56.43 397.305 ;
      VIA 55.66 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 391.515 56.45 391.845 ;
      VIA 55.66 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 391.495 56.43 391.865 ;
      VIA 55.66 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 386.075 56.45 386.405 ;
      VIA 55.66 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 386.055 56.43 386.425 ;
      VIA 55.66 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 380.635 56.45 380.965 ;
      VIA 55.66 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 380.615 56.43 380.985 ;
      VIA 55.66 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 375.195 56.45 375.525 ;
      VIA 55.66 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 375.175 56.43 375.545 ;
      VIA 55.66 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 369.755 56.45 370.085 ;
      VIA 55.66 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 369.735 56.43 370.105 ;
      VIA 55.66 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 364.315 56.45 364.645 ;
      VIA 55.66 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 364.295 56.43 364.665 ;
      VIA 55.66 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 358.875 56.45 359.205 ;
      VIA 55.66 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 358.855 56.43 359.225 ;
      VIA 55.66 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 353.435 56.45 353.765 ;
      VIA 55.66 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 353.415 56.43 353.785 ;
      VIA 55.66 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 347.995 56.45 348.325 ;
      VIA 55.66 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 347.975 56.43 348.345 ;
      VIA 55.66 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 342.555 56.45 342.885 ;
      VIA 55.66 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 342.535 56.43 342.905 ;
      VIA 55.66 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 337.115 56.45 337.445 ;
      VIA 55.66 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 337.095 56.43 337.465 ;
      VIA 55.66 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 331.675 56.45 332.005 ;
      VIA 55.66 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 331.655 56.43 332.025 ;
      VIA 55.66 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 326.235 56.45 326.565 ;
      VIA 55.66 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 326.215 56.43 326.585 ;
      VIA 55.66 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 320.795 56.45 321.125 ;
      VIA 55.66 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 320.775 56.43 321.145 ;
      VIA 55.66 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 315.355 56.45 315.685 ;
      VIA 55.66 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 315.335 56.43 315.705 ;
      VIA 55.66 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 309.915 56.45 310.245 ;
      VIA 55.66 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 309.895 56.43 310.265 ;
      VIA 55.66 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 304.475 56.45 304.805 ;
      VIA 55.66 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 304.455 56.43 304.825 ;
      VIA 55.66 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 299.035 56.45 299.365 ;
      VIA 55.66 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 299.015 56.43 299.385 ;
      VIA 55.66 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 293.595 56.45 293.925 ;
      VIA 55.66 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 293.575 56.43 293.945 ;
      VIA 55.66 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 288.155 56.45 288.485 ;
      VIA 55.66 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 288.135 56.43 288.505 ;
      VIA 55.66 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 282.715 56.45 283.045 ;
      VIA 55.66 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 282.695 56.43 283.065 ;
      VIA 55.66 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 277.275 56.45 277.605 ;
      VIA 55.66 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 277.255 56.43 277.625 ;
      VIA 55.66 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 271.835 56.45 272.165 ;
      VIA 55.66 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 271.815 56.43 272.185 ;
      VIA 55.66 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 266.395 56.45 266.725 ;
      VIA 55.66 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 266.375 56.43 266.745 ;
      VIA 55.66 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 260.955 56.45 261.285 ;
      VIA 55.66 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 260.935 56.43 261.305 ;
      VIA 55.66 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 255.515 56.45 255.845 ;
      VIA 55.66 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 255.495 56.43 255.865 ;
      VIA 55.66 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 250.075 56.45 250.405 ;
      VIA 55.66 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 250.055 56.43 250.425 ;
      VIA 55.66 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 244.635 56.45 244.965 ;
      VIA 55.66 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 244.615 56.43 244.985 ;
      VIA 55.66 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 239.195 56.45 239.525 ;
      VIA 55.66 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 239.175 56.43 239.545 ;
      VIA 55.66 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 233.755 56.45 234.085 ;
      VIA 55.66 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 233.735 56.43 234.105 ;
      VIA 55.66 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 228.315 56.45 228.645 ;
      VIA 55.66 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 228.295 56.43 228.665 ;
      VIA 55.66 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 222.875 56.45 223.205 ;
      VIA 55.66 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 222.855 56.43 223.225 ;
      VIA 55.66 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 217.435 56.45 217.765 ;
      VIA 55.66 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 217.415 56.43 217.785 ;
      VIA 55.66 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 211.995 56.45 212.325 ;
      VIA 55.66 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 211.975 56.43 212.345 ;
      VIA 55.66 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 206.555 56.45 206.885 ;
      VIA 55.66 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 206.535 56.43 206.905 ;
      VIA 55.66 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 201.115 56.45 201.445 ;
      VIA 55.66 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 201.095 56.43 201.465 ;
      VIA 55.66 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 195.675 56.45 196.005 ;
      VIA 55.66 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 195.655 56.43 196.025 ;
      VIA 55.66 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 190.235 56.45 190.565 ;
      VIA 55.66 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 190.215 56.43 190.585 ;
      VIA 55.66 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 184.795 56.45 185.125 ;
      VIA 55.66 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 184.775 56.43 185.145 ;
      VIA 55.66 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 179.355 56.45 179.685 ;
      VIA 55.66 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 179.335 56.43 179.705 ;
      VIA 55.66 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 173.915 56.45 174.245 ;
      VIA 55.66 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 173.895 56.43 174.265 ;
      VIA 55.66 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 168.475 56.45 168.805 ;
      VIA 55.66 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 168.455 56.43 168.825 ;
      VIA 55.66 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 163.035 56.45 163.365 ;
      VIA 55.66 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 163.015 56.43 163.385 ;
      VIA 55.66 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 157.595 56.45 157.925 ;
      VIA 55.66 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 157.575 56.43 157.945 ;
      VIA 55.66 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 152.155 56.45 152.485 ;
      VIA 55.66 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 152.135 56.43 152.505 ;
      VIA 55.66 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 146.715 56.45 147.045 ;
      VIA 55.66 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 146.695 56.43 147.065 ;
      VIA 55.66 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 141.275 56.45 141.605 ;
      VIA 55.66 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 141.255 56.43 141.625 ;
      VIA 55.66 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 135.835 56.45 136.165 ;
      VIA 55.66 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 135.815 56.43 136.185 ;
      VIA 55.66 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 130.395 56.45 130.725 ;
      VIA 55.66 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 130.375 56.43 130.745 ;
      VIA 55.66 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 124.955 56.45 125.285 ;
      VIA 55.66 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 124.935 56.43 125.305 ;
      VIA 55.66 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 119.515 56.45 119.845 ;
      VIA 55.66 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 119.495 56.43 119.865 ;
      VIA 55.66 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 114.075 56.45 114.405 ;
      VIA 55.66 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 114.055 56.43 114.425 ;
      VIA 55.66 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 108.635 56.45 108.965 ;
      VIA 55.66 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 108.615 56.43 108.985 ;
      VIA 55.66 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 103.195 56.45 103.525 ;
      VIA 55.66 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 103.175 56.43 103.545 ;
      VIA 55.66 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 97.755 56.45 98.085 ;
      VIA 55.66 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 97.735 56.43 98.105 ;
      VIA 55.66 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 92.315 56.45 92.645 ;
      VIA 55.66 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 92.295 56.43 92.665 ;
      VIA 55.66 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 86.875 56.45 87.205 ;
      VIA 55.66 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 86.855 56.43 87.225 ;
      VIA 55.66 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 81.435 56.45 81.765 ;
      VIA 55.66 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 81.415 56.43 81.785 ;
      VIA 55.66 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 75.995 56.45 76.325 ;
      VIA 55.66 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 75.975 56.43 76.345 ;
      VIA 55.66 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 70.555 56.45 70.885 ;
      VIA 55.66 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 70.535 56.43 70.905 ;
      VIA 55.66 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 65.115 56.45 65.445 ;
      VIA 55.66 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 65.095 56.43 65.465 ;
      VIA 55.66 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 59.675 56.45 60.005 ;
      VIA 55.66 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 59.655 56.43 60.025 ;
      VIA 55.66 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 54.235 56.45 54.565 ;
      VIA 55.66 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 54.215 56.43 54.585 ;
      VIA 55.66 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 48.795 56.45 49.125 ;
      VIA 55.66 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 48.775 56.43 49.145 ;
      VIA 55.66 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 43.355 56.45 43.685 ;
      VIA 55.66 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 43.335 56.43 43.705 ;
      VIA 55.66 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 37.915 56.45 38.245 ;
      VIA 55.66 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 37.895 56.43 38.265 ;
      VIA 55.66 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 32.475 56.45 32.805 ;
      VIA 55.66 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 32.455 56.43 32.825 ;
      VIA 55.66 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 27.035 56.45 27.365 ;
      VIA 55.66 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 27.015 56.43 27.385 ;
      VIA 55.66 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 21.595 56.45 21.925 ;
      VIA 55.66 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 21.575 56.43 21.945 ;
      VIA 55.66 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 16.155 56.45 16.485 ;
      VIA 55.66 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 16.135 56.43 16.505 ;
      VIA 55.66 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 10.715 56.45 11.045 ;
      VIA 55.66 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 10.695 56.43 11.065 ;
      VIA 55.66 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 5.275 56.45 5.605 ;
      VIA 55.66 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 5.255 56.43 5.625 ;
      VIA 55.66 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 418.715 29.31 419.045 ;
      VIA 28.52 418.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 418.695 29.29 419.065 ;
      VIA 28.52 418.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 418.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 413.275 29.31 413.605 ;
      VIA 28.52 413.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 413.255 29.29 413.625 ;
      VIA 28.52 413.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 413.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 407.835 29.31 408.165 ;
      VIA 28.52 408 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 407.815 29.29 408.185 ;
      VIA 28.52 408 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 408 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 402.395 29.31 402.725 ;
      VIA 28.52 402.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 402.375 29.29 402.745 ;
      VIA 28.52 402.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 402.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 396.955 29.31 397.285 ;
      VIA 28.52 397.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 396.935 29.29 397.305 ;
      VIA 28.52 397.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 397.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 391.515 29.31 391.845 ;
      VIA 28.52 391.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 391.495 29.29 391.865 ;
      VIA 28.52 391.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 391.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 386.075 29.31 386.405 ;
      VIA 28.52 386.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 386.055 29.29 386.425 ;
      VIA 28.52 386.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 386.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 380.635 29.31 380.965 ;
      VIA 28.52 380.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 380.615 29.29 380.985 ;
      VIA 28.52 380.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 380.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 375.195 29.31 375.525 ;
      VIA 28.52 375.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 375.175 29.29 375.545 ;
      VIA 28.52 375.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 375.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 369.755 29.31 370.085 ;
      VIA 28.52 369.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 369.735 29.29 370.105 ;
      VIA 28.52 369.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 369.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 364.315 29.31 364.645 ;
      VIA 28.52 364.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 364.295 29.29 364.665 ;
      VIA 28.52 364.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 364.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 358.875 29.31 359.205 ;
      VIA 28.52 359.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 358.855 29.29 359.225 ;
      VIA 28.52 359.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 359.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 353.435 29.31 353.765 ;
      VIA 28.52 353.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 353.415 29.29 353.785 ;
      VIA 28.52 353.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 353.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 347.995 29.31 348.325 ;
      VIA 28.52 348.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 347.975 29.29 348.345 ;
      VIA 28.52 348.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 348.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 342.555 29.31 342.885 ;
      VIA 28.52 342.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 342.535 29.29 342.905 ;
      VIA 28.52 342.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 342.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 337.115 29.31 337.445 ;
      VIA 28.52 337.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 337.095 29.29 337.465 ;
      VIA 28.52 337.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 337.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 331.675 29.31 332.005 ;
      VIA 28.52 331.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 331.655 29.29 332.025 ;
      VIA 28.52 331.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 331.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 326.235 29.31 326.565 ;
      VIA 28.52 326.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 326.215 29.29 326.585 ;
      VIA 28.52 326.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 326.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 320.795 29.31 321.125 ;
      VIA 28.52 320.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 320.775 29.29 321.145 ;
      VIA 28.52 320.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 320.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 315.355 29.31 315.685 ;
      VIA 28.52 315.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 315.335 29.29 315.705 ;
      VIA 28.52 315.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 315.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 309.915 29.31 310.245 ;
      VIA 28.52 310.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 309.895 29.29 310.265 ;
      VIA 28.52 310.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 310.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 304.475 29.31 304.805 ;
      VIA 28.52 304.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 304.455 29.29 304.825 ;
      VIA 28.52 304.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 304.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 299.035 29.31 299.365 ;
      VIA 28.52 299.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 299.015 29.29 299.385 ;
      VIA 28.52 299.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 299.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 293.595 29.31 293.925 ;
      VIA 28.52 293.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 293.575 29.29 293.945 ;
      VIA 28.52 293.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 293.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 288.155 29.31 288.485 ;
      VIA 28.52 288.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 288.135 29.29 288.505 ;
      VIA 28.52 288.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 288.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 282.715 29.31 283.045 ;
      VIA 28.52 282.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 282.695 29.29 283.065 ;
      VIA 28.52 282.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 282.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 277.275 29.31 277.605 ;
      VIA 28.52 277.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 277.255 29.29 277.625 ;
      VIA 28.52 277.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 277.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 271.835 29.31 272.165 ;
      VIA 28.52 272 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 271.815 29.29 272.185 ;
      VIA 28.52 272 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 272 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 266.395 29.31 266.725 ;
      VIA 28.52 266.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 266.375 29.29 266.745 ;
      VIA 28.52 266.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 266.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 260.955 29.31 261.285 ;
      VIA 28.52 261.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 260.935 29.29 261.305 ;
      VIA 28.52 261.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 261.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 255.515 29.31 255.845 ;
      VIA 28.52 255.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 255.495 29.29 255.865 ;
      VIA 28.52 255.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 255.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 250.075 29.31 250.405 ;
      VIA 28.52 250.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 250.055 29.29 250.425 ;
      VIA 28.52 250.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 250.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 244.635 29.31 244.965 ;
      VIA 28.52 244.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 244.615 29.29 244.985 ;
      VIA 28.52 244.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 244.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 239.195 29.31 239.525 ;
      VIA 28.52 239.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 239.175 29.29 239.545 ;
      VIA 28.52 239.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 239.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 233.755 29.31 234.085 ;
      VIA 28.52 233.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 233.735 29.29 234.105 ;
      VIA 28.52 233.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 233.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 228.315 29.31 228.645 ;
      VIA 28.52 228.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 228.295 29.29 228.665 ;
      VIA 28.52 228.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 228.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 222.875 29.31 223.205 ;
      VIA 28.52 223.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 222.855 29.29 223.225 ;
      VIA 28.52 223.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 223.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 217.435 29.31 217.765 ;
      VIA 28.52 217.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 217.415 29.29 217.785 ;
      VIA 28.52 217.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 217.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 211.995 29.31 212.325 ;
      VIA 28.52 212.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 211.975 29.29 212.345 ;
      VIA 28.52 212.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 212.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 206.555 29.31 206.885 ;
      VIA 28.52 206.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 206.535 29.29 206.905 ;
      VIA 28.52 206.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 206.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 201.115 29.31 201.445 ;
      VIA 28.52 201.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 201.095 29.29 201.465 ;
      VIA 28.52 201.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 201.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 195.675 29.31 196.005 ;
      VIA 28.52 195.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 195.655 29.29 196.025 ;
      VIA 28.52 195.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 195.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 190.235 29.31 190.565 ;
      VIA 28.52 190.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 190.215 29.29 190.585 ;
      VIA 28.52 190.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 190.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 184.795 29.31 185.125 ;
      VIA 28.52 184.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 184.775 29.29 185.145 ;
      VIA 28.52 184.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 184.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 179.355 29.31 179.685 ;
      VIA 28.52 179.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 179.335 29.29 179.705 ;
      VIA 28.52 179.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 179.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 173.915 29.31 174.245 ;
      VIA 28.52 174.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 173.895 29.29 174.265 ;
      VIA 28.52 174.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 174.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 168.475 29.31 168.805 ;
      VIA 28.52 168.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 168.455 29.29 168.825 ;
      VIA 28.52 168.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 168.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 163.035 29.31 163.365 ;
      VIA 28.52 163.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 163.015 29.29 163.385 ;
      VIA 28.52 163.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 163.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 157.595 29.31 157.925 ;
      VIA 28.52 157.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 157.575 29.29 157.945 ;
      VIA 28.52 157.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 157.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 152.155 29.31 152.485 ;
      VIA 28.52 152.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 152.135 29.29 152.505 ;
      VIA 28.52 152.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 152.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 146.715 29.31 147.045 ;
      VIA 28.52 146.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 146.695 29.29 147.065 ;
      VIA 28.52 146.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 146.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 141.275 29.31 141.605 ;
      VIA 28.52 141.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 141.255 29.29 141.625 ;
      VIA 28.52 141.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 141.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 135.835 29.31 136.165 ;
      VIA 28.52 136 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 135.815 29.29 136.185 ;
      VIA 28.52 136 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 136 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 130.395 29.31 130.725 ;
      VIA 28.52 130.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 130.375 29.29 130.745 ;
      VIA 28.52 130.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 130.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 124.955 29.31 125.285 ;
      VIA 28.52 125.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 124.935 29.29 125.305 ;
      VIA 28.52 125.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 125.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 119.515 29.31 119.845 ;
      VIA 28.52 119.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 119.495 29.29 119.865 ;
      VIA 28.52 119.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 119.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 114.075 29.31 114.405 ;
      VIA 28.52 114.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 114.055 29.29 114.425 ;
      VIA 28.52 114.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 114.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 108.635 29.31 108.965 ;
      VIA 28.52 108.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 108.615 29.29 108.985 ;
      VIA 28.52 108.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 108.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 103.195 29.31 103.525 ;
      VIA 28.52 103.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 103.175 29.29 103.545 ;
      VIA 28.52 103.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 103.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 97.755 29.31 98.085 ;
      VIA 28.52 97.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 97.735 29.29 98.105 ;
      VIA 28.52 97.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 97.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 92.315 29.31 92.645 ;
      VIA 28.52 92.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 92.295 29.29 92.665 ;
      VIA 28.52 92.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 92.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 86.875 29.31 87.205 ;
      VIA 28.52 87.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 86.855 29.29 87.225 ;
      VIA 28.52 87.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 87.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 81.435 29.31 81.765 ;
      VIA 28.52 81.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 81.415 29.29 81.785 ;
      VIA 28.52 81.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 81.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 75.995 29.31 76.325 ;
      VIA 28.52 76.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 75.975 29.29 76.345 ;
      VIA 28.52 76.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 76.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 70.555 29.31 70.885 ;
      VIA 28.52 70.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 70.535 29.29 70.905 ;
      VIA 28.52 70.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 70.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 65.115 29.31 65.445 ;
      VIA 28.52 65.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 65.095 29.29 65.465 ;
      VIA 28.52 65.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 65.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 59.675 29.31 60.005 ;
      VIA 28.52 59.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 59.655 29.29 60.025 ;
      VIA 28.52 59.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 59.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 54.235 29.31 54.565 ;
      VIA 28.52 54.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 54.215 29.29 54.585 ;
      VIA 28.52 54.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 54.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 48.795 29.31 49.125 ;
      VIA 28.52 48.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 48.775 29.29 49.145 ;
      VIA 28.52 48.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 48.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 43.355 29.31 43.685 ;
      VIA 28.52 43.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 43.335 29.29 43.705 ;
      VIA 28.52 43.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 43.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 37.915 29.31 38.245 ;
      VIA 28.52 38.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 37.895 29.29 38.265 ;
      VIA 28.52 38.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 38.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 32.475 29.31 32.805 ;
      VIA 28.52 32.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 32.455 29.29 32.825 ;
      VIA 28.52 32.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 32.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 27.035 29.31 27.365 ;
      VIA 28.52 27.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 27.015 29.29 27.385 ;
      VIA 28.52 27.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 27.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 21.595 29.31 21.925 ;
      VIA 28.52 21.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 21.575 29.29 21.945 ;
      VIA 28.52 21.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 21.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 16.155 29.31 16.485 ;
      VIA 28.52 16.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 16.135 29.29 16.505 ;
      VIA 28.52 16.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 16.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 10.715 29.31 11.045 ;
      VIA 28.52 10.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 10.695 29.29 11.065 ;
      VIA 28.52 10.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 10.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 5.275 29.31 5.605 ;
      VIA 28.52 5.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 5.255 29.29 5.625 ;
      VIA 28.52 5.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 5.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  14.15 396.32 395.71 397.92 ;
        RECT  14.15 369.12 395.71 370.72 ;
        RECT  14.15 341.92 395.71 343.52 ;
        RECT  14.15 314.72 395.71 316.32 ;
        RECT  14.15 287.52 395.71 289.12 ;
        RECT  14.15 260.32 395.71 261.92 ;
        RECT  14.15 233.12 395.71 234.72 ;
        RECT  14.15 205.92 395.71 207.52 ;
        RECT  14.15 178.72 395.71 180.32 ;
        RECT  14.15 151.52 395.71 153.12 ;
        RECT  14.15 124.32 395.71 125.92 ;
        RECT  14.15 97.12 395.71 98.72 ;
        RECT  14.15 69.92 395.71 71.52 ;
        RECT  14.15 42.72 395.71 44.32 ;
        RECT  14.15 15.52 395.71 17.12 ;
      LAYER met4 ;
        RECT  394.11 2.48 395.71 416.4 ;
        RECT  366.97 2.48 368.57 416.4 ;
        RECT  339.83 2.48 341.43 416.4 ;
        RECT  312.69 2.48 314.29 416.4 ;
        RECT  285.55 2.48 287.15 416.4 ;
        RECT  258.41 2.48 260.01 416.4 ;
        RECT  231.27 2.48 232.87 416.4 ;
        RECT  204.13 2.48 205.73 416.4 ;
        RECT  176.99 2.48 178.59 416.4 ;
        RECT  149.85 2.48 151.45 416.4 ;
        RECT  122.71 2.48 124.31 416.4 ;
        RECT  95.57 2.48 97.17 416.4 ;
        RECT  68.43 2.48 70.03 416.4 ;
        RECT  41.29 2.48 42.89 416.4 ;
        RECT  14.15 2.48 15.75 416.4 ;
      LAYER met1 ;
        RECT  1.38 415.92 420.9 416.4 ;
        RECT  1.38 410.48 420.9 410.96 ;
        RECT  1.38 405.04 420.9 405.52 ;
        RECT  1.38 399.6 420.9 400.08 ;
        RECT  1.38 394.16 420.9 394.64 ;
        RECT  1.38 388.72 420.9 389.2 ;
        RECT  1.38 383.28 420.9 383.76 ;
        RECT  1.38 377.84 420.9 378.32 ;
        RECT  1.38 372.4 420.9 372.88 ;
        RECT  1.38 366.96 420.9 367.44 ;
        RECT  1.38 361.52 420.9 362 ;
        RECT  1.38 356.08 420.9 356.56 ;
        RECT  1.38 350.64 420.9 351.12 ;
        RECT  1.38 345.2 420.9 345.68 ;
        RECT  1.38 339.76 420.9 340.24 ;
        RECT  1.38 334.32 420.9 334.8 ;
        RECT  1.38 328.88 420.9 329.36 ;
        RECT  1.38 323.44 420.9 323.92 ;
        RECT  1.38 318 420.9 318.48 ;
        RECT  1.38 312.56 420.9 313.04 ;
        RECT  1.38 307.12 420.9 307.6 ;
        RECT  1.38 301.68 420.9 302.16 ;
        RECT  1.38 296.24 420.9 296.72 ;
        RECT  1.38 290.8 420.9 291.28 ;
        RECT  1.38 285.36 420.9 285.84 ;
        RECT  1.38 279.92 420.9 280.4 ;
        RECT  1.38 274.48 420.9 274.96 ;
        RECT  1.38 269.04 420.9 269.52 ;
        RECT  1.38 263.6 420.9 264.08 ;
        RECT  1.38 258.16 420.9 258.64 ;
        RECT  1.38 252.72 420.9 253.2 ;
        RECT  1.38 247.28 420.9 247.76 ;
        RECT  1.38 241.84 420.9 242.32 ;
        RECT  1.38 236.4 420.9 236.88 ;
        RECT  1.38 230.96 420.9 231.44 ;
        RECT  1.38 225.52 420.9 226 ;
        RECT  1.38 220.08 420.9 220.56 ;
        RECT  1.38 214.64 420.9 215.12 ;
        RECT  1.38 209.2 420.9 209.68 ;
        RECT  1.38 203.76 420.9 204.24 ;
        RECT  1.38 198.32 420.9 198.8 ;
        RECT  1.38 192.88 420.9 193.36 ;
        RECT  1.38 187.44 420.9 187.92 ;
        RECT  1.38 182 420.9 182.48 ;
        RECT  1.38 176.56 420.9 177.04 ;
        RECT  1.38 171.12 420.9 171.6 ;
        RECT  1.38 165.68 420.9 166.16 ;
        RECT  1.38 160.24 420.9 160.72 ;
        RECT  1.38 154.8 420.9 155.28 ;
        RECT  1.38 149.36 420.9 149.84 ;
        RECT  1.38 143.92 420.9 144.4 ;
        RECT  1.38 138.48 420.9 138.96 ;
        RECT  1.38 133.04 420.9 133.52 ;
        RECT  1.38 127.6 420.9 128.08 ;
        RECT  1.38 122.16 420.9 122.64 ;
        RECT  1.38 116.72 420.9 117.2 ;
        RECT  1.38 111.28 420.9 111.76 ;
        RECT  1.38 105.84 420.9 106.32 ;
        RECT  1.38 100.4 420.9 100.88 ;
        RECT  1.38 94.96 420.9 95.44 ;
        RECT  1.38 89.52 420.9 90 ;
        RECT  1.38 84.08 420.9 84.56 ;
        RECT  1.38 78.64 420.9 79.12 ;
        RECT  1.38 73.2 420.9 73.68 ;
        RECT  1.38 67.76 420.9 68.24 ;
        RECT  1.38 62.32 420.9 62.8 ;
        RECT  1.38 56.88 420.9 57.36 ;
        RECT  1.38 51.44 420.9 51.92 ;
        RECT  1.38 46 420.9 46.48 ;
        RECT  1.38 40.56 420.9 41.04 ;
        RECT  1.38 35.12 420.9 35.6 ;
        RECT  1.38 29.68 420.9 30.16 ;
        RECT  1.38 24.24 420.9 24.72 ;
        RECT  1.38 18.8 420.9 19.28 ;
        RECT  1.38 13.36 420.9 13.84 ;
        RECT  1.38 7.92 420.9 8.4 ;
        RECT  1.38 2.48 420.9 2.96 ;
      VIA 394.91 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 394.91 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 367.77 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 340.63 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 313.49 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 397.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 369.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 342.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 315.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 288.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 261.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 233.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 206.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 179.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 152.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 125.12 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 97.92 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 70.72 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 43.52 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 16.32 ibex_register_file_ff_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  394.12 415.995 395.7 416.325 ;
      VIA 394.91 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 415.975 395.68 416.345 ;
      VIA 394.91 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 410.555 395.7 410.885 ;
      VIA 394.91 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 410.535 395.68 410.905 ;
      VIA 394.91 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 405.115 395.7 405.445 ;
      VIA 394.91 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 405.095 395.68 405.465 ;
      VIA 394.91 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 399.675 395.7 400.005 ;
      VIA 394.91 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 399.655 395.68 400.025 ;
      VIA 394.91 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 394.235 395.7 394.565 ;
      VIA 394.91 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 394.215 395.68 394.585 ;
      VIA 394.91 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 388.795 395.7 389.125 ;
      VIA 394.91 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 388.775 395.68 389.145 ;
      VIA 394.91 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 383.355 395.7 383.685 ;
      VIA 394.91 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 383.335 395.68 383.705 ;
      VIA 394.91 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 377.915 395.7 378.245 ;
      VIA 394.91 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 377.895 395.68 378.265 ;
      VIA 394.91 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 372.475 395.7 372.805 ;
      VIA 394.91 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 372.455 395.68 372.825 ;
      VIA 394.91 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 367.035 395.7 367.365 ;
      VIA 394.91 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 367.015 395.68 367.385 ;
      VIA 394.91 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 361.595 395.7 361.925 ;
      VIA 394.91 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 361.575 395.68 361.945 ;
      VIA 394.91 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 356.155 395.7 356.485 ;
      VIA 394.91 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 356.135 395.68 356.505 ;
      VIA 394.91 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 350.715 395.7 351.045 ;
      VIA 394.91 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 350.695 395.68 351.065 ;
      VIA 394.91 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 345.275 395.7 345.605 ;
      VIA 394.91 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 345.255 395.68 345.625 ;
      VIA 394.91 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 339.835 395.7 340.165 ;
      VIA 394.91 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 339.815 395.68 340.185 ;
      VIA 394.91 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 334.395 395.7 334.725 ;
      VIA 394.91 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 334.375 395.68 334.745 ;
      VIA 394.91 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 328.955 395.7 329.285 ;
      VIA 394.91 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 328.935 395.68 329.305 ;
      VIA 394.91 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 323.515 395.7 323.845 ;
      VIA 394.91 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 323.495 395.68 323.865 ;
      VIA 394.91 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 318.075 395.7 318.405 ;
      VIA 394.91 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 318.055 395.68 318.425 ;
      VIA 394.91 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 312.635 395.7 312.965 ;
      VIA 394.91 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 312.615 395.68 312.985 ;
      VIA 394.91 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 307.195 395.7 307.525 ;
      VIA 394.91 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 307.175 395.68 307.545 ;
      VIA 394.91 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 301.755 395.7 302.085 ;
      VIA 394.91 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 301.735 395.68 302.105 ;
      VIA 394.91 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 296.315 395.7 296.645 ;
      VIA 394.91 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 296.295 395.68 296.665 ;
      VIA 394.91 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 290.875 395.7 291.205 ;
      VIA 394.91 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 290.855 395.68 291.225 ;
      VIA 394.91 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 285.435 395.7 285.765 ;
      VIA 394.91 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 285.415 395.68 285.785 ;
      VIA 394.91 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 279.995 395.7 280.325 ;
      VIA 394.91 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 279.975 395.68 280.345 ;
      VIA 394.91 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 274.555 395.7 274.885 ;
      VIA 394.91 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 274.535 395.68 274.905 ;
      VIA 394.91 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 269.115 395.7 269.445 ;
      VIA 394.91 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 269.095 395.68 269.465 ;
      VIA 394.91 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 263.675 395.7 264.005 ;
      VIA 394.91 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 263.655 395.68 264.025 ;
      VIA 394.91 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 258.235 395.7 258.565 ;
      VIA 394.91 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 258.215 395.68 258.585 ;
      VIA 394.91 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 252.795 395.7 253.125 ;
      VIA 394.91 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 252.775 395.68 253.145 ;
      VIA 394.91 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 247.355 395.7 247.685 ;
      VIA 394.91 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 247.335 395.68 247.705 ;
      VIA 394.91 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 241.915 395.7 242.245 ;
      VIA 394.91 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 241.895 395.68 242.265 ;
      VIA 394.91 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 236.475 395.7 236.805 ;
      VIA 394.91 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 236.455 395.68 236.825 ;
      VIA 394.91 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 231.035 395.7 231.365 ;
      VIA 394.91 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 231.015 395.68 231.385 ;
      VIA 394.91 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 225.595 395.7 225.925 ;
      VIA 394.91 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 225.575 395.68 225.945 ;
      VIA 394.91 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 220.155 395.7 220.485 ;
      VIA 394.91 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 220.135 395.68 220.505 ;
      VIA 394.91 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 214.715 395.7 215.045 ;
      VIA 394.91 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 214.695 395.68 215.065 ;
      VIA 394.91 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 209.275 395.7 209.605 ;
      VIA 394.91 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 209.255 395.68 209.625 ;
      VIA 394.91 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 203.835 395.7 204.165 ;
      VIA 394.91 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 203.815 395.68 204.185 ;
      VIA 394.91 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 198.395 395.7 198.725 ;
      VIA 394.91 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 198.375 395.68 198.745 ;
      VIA 394.91 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 192.955 395.7 193.285 ;
      VIA 394.91 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 192.935 395.68 193.305 ;
      VIA 394.91 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 187.515 395.7 187.845 ;
      VIA 394.91 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 187.495 395.68 187.865 ;
      VIA 394.91 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 182.075 395.7 182.405 ;
      VIA 394.91 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 182.055 395.68 182.425 ;
      VIA 394.91 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 176.635 395.7 176.965 ;
      VIA 394.91 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 176.615 395.68 176.985 ;
      VIA 394.91 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 171.195 395.7 171.525 ;
      VIA 394.91 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 171.175 395.68 171.545 ;
      VIA 394.91 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 165.755 395.7 166.085 ;
      VIA 394.91 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 165.735 395.68 166.105 ;
      VIA 394.91 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 160.315 395.7 160.645 ;
      VIA 394.91 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 160.295 395.68 160.665 ;
      VIA 394.91 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 154.875 395.7 155.205 ;
      VIA 394.91 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 154.855 395.68 155.225 ;
      VIA 394.91 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 149.435 395.7 149.765 ;
      VIA 394.91 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 149.415 395.68 149.785 ;
      VIA 394.91 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 143.995 395.7 144.325 ;
      VIA 394.91 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 143.975 395.68 144.345 ;
      VIA 394.91 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 138.555 395.7 138.885 ;
      VIA 394.91 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 138.535 395.68 138.905 ;
      VIA 394.91 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 133.115 395.7 133.445 ;
      VIA 394.91 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 133.095 395.68 133.465 ;
      VIA 394.91 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 127.675 395.7 128.005 ;
      VIA 394.91 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 127.655 395.68 128.025 ;
      VIA 394.91 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 122.235 395.7 122.565 ;
      VIA 394.91 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 122.215 395.68 122.585 ;
      VIA 394.91 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 116.795 395.7 117.125 ;
      VIA 394.91 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 116.775 395.68 117.145 ;
      VIA 394.91 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 111.355 395.7 111.685 ;
      VIA 394.91 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 111.335 395.68 111.705 ;
      VIA 394.91 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 105.915 395.7 106.245 ;
      VIA 394.91 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 105.895 395.68 106.265 ;
      VIA 394.91 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 100.475 395.7 100.805 ;
      VIA 394.91 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 100.455 395.68 100.825 ;
      VIA 394.91 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 95.035 395.7 95.365 ;
      VIA 394.91 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 95.015 395.68 95.385 ;
      VIA 394.91 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 89.595 395.7 89.925 ;
      VIA 394.91 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 89.575 395.68 89.945 ;
      VIA 394.91 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 84.155 395.7 84.485 ;
      VIA 394.91 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 84.135 395.68 84.505 ;
      VIA 394.91 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 78.715 395.7 79.045 ;
      VIA 394.91 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 78.695 395.68 79.065 ;
      VIA 394.91 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 73.275 395.7 73.605 ;
      VIA 394.91 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 73.255 395.68 73.625 ;
      VIA 394.91 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 67.835 395.7 68.165 ;
      VIA 394.91 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 67.815 395.68 68.185 ;
      VIA 394.91 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 62.395 395.7 62.725 ;
      VIA 394.91 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 62.375 395.68 62.745 ;
      VIA 394.91 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 56.955 395.7 57.285 ;
      VIA 394.91 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 56.935 395.68 57.305 ;
      VIA 394.91 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 51.515 395.7 51.845 ;
      VIA 394.91 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 51.495 395.68 51.865 ;
      VIA 394.91 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 46.075 395.7 46.405 ;
      VIA 394.91 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 46.055 395.68 46.425 ;
      VIA 394.91 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 40.635 395.7 40.965 ;
      VIA 394.91 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 40.615 395.68 40.985 ;
      VIA 394.91 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 35.195 395.7 35.525 ;
      VIA 394.91 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 35.175 395.68 35.545 ;
      VIA 394.91 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 29.755 395.7 30.085 ;
      VIA 394.91 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 29.735 395.68 30.105 ;
      VIA 394.91 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 24.315 395.7 24.645 ;
      VIA 394.91 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 24.295 395.68 24.665 ;
      VIA 394.91 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 18.875 395.7 19.205 ;
      VIA 394.91 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 18.855 395.68 19.225 ;
      VIA 394.91 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 13.435 395.7 13.765 ;
      VIA 394.91 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 13.415 395.68 13.785 ;
      VIA 394.91 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 7.995 395.7 8.325 ;
      VIA 394.91 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 7.975 395.68 8.345 ;
      VIA 394.91 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  394.12 2.555 395.7 2.885 ;
      VIA 394.91 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  394.14 2.535 395.68 2.905 ;
      VIA 394.91 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 394.91 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 415.995 368.56 416.325 ;
      VIA 367.77 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 415.975 368.54 416.345 ;
      VIA 367.77 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 410.555 368.56 410.885 ;
      VIA 367.77 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 410.535 368.54 410.905 ;
      VIA 367.77 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 405.115 368.56 405.445 ;
      VIA 367.77 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 405.095 368.54 405.465 ;
      VIA 367.77 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 399.675 368.56 400.005 ;
      VIA 367.77 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 399.655 368.54 400.025 ;
      VIA 367.77 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 394.235 368.56 394.565 ;
      VIA 367.77 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 394.215 368.54 394.585 ;
      VIA 367.77 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 388.795 368.56 389.125 ;
      VIA 367.77 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 388.775 368.54 389.145 ;
      VIA 367.77 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 383.355 368.56 383.685 ;
      VIA 367.77 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 383.335 368.54 383.705 ;
      VIA 367.77 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 377.915 368.56 378.245 ;
      VIA 367.77 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 377.895 368.54 378.265 ;
      VIA 367.77 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 372.475 368.56 372.805 ;
      VIA 367.77 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 372.455 368.54 372.825 ;
      VIA 367.77 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 367.035 368.56 367.365 ;
      VIA 367.77 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 367.015 368.54 367.385 ;
      VIA 367.77 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 361.595 368.56 361.925 ;
      VIA 367.77 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 361.575 368.54 361.945 ;
      VIA 367.77 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 356.155 368.56 356.485 ;
      VIA 367.77 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 356.135 368.54 356.505 ;
      VIA 367.77 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 350.715 368.56 351.045 ;
      VIA 367.77 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 350.695 368.54 351.065 ;
      VIA 367.77 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 345.275 368.56 345.605 ;
      VIA 367.77 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 345.255 368.54 345.625 ;
      VIA 367.77 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 339.835 368.56 340.165 ;
      VIA 367.77 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 339.815 368.54 340.185 ;
      VIA 367.77 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 334.395 368.56 334.725 ;
      VIA 367.77 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 334.375 368.54 334.745 ;
      VIA 367.77 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 328.955 368.56 329.285 ;
      VIA 367.77 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 328.935 368.54 329.305 ;
      VIA 367.77 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 323.515 368.56 323.845 ;
      VIA 367.77 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 323.495 368.54 323.865 ;
      VIA 367.77 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 318.075 368.56 318.405 ;
      VIA 367.77 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 318.055 368.54 318.425 ;
      VIA 367.77 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 312.635 368.56 312.965 ;
      VIA 367.77 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 312.615 368.54 312.985 ;
      VIA 367.77 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 307.195 368.56 307.525 ;
      VIA 367.77 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 307.175 368.54 307.545 ;
      VIA 367.77 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 301.755 368.56 302.085 ;
      VIA 367.77 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 301.735 368.54 302.105 ;
      VIA 367.77 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 296.315 368.56 296.645 ;
      VIA 367.77 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 296.295 368.54 296.665 ;
      VIA 367.77 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 290.875 368.56 291.205 ;
      VIA 367.77 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 290.855 368.54 291.225 ;
      VIA 367.77 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 285.435 368.56 285.765 ;
      VIA 367.77 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 285.415 368.54 285.785 ;
      VIA 367.77 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 279.995 368.56 280.325 ;
      VIA 367.77 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 279.975 368.54 280.345 ;
      VIA 367.77 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 274.555 368.56 274.885 ;
      VIA 367.77 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 274.535 368.54 274.905 ;
      VIA 367.77 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 269.115 368.56 269.445 ;
      VIA 367.77 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 269.095 368.54 269.465 ;
      VIA 367.77 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 263.675 368.56 264.005 ;
      VIA 367.77 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 263.655 368.54 264.025 ;
      VIA 367.77 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 258.235 368.56 258.565 ;
      VIA 367.77 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 258.215 368.54 258.585 ;
      VIA 367.77 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 252.795 368.56 253.125 ;
      VIA 367.77 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 252.775 368.54 253.145 ;
      VIA 367.77 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 247.355 368.56 247.685 ;
      VIA 367.77 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 247.335 368.54 247.705 ;
      VIA 367.77 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 241.915 368.56 242.245 ;
      VIA 367.77 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 241.895 368.54 242.265 ;
      VIA 367.77 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 236.475 368.56 236.805 ;
      VIA 367.77 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 236.455 368.54 236.825 ;
      VIA 367.77 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 231.035 368.56 231.365 ;
      VIA 367.77 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 231.015 368.54 231.385 ;
      VIA 367.77 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 225.595 368.56 225.925 ;
      VIA 367.77 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 225.575 368.54 225.945 ;
      VIA 367.77 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 220.155 368.56 220.485 ;
      VIA 367.77 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 220.135 368.54 220.505 ;
      VIA 367.77 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 214.715 368.56 215.045 ;
      VIA 367.77 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 214.695 368.54 215.065 ;
      VIA 367.77 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 209.275 368.56 209.605 ;
      VIA 367.77 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 209.255 368.54 209.625 ;
      VIA 367.77 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 203.835 368.56 204.165 ;
      VIA 367.77 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 203.815 368.54 204.185 ;
      VIA 367.77 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 198.395 368.56 198.725 ;
      VIA 367.77 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 198.375 368.54 198.745 ;
      VIA 367.77 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 192.955 368.56 193.285 ;
      VIA 367.77 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 192.935 368.54 193.305 ;
      VIA 367.77 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 187.515 368.56 187.845 ;
      VIA 367.77 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 187.495 368.54 187.865 ;
      VIA 367.77 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 182.075 368.56 182.405 ;
      VIA 367.77 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 182.055 368.54 182.425 ;
      VIA 367.77 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 176.635 368.56 176.965 ;
      VIA 367.77 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 176.615 368.54 176.985 ;
      VIA 367.77 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 171.195 368.56 171.525 ;
      VIA 367.77 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 171.175 368.54 171.545 ;
      VIA 367.77 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 165.755 368.56 166.085 ;
      VIA 367.77 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 165.735 368.54 166.105 ;
      VIA 367.77 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 160.315 368.56 160.645 ;
      VIA 367.77 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 160.295 368.54 160.665 ;
      VIA 367.77 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 154.875 368.56 155.205 ;
      VIA 367.77 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 154.855 368.54 155.225 ;
      VIA 367.77 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 149.435 368.56 149.765 ;
      VIA 367.77 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 149.415 368.54 149.785 ;
      VIA 367.77 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 143.995 368.56 144.325 ;
      VIA 367.77 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 143.975 368.54 144.345 ;
      VIA 367.77 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 138.555 368.56 138.885 ;
      VIA 367.77 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 138.535 368.54 138.905 ;
      VIA 367.77 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 133.115 368.56 133.445 ;
      VIA 367.77 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 133.095 368.54 133.465 ;
      VIA 367.77 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 127.675 368.56 128.005 ;
      VIA 367.77 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 127.655 368.54 128.025 ;
      VIA 367.77 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 122.235 368.56 122.565 ;
      VIA 367.77 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 122.215 368.54 122.585 ;
      VIA 367.77 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 116.795 368.56 117.125 ;
      VIA 367.77 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 116.775 368.54 117.145 ;
      VIA 367.77 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 111.355 368.56 111.685 ;
      VIA 367.77 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 111.335 368.54 111.705 ;
      VIA 367.77 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 105.915 368.56 106.245 ;
      VIA 367.77 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 105.895 368.54 106.265 ;
      VIA 367.77 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 100.475 368.56 100.805 ;
      VIA 367.77 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 100.455 368.54 100.825 ;
      VIA 367.77 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 95.035 368.56 95.365 ;
      VIA 367.77 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 95.015 368.54 95.385 ;
      VIA 367.77 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 89.595 368.56 89.925 ;
      VIA 367.77 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 89.575 368.54 89.945 ;
      VIA 367.77 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 84.155 368.56 84.485 ;
      VIA 367.77 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 84.135 368.54 84.505 ;
      VIA 367.77 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 78.715 368.56 79.045 ;
      VIA 367.77 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 78.695 368.54 79.065 ;
      VIA 367.77 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 73.275 368.56 73.605 ;
      VIA 367.77 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 73.255 368.54 73.625 ;
      VIA 367.77 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 67.835 368.56 68.165 ;
      VIA 367.77 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 67.815 368.54 68.185 ;
      VIA 367.77 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 62.395 368.56 62.725 ;
      VIA 367.77 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 62.375 368.54 62.745 ;
      VIA 367.77 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 56.955 368.56 57.285 ;
      VIA 367.77 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 56.935 368.54 57.305 ;
      VIA 367.77 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 51.515 368.56 51.845 ;
      VIA 367.77 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 51.495 368.54 51.865 ;
      VIA 367.77 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 46.075 368.56 46.405 ;
      VIA 367.77 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 46.055 368.54 46.425 ;
      VIA 367.77 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 40.635 368.56 40.965 ;
      VIA 367.77 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 40.615 368.54 40.985 ;
      VIA 367.77 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 35.195 368.56 35.525 ;
      VIA 367.77 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 35.175 368.54 35.545 ;
      VIA 367.77 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 29.755 368.56 30.085 ;
      VIA 367.77 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 29.735 368.54 30.105 ;
      VIA 367.77 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 24.315 368.56 24.645 ;
      VIA 367.77 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 24.295 368.54 24.665 ;
      VIA 367.77 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 18.875 368.56 19.205 ;
      VIA 367.77 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 18.855 368.54 19.225 ;
      VIA 367.77 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 13.435 368.56 13.765 ;
      VIA 367.77 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 13.415 368.54 13.785 ;
      VIA 367.77 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 7.995 368.56 8.325 ;
      VIA 367.77 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 7.975 368.54 8.345 ;
      VIA 367.77 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  366.98 2.555 368.56 2.885 ;
      VIA 367.77 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  367 2.535 368.54 2.905 ;
      VIA 367.77 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 367.77 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 415.995 341.42 416.325 ;
      VIA 340.63 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 415.975 341.4 416.345 ;
      VIA 340.63 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 410.555 341.42 410.885 ;
      VIA 340.63 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 410.535 341.4 410.905 ;
      VIA 340.63 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 405.115 341.42 405.445 ;
      VIA 340.63 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 405.095 341.4 405.465 ;
      VIA 340.63 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 399.675 341.42 400.005 ;
      VIA 340.63 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 399.655 341.4 400.025 ;
      VIA 340.63 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 394.235 341.42 394.565 ;
      VIA 340.63 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 394.215 341.4 394.585 ;
      VIA 340.63 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 388.795 341.42 389.125 ;
      VIA 340.63 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 388.775 341.4 389.145 ;
      VIA 340.63 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 383.355 341.42 383.685 ;
      VIA 340.63 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 383.335 341.4 383.705 ;
      VIA 340.63 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 377.915 341.42 378.245 ;
      VIA 340.63 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 377.895 341.4 378.265 ;
      VIA 340.63 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 372.475 341.42 372.805 ;
      VIA 340.63 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 372.455 341.4 372.825 ;
      VIA 340.63 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 367.035 341.42 367.365 ;
      VIA 340.63 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 367.015 341.4 367.385 ;
      VIA 340.63 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 361.595 341.42 361.925 ;
      VIA 340.63 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 361.575 341.4 361.945 ;
      VIA 340.63 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 356.155 341.42 356.485 ;
      VIA 340.63 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 356.135 341.4 356.505 ;
      VIA 340.63 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 350.715 341.42 351.045 ;
      VIA 340.63 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 350.695 341.4 351.065 ;
      VIA 340.63 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 345.275 341.42 345.605 ;
      VIA 340.63 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 345.255 341.4 345.625 ;
      VIA 340.63 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 339.835 341.42 340.165 ;
      VIA 340.63 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 339.815 341.4 340.185 ;
      VIA 340.63 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 334.395 341.42 334.725 ;
      VIA 340.63 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 334.375 341.4 334.745 ;
      VIA 340.63 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 328.955 341.42 329.285 ;
      VIA 340.63 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 328.935 341.4 329.305 ;
      VIA 340.63 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 323.515 341.42 323.845 ;
      VIA 340.63 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 323.495 341.4 323.865 ;
      VIA 340.63 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 318.075 341.42 318.405 ;
      VIA 340.63 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 318.055 341.4 318.425 ;
      VIA 340.63 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 312.635 341.42 312.965 ;
      VIA 340.63 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 312.615 341.4 312.985 ;
      VIA 340.63 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 307.195 341.42 307.525 ;
      VIA 340.63 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 307.175 341.4 307.545 ;
      VIA 340.63 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 301.755 341.42 302.085 ;
      VIA 340.63 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 301.735 341.4 302.105 ;
      VIA 340.63 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 296.315 341.42 296.645 ;
      VIA 340.63 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 296.295 341.4 296.665 ;
      VIA 340.63 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 290.875 341.42 291.205 ;
      VIA 340.63 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 290.855 341.4 291.225 ;
      VIA 340.63 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 285.435 341.42 285.765 ;
      VIA 340.63 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 285.415 341.4 285.785 ;
      VIA 340.63 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 279.995 341.42 280.325 ;
      VIA 340.63 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 279.975 341.4 280.345 ;
      VIA 340.63 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 274.555 341.42 274.885 ;
      VIA 340.63 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 274.535 341.4 274.905 ;
      VIA 340.63 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 269.115 341.42 269.445 ;
      VIA 340.63 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 269.095 341.4 269.465 ;
      VIA 340.63 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 263.675 341.42 264.005 ;
      VIA 340.63 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 263.655 341.4 264.025 ;
      VIA 340.63 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 258.235 341.42 258.565 ;
      VIA 340.63 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 258.215 341.4 258.585 ;
      VIA 340.63 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 252.795 341.42 253.125 ;
      VIA 340.63 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 252.775 341.4 253.145 ;
      VIA 340.63 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 247.355 341.42 247.685 ;
      VIA 340.63 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 247.335 341.4 247.705 ;
      VIA 340.63 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 241.915 341.42 242.245 ;
      VIA 340.63 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 241.895 341.4 242.265 ;
      VIA 340.63 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 236.475 341.42 236.805 ;
      VIA 340.63 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 236.455 341.4 236.825 ;
      VIA 340.63 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 231.035 341.42 231.365 ;
      VIA 340.63 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 231.015 341.4 231.385 ;
      VIA 340.63 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 225.595 341.42 225.925 ;
      VIA 340.63 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 225.575 341.4 225.945 ;
      VIA 340.63 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 220.155 341.42 220.485 ;
      VIA 340.63 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 220.135 341.4 220.505 ;
      VIA 340.63 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 214.715 341.42 215.045 ;
      VIA 340.63 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 214.695 341.4 215.065 ;
      VIA 340.63 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 209.275 341.42 209.605 ;
      VIA 340.63 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 209.255 341.4 209.625 ;
      VIA 340.63 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 203.835 341.42 204.165 ;
      VIA 340.63 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 203.815 341.4 204.185 ;
      VIA 340.63 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 198.395 341.42 198.725 ;
      VIA 340.63 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 198.375 341.4 198.745 ;
      VIA 340.63 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 192.955 341.42 193.285 ;
      VIA 340.63 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 192.935 341.4 193.305 ;
      VIA 340.63 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 187.515 341.42 187.845 ;
      VIA 340.63 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 187.495 341.4 187.865 ;
      VIA 340.63 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 182.075 341.42 182.405 ;
      VIA 340.63 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 182.055 341.4 182.425 ;
      VIA 340.63 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 176.635 341.42 176.965 ;
      VIA 340.63 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 176.615 341.4 176.985 ;
      VIA 340.63 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 171.195 341.42 171.525 ;
      VIA 340.63 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 171.175 341.4 171.545 ;
      VIA 340.63 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 165.755 341.42 166.085 ;
      VIA 340.63 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 165.735 341.4 166.105 ;
      VIA 340.63 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 160.315 341.42 160.645 ;
      VIA 340.63 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 160.295 341.4 160.665 ;
      VIA 340.63 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 154.875 341.42 155.205 ;
      VIA 340.63 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 154.855 341.4 155.225 ;
      VIA 340.63 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 149.435 341.42 149.765 ;
      VIA 340.63 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 149.415 341.4 149.785 ;
      VIA 340.63 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 143.995 341.42 144.325 ;
      VIA 340.63 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 143.975 341.4 144.345 ;
      VIA 340.63 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 138.555 341.42 138.885 ;
      VIA 340.63 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 138.535 341.4 138.905 ;
      VIA 340.63 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 133.115 341.42 133.445 ;
      VIA 340.63 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 133.095 341.4 133.465 ;
      VIA 340.63 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 127.675 341.42 128.005 ;
      VIA 340.63 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 127.655 341.4 128.025 ;
      VIA 340.63 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 122.235 341.42 122.565 ;
      VIA 340.63 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 122.215 341.4 122.585 ;
      VIA 340.63 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 116.795 341.42 117.125 ;
      VIA 340.63 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 116.775 341.4 117.145 ;
      VIA 340.63 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 111.355 341.42 111.685 ;
      VIA 340.63 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 111.335 341.4 111.705 ;
      VIA 340.63 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 105.915 341.42 106.245 ;
      VIA 340.63 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 105.895 341.4 106.265 ;
      VIA 340.63 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 100.475 341.42 100.805 ;
      VIA 340.63 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 100.455 341.4 100.825 ;
      VIA 340.63 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 95.035 341.42 95.365 ;
      VIA 340.63 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 95.015 341.4 95.385 ;
      VIA 340.63 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 89.595 341.42 89.925 ;
      VIA 340.63 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 89.575 341.4 89.945 ;
      VIA 340.63 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 84.155 341.42 84.485 ;
      VIA 340.63 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 84.135 341.4 84.505 ;
      VIA 340.63 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 78.715 341.42 79.045 ;
      VIA 340.63 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 78.695 341.4 79.065 ;
      VIA 340.63 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 73.275 341.42 73.605 ;
      VIA 340.63 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 73.255 341.4 73.625 ;
      VIA 340.63 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 67.835 341.42 68.165 ;
      VIA 340.63 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 67.815 341.4 68.185 ;
      VIA 340.63 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 62.395 341.42 62.725 ;
      VIA 340.63 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 62.375 341.4 62.745 ;
      VIA 340.63 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 56.955 341.42 57.285 ;
      VIA 340.63 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 56.935 341.4 57.305 ;
      VIA 340.63 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 51.515 341.42 51.845 ;
      VIA 340.63 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 51.495 341.4 51.865 ;
      VIA 340.63 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 46.075 341.42 46.405 ;
      VIA 340.63 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 46.055 341.4 46.425 ;
      VIA 340.63 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 40.635 341.42 40.965 ;
      VIA 340.63 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 40.615 341.4 40.985 ;
      VIA 340.63 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 35.195 341.42 35.525 ;
      VIA 340.63 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 35.175 341.4 35.545 ;
      VIA 340.63 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 29.755 341.42 30.085 ;
      VIA 340.63 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 29.735 341.4 30.105 ;
      VIA 340.63 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 24.315 341.42 24.645 ;
      VIA 340.63 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 24.295 341.4 24.665 ;
      VIA 340.63 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 18.875 341.42 19.205 ;
      VIA 340.63 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 18.855 341.4 19.225 ;
      VIA 340.63 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 13.435 341.42 13.765 ;
      VIA 340.63 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 13.415 341.4 13.785 ;
      VIA 340.63 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 7.995 341.42 8.325 ;
      VIA 340.63 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 7.975 341.4 8.345 ;
      VIA 340.63 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  339.84 2.555 341.42 2.885 ;
      VIA 340.63 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  339.86 2.535 341.4 2.905 ;
      VIA 340.63 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 340.63 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 415.995 314.28 416.325 ;
      VIA 313.49 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 415.975 314.26 416.345 ;
      VIA 313.49 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 410.555 314.28 410.885 ;
      VIA 313.49 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 410.535 314.26 410.905 ;
      VIA 313.49 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 405.115 314.28 405.445 ;
      VIA 313.49 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 405.095 314.26 405.465 ;
      VIA 313.49 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 399.675 314.28 400.005 ;
      VIA 313.49 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 399.655 314.26 400.025 ;
      VIA 313.49 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 394.235 314.28 394.565 ;
      VIA 313.49 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 394.215 314.26 394.585 ;
      VIA 313.49 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 388.795 314.28 389.125 ;
      VIA 313.49 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 388.775 314.26 389.145 ;
      VIA 313.49 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 383.355 314.28 383.685 ;
      VIA 313.49 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 383.335 314.26 383.705 ;
      VIA 313.49 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 377.915 314.28 378.245 ;
      VIA 313.49 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 377.895 314.26 378.265 ;
      VIA 313.49 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 372.475 314.28 372.805 ;
      VIA 313.49 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 372.455 314.26 372.825 ;
      VIA 313.49 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 367.035 314.28 367.365 ;
      VIA 313.49 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 367.015 314.26 367.385 ;
      VIA 313.49 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 361.595 314.28 361.925 ;
      VIA 313.49 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 361.575 314.26 361.945 ;
      VIA 313.49 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 356.155 314.28 356.485 ;
      VIA 313.49 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 356.135 314.26 356.505 ;
      VIA 313.49 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 350.715 314.28 351.045 ;
      VIA 313.49 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 350.695 314.26 351.065 ;
      VIA 313.49 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 345.275 314.28 345.605 ;
      VIA 313.49 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 345.255 314.26 345.625 ;
      VIA 313.49 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 339.835 314.28 340.165 ;
      VIA 313.49 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 339.815 314.26 340.185 ;
      VIA 313.49 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 334.395 314.28 334.725 ;
      VIA 313.49 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 334.375 314.26 334.745 ;
      VIA 313.49 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 328.955 314.28 329.285 ;
      VIA 313.49 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 328.935 314.26 329.305 ;
      VIA 313.49 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 323.515 314.28 323.845 ;
      VIA 313.49 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 323.495 314.26 323.865 ;
      VIA 313.49 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 318.075 314.28 318.405 ;
      VIA 313.49 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 318.055 314.26 318.425 ;
      VIA 313.49 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 312.635 314.28 312.965 ;
      VIA 313.49 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 312.615 314.26 312.985 ;
      VIA 313.49 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 307.195 314.28 307.525 ;
      VIA 313.49 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 307.175 314.26 307.545 ;
      VIA 313.49 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 301.755 314.28 302.085 ;
      VIA 313.49 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 301.735 314.26 302.105 ;
      VIA 313.49 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 296.315 314.28 296.645 ;
      VIA 313.49 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 296.295 314.26 296.665 ;
      VIA 313.49 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 290.875 314.28 291.205 ;
      VIA 313.49 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 290.855 314.26 291.225 ;
      VIA 313.49 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 285.435 314.28 285.765 ;
      VIA 313.49 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 285.415 314.26 285.785 ;
      VIA 313.49 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 279.995 314.28 280.325 ;
      VIA 313.49 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 279.975 314.26 280.345 ;
      VIA 313.49 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 274.555 314.28 274.885 ;
      VIA 313.49 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 274.535 314.26 274.905 ;
      VIA 313.49 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 269.115 314.28 269.445 ;
      VIA 313.49 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 269.095 314.26 269.465 ;
      VIA 313.49 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 263.675 314.28 264.005 ;
      VIA 313.49 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 263.655 314.26 264.025 ;
      VIA 313.49 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 258.235 314.28 258.565 ;
      VIA 313.49 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 258.215 314.26 258.585 ;
      VIA 313.49 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 252.795 314.28 253.125 ;
      VIA 313.49 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 252.775 314.26 253.145 ;
      VIA 313.49 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 247.355 314.28 247.685 ;
      VIA 313.49 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 247.335 314.26 247.705 ;
      VIA 313.49 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 241.915 314.28 242.245 ;
      VIA 313.49 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 241.895 314.26 242.265 ;
      VIA 313.49 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 236.475 314.28 236.805 ;
      VIA 313.49 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 236.455 314.26 236.825 ;
      VIA 313.49 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 231.035 314.28 231.365 ;
      VIA 313.49 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 231.015 314.26 231.385 ;
      VIA 313.49 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 225.595 314.28 225.925 ;
      VIA 313.49 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 225.575 314.26 225.945 ;
      VIA 313.49 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 220.155 314.28 220.485 ;
      VIA 313.49 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 220.135 314.26 220.505 ;
      VIA 313.49 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 214.715 314.28 215.045 ;
      VIA 313.49 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 214.695 314.26 215.065 ;
      VIA 313.49 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 209.275 314.28 209.605 ;
      VIA 313.49 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 209.255 314.26 209.625 ;
      VIA 313.49 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 203.835 314.28 204.165 ;
      VIA 313.49 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 203.815 314.26 204.185 ;
      VIA 313.49 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 198.395 314.28 198.725 ;
      VIA 313.49 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 198.375 314.26 198.745 ;
      VIA 313.49 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 192.955 314.28 193.285 ;
      VIA 313.49 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 192.935 314.26 193.305 ;
      VIA 313.49 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 187.515 314.28 187.845 ;
      VIA 313.49 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 187.495 314.26 187.865 ;
      VIA 313.49 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 182.075 314.28 182.405 ;
      VIA 313.49 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 182.055 314.26 182.425 ;
      VIA 313.49 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 176.635 314.28 176.965 ;
      VIA 313.49 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 176.615 314.26 176.985 ;
      VIA 313.49 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 171.195 314.28 171.525 ;
      VIA 313.49 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 171.175 314.26 171.545 ;
      VIA 313.49 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 165.755 314.28 166.085 ;
      VIA 313.49 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 165.735 314.26 166.105 ;
      VIA 313.49 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 160.315 314.28 160.645 ;
      VIA 313.49 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 160.295 314.26 160.665 ;
      VIA 313.49 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 154.875 314.28 155.205 ;
      VIA 313.49 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 154.855 314.26 155.225 ;
      VIA 313.49 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 149.435 314.28 149.765 ;
      VIA 313.49 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 149.415 314.26 149.785 ;
      VIA 313.49 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 143.995 314.28 144.325 ;
      VIA 313.49 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 143.975 314.26 144.345 ;
      VIA 313.49 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 138.555 314.28 138.885 ;
      VIA 313.49 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 138.535 314.26 138.905 ;
      VIA 313.49 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 133.115 314.28 133.445 ;
      VIA 313.49 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 133.095 314.26 133.465 ;
      VIA 313.49 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 127.675 314.28 128.005 ;
      VIA 313.49 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 127.655 314.26 128.025 ;
      VIA 313.49 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 122.235 314.28 122.565 ;
      VIA 313.49 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 122.215 314.26 122.585 ;
      VIA 313.49 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 116.795 314.28 117.125 ;
      VIA 313.49 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 116.775 314.26 117.145 ;
      VIA 313.49 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 111.355 314.28 111.685 ;
      VIA 313.49 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 111.335 314.26 111.705 ;
      VIA 313.49 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 105.915 314.28 106.245 ;
      VIA 313.49 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 105.895 314.26 106.265 ;
      VIA 313.49 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 100.475 314.28 100.805 ;
      VIA 313.49 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 100.455 314.26 100.825 ;
      VIA 313.49 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 95.035 314.28 95.365 ;
      VIA 313.49 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 95.015 314.26 95.385 ;
      VIA 313.49 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 89.595 314.28 89.925 ;
      VIA 313.49 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 89.575 314.26 89.945 ;
      VIA 313.49 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 84.155 314.28 84.485 ;
      VIA 313.49 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 84.135 314.26 84.505 ;
      VIA 313.49 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 78.715 314.28 79.045 ;
      VIA 313.49 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 78.695 314.26 79.065 ;
      VIA 313.49 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 73.275 314.28 73.605 ;
      VIA 313.49 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 73.255 314.26 73.625 ;
      VIA 313.49 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 67.835 314.28 68.165 ;
      VIA 313.49 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 67.815 314.26 68.185 ;
      VIA 313.49 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 62.395 314.28 62.725 ;
      VIA 313.49 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 62.375 314.26 62.745 ;
      VIA 313.49 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 56.955 314.28 57.285 ;
      VIA 313.49 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 56.935 314.26 57.305 ;
      VIA 313.49 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 51.515 314.28 51.845 ;
      VIA 313.49 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 51.495 314.26 51.865 ;
      VIA 313.49 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 46.075 314.28 46.405 ;
      VIA 313.49 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 46.055 314.26 46.425 ;
      VIA 313.49 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 40.635 314.28 40.965 ;
      VIA 313.49 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 40.615 314.26 40.985 ;
      VIA 313.49 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 35.195 314.28 35.525 ;
      VIA 313.49 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 35.175 314.26 35.545 ;
      VIA 313.49 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 29.755 314.28 30.085 ;
      VIA 313.49 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 29.735 314.26 30.105 ;
      VIA 313.49 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 24.315 314.28 24.645 ;
      VIA 313.49 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 24.295 314.26 24.665 ;
      VIA 313.49 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 18.875 314.28 19.205 ;
      VIA 313.49 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 18.855 314.26 19.225 ;
      VIA 313.49 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 13.435 314.28 13.765 ;
      VIA 313.49 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 13.415 314.26 13.785 ;
      VIA 313.49 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 7.995 314.28 8.325 ;
      VIA 313.49 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 7.975 314.26 8.345 ;
      VIA 313.49 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  312.7 2.555 314.28 2.885 ;
      VIA 313.49 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  312.72 2.535 314.26 2.905 ;
      VIA 313.49 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 313.49 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 415.995 287.14 416.325 ;
      VIA 286.35 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 415.975 287.12 416.345 ;
      VIA 286.35 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 410.555 287.14 410.885 ;
      VIA 286.35 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 410.535 287.12 410.905 ;
      VIA 286.35 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 405.115 287.14 405.445 ;
      VIA 286.35 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 405.095 287.12 405.465 ;
      VIA 286.35 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 399.675 287.14 400.005 ;
      VIA 286.35 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 399.655 287.12 400.025 ;
      VIA 286.35 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 394.235 287.14 394.565 ;
      VIA 286.35 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 394.215 287.12 394.585 ;
      VIA 286.35 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 388.795 287.14 389.125 ;
      VIA 286.35 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 388.775 287.12 389.145 ;
      VIA 286.35 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 383.355 287.14 383.685 ;
      VIA 286.35 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 383.335 287.12 383.705 ;
      VIA 286.35 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 377.915 287.14 378.245 ;
      VIA 286.35 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 377.895 287.12 378.265 ;
      VIA 286.35 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 372.475 287.14 372.805 ;
      VIA 286.35 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 372.455 287.12 372.825 ;
      VIA 286.35 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 367.035 287.14 367.365 ;
      VIA 286.35 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 367.015 287.12 367.385 ;
      VIA 286.35 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 361.595 287.14 361.925 ;
      VIA 286.35 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 361.575 287.12 361.945 ;
      VIA 286.35 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 356.155 287.14 356.485 ;
      VIA 286.35 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 356.135 287.12 356.505 ;
      VIA 286.35 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 350.715 287.14 351.045 ;
      VIA 286.35 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 350.695 287.12 351.065 ;
      VIA 286.35 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 345.275 287.14 345.605 ;
      VIA 286.35 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 345.255 287.12 345.625 ;
      VIA 286.35 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 339.835 287.14 340.165 ;
      VIA 286.35 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 339.815 287.12 340.185 ;
      VIA 286.35 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 334.395 287.14 334.725 ;
      VIA 286.35 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 334.375 287.12 334.745 ;
      VIA 286.35 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 328.955 287.14 329.285 ;
      VIA 286.35 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 328.935 287.12 329.305 ;
      VIA 286.35 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 323.515 287.14 323.845 ;
      VIA 286.35 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 323.495 287.12 323.865 ;
      VIA 286.35 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 318.075 287.14 318.405 ;
      VIA 286.35 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 318.055 287.12 318.425 ;
      VIA 286.35 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 312.635 287.14 312.965 ;
      VIA 286.35 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 312.615 287.12 312.985 ;
      VIA 286.35 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 307.195 287.14 307.525 ;
      VIA 286.35 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 307.175 287.12 307.545 ;
      VIA 286.35 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 301.755 287.14 302.085 ;
      VIA 286.35 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 301.735 287.12 302.105 ;
      VIA 286.35 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 296.315 287.14 296.645 ;
      VIA 286.35 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 296.295 287.12 296.665 ;
      VIA 286.35 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 290.875 287.14 291.205 ;
      VIA 286.35 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 290.855 287.12 291.225 ;
      VIA 286.35 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 285.435 287.14 285.765 ;
      VIA 286.35 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 285.415 287.12 285.785 ;
      VIA 286.35 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 279.995 287.14 280.325 ;
      VIA 286.35 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 279.975 287.12 280.345 ;
      VIA 286.35 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 274.555 287.14 274.885 ;
      VIA 286.35 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 274.535 287.12 274.905 ;
      VIA 286.35 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 269.115 287.14 269.445 ;
      VIA 286.35 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 269.095 287.12 269.465 ;
      VIA 286.35 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 263.675 287.14 264.005 ;
      VIA 286.35 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 263.655 287.12 264.025 ;
      VIA 286.35 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 258.235 287.14 258.565 ;
      VIA 286.35 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 258.215 287.12 258.585 ;
      VIA 286.35 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 252.795 287.14 253.125 ;
      VIA 286.35 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 252.775 287.12 253.145 ;
      VIA 286.35 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 247.355 287.14 247.685 ;
      VIA 286.35 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 247.335 287.12 247.705 ;
      VIA 286.35 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 241.915 287.14 242.245 ;
      VIA 286.35 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 241.895 287.12 242.265 ;
      VIA 286.35 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 236.475 287.14 236.805 ;
      VIA 286.35 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 236.455 287.12 236.825 ;
      VIA 286.35 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 231.035 287.14 231.365 ;
      VIA 286.35 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 231.015 287.12 231.385 ;
      VIA 286.35 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 225.595 287.14 225.925 ;
      VIA 286.35 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 225.575 287.12 225.945 ;
      VIA 286.35 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 220.155 287.14 220.485 ;
      VIA 286.35 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 220.135 287.12 220.505 ;
      VIA 286.35 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 214.715 287.14 215.045 ;
      VIA 286.35 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 214.695 287.12 215.065 ;
      VIA 286.35 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 209.275 287.14 209.605 ;
      VIA 286.35 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 209.255 287.12 209.625 ;
      VIA 286.35 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 203.835 287.14 204.165 ;
      VIA 286.35 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 203.815 287.12 204.185 ;
      VIA 286.35 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 198.395 287.14 198.725 ;
      VIA 286.35 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 198.375 287.12 198.745 ;
      VIA 286.35 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 192.955 287.14 193.285 ;
      VIA 286.35 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 192.935 287.12 193.305 ;
      VIA 286.35 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 187.515 287.14 187.845 ;
      VIA 286.35 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 187.495 287.12 187.865 ;
      VIA 286.35 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 182.075 287.14 182.405 ;
      VIA 286.35 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 182.055 287.12 182.425 ;
      VIA 286.35 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 176.635 287.14 176.965 ;
      VIA 286.35 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 176.615 287.12 176.985 ;
      VIA 286.35 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 171.195 287.14 171.525 ;
      VIA 286.35 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 171.175 287.12 171.545 ;
      VIA 286.35 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 165.755 287.14 166.085 ;
      VIA 286.35 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 165.735 287.12 166.105 ;
      VIA 286.35 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 160.315 287.14 160.645 ;
      VIA 286.35 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 160.295 287.12 160.665 ;
      VIA 286.35 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 154.875 287.14 155.205 ;
      VIA 286.35 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 154.855 287.12 155.225 ;
      VIA 286.35 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 149.435 287.14 149.765 ;
      VIA 286.35 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 149.415 287.12 149.785 ;
      VIA 286.35 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 143.995 287.14 144.325 ;
      VIA 286.35 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 143.975 287.12 144.345 ;
      VIA 286.35 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 138.555 287.14 138.885 ;
      VIA 286.35 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 138.535 287.12 138.905 ;
      VIA 286.35 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 133.115 287.14 133.445 ;
      VIA 286.35 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 133.095 287.12 133.465 ;
      VIA 286.35 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 127.675 287.14 128.005 ;
      VIA 286.35 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 127.655 287.12 128.025 ;
      VIA 286.35 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 122.235 287.14 122.565 ;
      VIA 286.35 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 122.215 287.12 122.585 ;
      VIA 286.35 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 116.795 287.14 117.125 ;
      VIA 286.35 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 116.775 287.12 117.145 ;
      VIA 286.35 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 111.355 287.14 111.685 ;
      VIA 286.35 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 111.335 287.12 111.705 ;
      VIA 286.35 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 105.915 287.14 106.245 ;
      VIA 286.35 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 105.895 287.12 106.265 ;
      VIA 286.35 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 100.475 287.14 100.805 ;
      VIA 286.35 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 100.455 287.12 100.825 ;
      VIA 286.35 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 95.035 287.14 95.365 ;
      VIA 286.35 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 95.015 287.12 95.385 ;
      VIA 286.35 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 89.595 287.14 89.925 ;
      VIA 286.35 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 89.575 287.12 89.945 ;
      VIA 286.35 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 84.155 287.14 84.485 ;
      VIA 286.35 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 84.135 287.12 84.505 ;
      VIA 286.35 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 78.715 287.14 79.045 ;
      VIA 286.35 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 78.695 287.12 79.065 ;
      VIA 286.35 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 73.275 287.14 73.605 ;
      VIA 286.35 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 73.255 287.12 73.625 ;
      VIA 286.35 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 67.835 287.14 68.165 ;
      VIA 286.35 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 67.815 287.12 68.185 ;
      VIA 286.35 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 62.395 287.14 62.725 ;
      VIA 286.35 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 62.375 287.12 62.745 ;
      VIA 286.35 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 56.955 287.14 57.285 ;
      VIA 286.35 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 56.935 287.12 57.305 ;
      VIA 286.35 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 51.515 287.14 51.845 ;
      VIA 286.35 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 51.495 287.12 51.865 ;
      VIA 286.35 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 46.075 287.14 46.405 ;
      VIA 286.35 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 46.055 287.12 46.425 ;
      VIA 286.35 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 40.635 287.14 40.965 ;
      VIA 286.35 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 40.615 287.12 40.985 ;
      VIA 286.35 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 35.195 287.14 35.525 ;
      VIA 286.35 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 35.175 287.12 35.545 ;
      VIA 286.35 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 29.755 287.14 30.085 ;
      VIA 286.35 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 29.735 287.12 30.105 ;
      VIA 286.35 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 24.315 287.14 24.645 ;
      VIA 286.35 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 24.295 287.12 24.665 ;
      VIA 286.35 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 18.875 287.14 19.205 ;
      VIA 286.35 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 18.855 287.12 19.225 ;
      VIA 286.35 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 13.435 287.14 13.765 ;
      VIA 286.35 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 13.415 287.12 13.785 ;
      VIA 286.35 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 7.995 287.14 8.325 ;
      VIA 286.35 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 7.975 287.12 8.345 ;
      VIA 286.35 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 2.555 287.14 2.885 ;
      VIA 286.35 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 2.535 287.12 2.905 ;
      VIA 286.35 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 415.995 260 416.325 ;
      VIA 259.21 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 415.975 259.98 416.345 ;
      VIA 259.21 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 410.555 260 410.885 ;
      VIA 259.21 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 410.535 259.98 410.905 ;
      VIA 259.21 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 405.115 260 405.445 ;
      VIA 259.21 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 405.095 259.98 405.465 ;
      VIA 259.21 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 399.675 260 400.005 ;
      VIA 259.21 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 399.655 259.98 400.025 ;
      VIA 259.21 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 394.235 260 394.565 ;
      VIA 259.21 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 394.215 259.98 394.585 ;
      VIA 259.21 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 388.795 260 389.125 ;
      VIA 259.21 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 388.775 259.98 389.145 ;
      VIA 259.21 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 383.355 260 383.685 ;
      VIA 259.21 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 383.335 259.98 383.705 ;
      VIA 259.21 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 377.915 260 378.245 ;
      VIA 259.21 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 377.895 259.98 378.265 ;
      VIA 259.21 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 372.475 260 372.805 ;
      VIA 259.21 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 372.455 259.98 372.825 ;
      VIA 259.21 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 367.035 260 367.365 ;
      VIA 259.21 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 367.015 259.98 367.385 ;
      VIA 259.21 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 361.595 260 361.925 ;
      VIA 259.21 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 361.575 259.98 361.945 ;
      VIA 259.21 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 356.155 260 356.485 ;
      VIA 259.21 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 356.135 259.98 356.505 ;
      VIA 259.21 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 350.715 260 351.045 ;
      VIA 259.21 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 350.695 259.98 351.065 ;
      VIA 259.21 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 345.275 260 345.605 ;
      VIA 259.21 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 345.255 259.98 345.625 ;
      VIA 259.21 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 339.835 260 340.165 ;
      VIA 259.21 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 339.815 259.98 340.185 ;
      VIA 259.21 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 334.395 260 334.725 ;
      VIA 259.21 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 334.375 259.98 334.745 ;
      VIA 259.21 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 328.955 260 329.285 ;
      VIA 259.21 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 328.935 259.98 329.305 ;
      VIA 259.21 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 323.515 260 323.845 ;
      VIA 259.21 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 323.495 259.98 323.865 ;
      VIA 259.21 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 318.075 260 318.405 ;
      VIA 259.21 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 318.055 259.98 318.425 ;
      VIA 259.21 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 312.635 260 312.965 ;
      VIA 259.21 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 312.615 259.98 312.985 ;
      VIA 259.21 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 307.195 260 307.525 ;
      VIA 259.21 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 307.175 259.98 307.545 ;
      VIA 259.21 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 301.755 260 302.085 ;
      VIA 259.21 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 301.735 259.98 302.105 ;
      VIA 259.21 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 296.315 260 296.645 ;
      VIA 259.21 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 296.295 259.98 296.665 ;
      VIA 259.21 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 290.875 260 291.205 ;
      VIA 259.21 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 290.855 259.98 291.225 ;
      VIA 259.21 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 285.435 260 285.765 ;
      VIA 259.21 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 285.415 259.98 285.785 ;
      VIA 259.21 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 279.995 260 280.325 ;
      VIA 259.21 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 279.975 259.98 280.345 ;
      VIA 259.21 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 274.555 260 274.885 ;
      VIA 259.21 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 274.535 259.98 274.905 ;
      VIA 259.21 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 269.115 260 269.445 ;
      VIA 259.21 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 269.095 259.98 269.465 ;
      VIA 259.21 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 263.675 260 264.005 ;
      VIA 259.21 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 263.655 259.98 264.025 ;
      VIA 259.21 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 258.235 260 258.565 ;
      VIA 259.21 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 258.215 259.98 258.585 ;
      VIA 259.21 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 252.795 260 253.125 ;
      VIA 259.21 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 252.775 259.98 253.145 ;
      VIA 259.21 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 247.355 260 247.685 ;
      VIA 259.21 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 247.335 259.98 247.705 ;
      VIA 259.21 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 241.915 260 242.245 ;
      VIA 259.21 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 241.895 259.98 242.265 ;
      VIA 259.21 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 236.475 260 236.805 ;
      VIA 259.21 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 236.455 259.98 236.825 ;
      VIA 259.21 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 231.035 260 231.365 ;
      VIA 259.21 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 231.015 259.98 231.385 ;
      VIA 259.21 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 225.595 260 225.925 ;
      VIA 259.21 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 225.575 259.98 225.945 ;
      VIA 259.21 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 220.155 260 220.485 ;
      VIA 259.21 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 220.135 259.98 220.505 ;
      VIA 259.21 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 214.715 260 215.045 ;
      VIA 259.21 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 214.695 259.98 215.065 ;
      VIA 259.21 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 209.275 260 209.605 ;
      VIA 259.21 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 209.255 259.98 209.625 ;
      VIA 259.21 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 203.835 260 204.165 ;
      VIA 259.21 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 203.815 259.98 204.185 ;
      VIA 259.21 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 198.395 260 198.725 ;
      VIA 259.21 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 198.375 259.98 198.745 ;
      VIA 259.21 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 192.955 260 193.285 ;
      VIA 259.21 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 192.935 259.98 193.305 ;
      VIA 259.21 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 187.515 260 187.845 ;
      VIA 259.21 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 187.495 259.98 187.865 ;
      VIA 259.21 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 182.075 260 182.405 ;
      VIA 259.21 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 182.055 259.98 182.425 ;
      VIA 259.21 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 176.635 260 176.965 ;
      VIA 259.21 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 176.615 259.98 176.985 ;
      VIA 259.21 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 171.195 260 171.525 ;
      VIA 259.21 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 171.175 259.98 171.545 ;
      VIA 259.21 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 165.755 260 166.085 ;
      VIA 259.21 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 165.735 259.98 166.105 ;
      VIA 259.21 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 160.315 260 160.645 ;
      VIA 259.21 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 160.295 259.98 160.665 ;
      VIA 259.21 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 154.875 260 155.205 ;
      VIA 259.21 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 154.855 259.98 155.225 ;
      VIA 259.21 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 149.435 260 149.765 ;
      VIA 259.21 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 149.415 259.98 149.785 ;
      VIA 259.21 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 143.995 260 144.325 ;
      VIA 259.21 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 143.975 259.98 144.345 ;
      VIA 259.21 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 138.555 260 138.885 ;
      VIA 259.21 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 138.535 259.98 138.905 ;
      VIA 259.21 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 133.115 260 133.445 ;
      VIA 259.21 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 133.095 259.98 133.465 ;
      VIA 259.21 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 127.675 260 128.005 ;
      VIA 259.21 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 127.655 259.98 128.025 ;
      VIA 259.21 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 122.235 260 122.565 ;
      VIA 259.21 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 122.215 259.98 122.585 ;
      VIA 259.21 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 116.795 260 117.125 ;
      VIA 259.21 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 116.775 259.98 117.145 ;
      VIA 259.21 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 111.355 260 111.685 ;
      VIA 259.21 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 111.335 259.98 111.705 ;
      VIA 259.21 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 105.915 260 106.245 ;
      VIA 259.21 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 105.895 259.98 106.265 ;
      VIA 259.21 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 100.475 260 100.805 ;
      VIA 259.21 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 100.455 259.98 100.825 ;
      VIA 259.21 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 95.035 260 95.365 ;
      VIA 259.21 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 95.015 259.98 95.385 ;
      VIA 259.21 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 89.595 260 89.925 ;
      VIA 259.21 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 89.575 259.98 89.945 ;
      VIA 259.21 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 84.155 260 84.485 ;
      VIA 259.21 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 84.135 259.98 84.505 ;
      VIA 259.21 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 78.715 260 79.045 ;
      VIA 259.21 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 78.695 259.98 79.065 ;
      VIA 259.21 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 73.275 260 73.605 ;
      VIA 259.21 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 73.255 259.98 73.625 ;
      VIA 259.21 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 67.835 260 68.165 ;
      VIA 259.21 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 67.815 259.98 68.185 ;
      VIA 259.21 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 62.395 260 62.725 ;
      VIA 259.21 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 62.375 259.98 62.745 ;
      VIA 259.21 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 56.955 260 57.285 ;
      VIA 259.21 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 56.935 259.98 57.305 ;
      VIA 259.21 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 51.515 260 51.845 ;
      VIA 259.21 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 51.495 259.98 51.865 ;
      VIA 259.21 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 46.075 260 46.405 ;
      VIA 259.21 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 46.055 259.98 46.425 ;
      VIA 259.21 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 40.635 260 40.965 ;
      VIA 259.21 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 40.615 259.98 40.985 ;
      VIA 259.21 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 35.195 260 35.525 ;
      VIA 259.21 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 35.175 259.98 35.545 ;
      VIA 259.21 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 29.755 260 30.085 ;
      VIA 259.21 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 29.735 259.98 30.105 ;
      VIA 259.21 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 24.315 260 24.645 ;
      VIA 259.21 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 24.295 259.98 24.665 ;
      VIA 259.21 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 18.875 260 19.205 ;
      VIA 259.21 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 18.855 259.98 19.225 ;
      VIA 259.21 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 13.435 260 13.765 ;
      VIA 259.21 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 13.415 259.98 13.785 ;
      VIA 259.21 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 7.995 260 8.325 ;
      VIA 259.21 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 7.975 259.98 8.345 ;
      VIA 259.21 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 2.555 260 2.885 ;
      VIA 259.21 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 2.535 259.98 2.905 ;
      VIA 259.21 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 415.995 232.86 416.325 ;
      VIA 232.07 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 415.975 232.84 416.345 ;
      VIA 232.07 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 410.555 232.86 410.885 ;
      VIA 232.07 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 410.535 232.84 410.905 ;
      VIA 232.07 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 405.115 232.86 405.445 ;
      VIA 232.07 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 405.095 232.84 405.465 ;
      VIA 232.07 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 399.675 232.86 400.005 ;
      VIA 232.07 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 399.655 232.84 400.025 ;
      VIA 232.07 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 394.235 232.86 394.565 ;
      VIA 232.07 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 394.215 232.84 394.585 ;
      VIA 232.07 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 388.795 232.86 389.125 ;
      VIA 232.07 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 388.775 232.84 389.145 ;
      VIA 232.07 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 383.355 232.86 383.685 ;
      VIA 232.07 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 383.335 232.84 383.705 ;
      VIA 232.07 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 377.915 232.86 378.245 ;
      VIA 232.07 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 377.895 232.84 378.265 ;
      VIA 232.07 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 372.475 232.86 372.805 ;
      VIA 232.07 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 372.455 232.84 372.825 ;
      VIA 232.07 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 367.035 232.86 367.365 ;
      VIA 232.07 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 367.015 232.84 367.385 ;
      VIA 232.07 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 361.595 232.86 361.925 ;
      VIA 232.07 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 361.575 232.84 361.945 ;
      VIA 232.07 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 356.155 232.86 356.485 ;
      VIA 232.07 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 356.135 232.84 356.505 ;
      VIA 232.07 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 350.715 232.86 351.045 ;
      VIA 232.07 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 350.695 232.84 351.065 ;
      VIA 232.07 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 345.275 232.86 345.605 ;
      VIA 232.07 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 345.255 232.84 345.625 ;
      VIA 232.07 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 339.835 232.86 340.165 ;
      VIA 232.07 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 339.815 232.84 340.185 ;
      VIA 232.07 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 334.395 232.86 334.725 ;
      VIA 232.07 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 334.375 232.84 334.745 ;
      VIA 232.07 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 328.955 232.86 329.285 ;
      VIA 232.07 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 328.935 232.84 329.305 ;
      VIA 232.07 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 323.515 232.86 323.845 ;
      VIA 232.07 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 323.495 232.84 323.865 ;
      VIA 232.07 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 318.075 232.86 318.405 ;
      VIA 232.07 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 318.055 232.84 318.425 ;
      VIA 232.07 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 312.635 232.86 312.965 ;
      VIA 232.07 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 312.615 232.84 312.985 ;
      VIA 232.07 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 307.195 232.86 307.525 ;
      VIA 232.07 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 307.175 232.84 307.545 ;
      VIA 232.07 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 301.755 232.86 302.085 ;
      VIA 232.07 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 301.735 232.84 302.105 ;
      VIA 232.07 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 296.315 232.86 296.645 ;
      VIA 232.07 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 296.295 232.84 296.665 ;
      VIA 232.07 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 290.875 232.86 291.205 ;
      VIA 232.07 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 290.855 232.84 291.225 ;
      VIA 232.07 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 285.435 232.86 285.765 ;
      VIA 232.07 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 285.415 232.84 285.785 ;
      VIA 232.07 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 279.995 232.86 280.325 ;
      VIA 232.07 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 279.975 232.84 280.345 ;
      VIA 232.07 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 274.555 232.86 274.885 ;
      VIA 232.07 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 274.535 232.84 274.905 ;
      VIA 232.07 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 269.115 232.86 269.445 ;
      VIA 232.07 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 269.095 232.84 269.465 ;
      VIA 232.07 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 263.675 232.86 264.005 ;
      VIA 232.07 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 263.655 232.84 264.025 ;
      VIA 232.07 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 258.235 232.86 258.565 ;
      VIA 232.07 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 258.215 232.84 258.585 ;
      VIA 232.07 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 252.795 232.86 253.125 ;
      VIA 232.07 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 252.775 232.84 253.145 ;
      VIA 232.07 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 247.355 232.86 247.685 ;
      VIA 232.07 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 247.335 232.84 247.705 ;
      VIA 232.07 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 241.915 232.86 242.245 ;
      VIA 232.07 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 241.895 232.84 242.265 ;
      VIA 232.07 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 236.475 232.86 236.805 ;
      VIA 232.07 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 236.455 232.84 236.825 ;
      VIA 232.07 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 231.035 232.86 231.365 ;
      VIA 232.07 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 231.015 232.84 231.385 ;
      VIA 232.07 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 225.595 232.86 225.925 ;
      VIA 232.07 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 225.575 232.84 225.945 ;
      VIA 232.07 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 220.155 232.86 220.485 ;
      VIA 232.07 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 220.135 232.84 220.505 ;
      VIA 232.07 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 214.715 232.86 215.045 ;
      VIA 232.07 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 214.695 232.84 215.065 ;
      VIA 232.07 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 209.275 232.86 209.605 ;
      VIA 232.07 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 209.255 232.84 209.625 ;
      VIA 232.07 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 203.835 232.86 204.165 ;
      VIA 232.07 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 203.815 232.84 204.185 ;
      VIA 232.07 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 198.395 232.86 198.725 ;
      VIA 232.07 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 198.375 232.84 198.745 ;
      VIA 232.07 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 192.955 232.86 193.285 ;
      VIA 232.07 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 192.935 232.84 193.305 ;
      VIA 232.07 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 187.515 232.86 187.845 ;
      VIA 232.07 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 187.495 232.84 187.865 ;
      VIA 232.07 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 182.075 232.86 182.405 ;
      VIA 232.07 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 182.055 232.84 182.425 ;
      VIA 232.07 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 176.635 232.86 176.965 ;
      VIA 232.07 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 176.615 232.84 176.985 ;
      VIA 232.07 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 171.195 232.86 171.525 ;
      VIA 232.07 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 171.175 232.84 171.545 ;
      VIA 232.07 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 165.755 232.86 166.085 ;
      VIA 232.07 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 165.735 232.84 166.105 ;
      VIA 232.07 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 160.315 232.86 160.645 ;
      VIA 232.07 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 160.295 232.84 160.665 ;
      VIA 232.07 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 154.875 232.86 155.205 ;
      VIA 232.07 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 154.855 232.84 155.225 ;
      VIA 232.07 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 149.435 232.86 149.765 ;
      VIA 232.07 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 149.415 232.84 149.785 ;
      VIA 232.07 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 143.995 232.86 144.325 ;
      VIA 232.07 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 143.975 232.84 144.345 ;
      VIA 232.07 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 138.555 232.86 138.885 ;
      VIA 232.07 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 138.535 232.84 138.905 ;
      VIA 232.07 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 133.115 232.86 133.445 ;
      VIA 232.07 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 133.095 232.84 133.465 ;
      VIA 232.07 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 127.675 232.86 128.005 ;
      VIA 232.07 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 127.655 232.84 128.025 ;
      VIA 232.07 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 122.235 232.86 122.565 ;
      VIA 232.07 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 122.215 232.84 122.585 ;
      VIA 232.07 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 116.795 232.86 117.125 ;
      VIA 232.07 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 116.775 232.84 117.145 ;
      VIA 232.07 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 111.355 232.86 111.685 ;
      VIA 232.07 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 111.335 232.84 111.705 ;
      VIA 232.07 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 105.915 232.86 106.245 ;
      VIA 232.07 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 105.895 232.84 106.265 ;
      VIA 232.07 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 100.475 232.86 100.805 ;
      VIA 232.07 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 100.455 232.84 100.825 ;
      VIA 232.07 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 95.035 232.86 95.365 ;
      VIA 232.07 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 95.015 232.84 95.385 ;
      VIA 232.07 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 89.595 232.86 89.925 ;
      VIA 232.07 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 89.575 232.84 89.945 ;
      VIA 232.07 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 84.155 232.86 84.485 ;
      VIA 232.07 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 84.135 232.84 84.505 ;
      VIA 232.07 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 78.715 232.86 79.045 ;
      VIA 232.07 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 78.695 232.84 79.065 ;
      VIA 232.07 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 73.275 232.86 73.605 ;
      VIA 232.07 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 73.255 232.84 73.625 ;
      VIA 232.07 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 67.835 232.86 68.165 ;
      VIA 232.07 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 67.815 232.84 68.185 ;
      VIA 232.07 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 62.395 232.86 62.725 ;
      VIA 232.07 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 62.375 232.84 62.745 ;
      VIA 232.07 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 56.955 232.86 57.285 ;
      VIA 232.07 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 56.935 232.84 57.305 ;
      VIA 232.07 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 51.515 232.86 51.845 ;
      VIA 232.07 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 51.495 232.84 51.865 ;
      VIA 232.07 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 46.075 232.86 46.405 ;
      VIA 232.07 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 46.055 232.84 46.425 ;
      VIA 232.07 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 40.635 232.86 40.965 ;
      VIA 232.07 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 40.615 232.84 40.985 ;
      VIA 232.07 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 35.195 232.86 35.525 ;
      VIA 232.07 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 35.175 232.84 35.545 ;
      VIA 232.07 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 29.755 232.86 30.085 ;
      VIA 232.07 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 29.735 232.84 30.105 ;
      VIA 232.07 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 24.315 232.86 24.645 ;
      VIA 232.07 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 24.295 232.84 24.665 ;
      VIA 232.07 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 18.875 232.86 19.205 ;
      VIA 232.07 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 18.855 232.84 19.225 ;
      VIA 232.07 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 13.435 232.86 13.765 ;
      VIA 232.07 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 13.415 232.84 13.785 ;
      VIA 232.07 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 7.995 232.86 8.325 ;
      VIA 232.07 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 7.975 232.84 8.345 ;
      VIA 232.07 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 2.555 232.86 2.885 ;
      VIA 232.07 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 2.535 232.84 2.905 ;
      VIA 232.07 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 415.995 205.72 416.325 ;
      VIA 204.93 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 415.975 205.7 416.345 ;
      VIA 204.93 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 410.555 205.72 410.885 ;
      VIA 204.93 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 410.535 205.7 410.905 ;
      VIA 204.93 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 405.115 205.72 405.445 ;
      VIA 204.93 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 405.095 205.7 405.465 ;
      VIA 204.93 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 399.675 205.72 400.005 ;
      VIA 204.93 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 399.655 205.7 400.025 ;
      VIA 204.93 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 394.235 205.72 394.565 ;
      VIA 204.93 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 394.215 205.7 394.585 ;
      VIA 204.93 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 388.795 205.72 389.125 ;
      VIA 204.93 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 388.775 205.7 389.145 ;
      VIA 204.93 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 383.355 205.72 383.685 ;
      VIA 204.93 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 383.335 205.7 383.705 ;
      VIA 204.93 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 377.915 205.72 378.245 ;
      VIA 204.93 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 377.895 205.7 378.265 ;
      VIA 204.93 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 372.475 205.72 372.805 ;
      VIA 204.93 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 372.455 205.7 372.825 ;
      VIA 204.93 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 367.035 205.72 367.365 ;
      VIA 204.93 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 367.015 205.7 367.385 ;
      VIA 204.93 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 361.595 205.72 361.925 ;
      VIA 204.93 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 361.575 205.7 361.945 ;
      VIA 204.93 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 356.155 205.72 356.485 ;
      VIA 204.93 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 356.135 205.7 356.505 ;
      VIA 204.93 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 350.715 205.72 351.045 ;
      VIA 204.93 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 350.695 205.7 351.065 ;
      VIA 204.93 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 345.275 205.72 345.605 ;
      VIA 204.93 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 345.255 205.7 345.625 ;
      VIA 204.93 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 339.835 205.72 340.165 ;
      VIA 204.93 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 339.815 205.7 340.185 ;
      VIA 204.93 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 334.395 205.72 334.725 ;
      VIA 204.93 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 334.375 205.7 334.745 ;
      VIA 204.93 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 328.955 205.72 329.285 ;
      VIA 204.93 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 328.935 205.7 329.305 ;
      VIA 204.93 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 323.515 205.72 323.845 ;
      VIA 204.93 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 323.495 205.7 323.865 ;
      VIA 204.93 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 318.075 205.72 318.405 ;
      VIA 204.93 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 318.055 205.7 318.425 ;
      VIA 204.93 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 312.635 205.72 312.965 ;
      VIA 204.93 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 312.615 205.7 312.985 ;
      VIA 204.93 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 307.195 205.72 307.525 ;
      VIA 204.93 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 307.175 205.7 307.545 ;
      VIA 204.93 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 301.755 205.72 302.085 ;
      VIA 204.93 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 301.735 205.7 302.105 ;
      VIA 204.93 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 296.315 205.72 296.645 ;
      VIA 204.93 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 296.295 205.7 296.665 ;
      VIA 204.93 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 290.875 205.72 291.205 ;
      VIA 204.93 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 290.855 205.7 291.225 ;
      VIA 204.93 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 285.435 205.72 285.765 ;
      VIA 204.93 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 285.415 205.7 285.785 ;
      VIA 204.93 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 279.995 205.72 280.325 ;
      VIA 204.93 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 279.975 205.7 280.345 ;
      VIA 204.93 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 274.555 205.72 274.885 ;
      VIA 204.93 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 274.535 205.7 274.905 ;
      VIA 204.93 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 269.115 205.72 269.445 ;
      VIA 204.93 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 269.095 205.7 269.465 ;
      VIA 204.93 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 263.675 205.72 264.005 ;
      VIA 204.93 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 263.655 205.7 264.025 ;
      VIA 204.93 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 258.235 205.72 258.565 ;
      VIA 204.93 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 258.215 205.7 258.585 ;
      VIA 204.93 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 252.795 205.72 253.125 ;
      VIA 204.93 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 252.775 205.7 253.145 ;
      VIA 204.93 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 247.355 205.72 247.685 ;
      VIA 204.93 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 247.335 205.7 247.705 ;
      VIA 204.93 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 241.915 205.72 242.245 ;
      VIA 204.93 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 241.895 205.7 242.265 ;
      VIA 204.93 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 236.475 205.72 236.805 ;
      VIA 204.93 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 236.455 205.7 236.825 ;
      VIA 204.93 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 231.035 205.72 231.365 ;
      VIA 204.93 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 231.015 205.7 231.385 ;
      VIA 204.93 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 225.595 205.72 225.925 ;
      VIA 204.93 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 225.575 205.7 225.945 ;
      VIA 204.93 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 220.155 205.72 220.485 ;
      VIA 204.93 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 220.135 205.7 220.505 ;
      VIA 204.93 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 214.715 205.72 215.045 ;
      VIA 204.93 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 214.695 205.7 215.065 ;
      VIA 204.93 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 209.275 205.72 209.605 ;
      VIA 204.93 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 209.255 205.7 209.625 ;
      VIA 204.93 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 203.835 205.72 204.165 ;
      VIA 204.93 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 203.815 205.7 204.185 ;
      VIA 204.93 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 198.395 205.72 198.725 ;
      VIA 204.93 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 198.375 205.7 198.745 ;
      VIA 204.93 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 192.955 205.72 193.285 ;
      VIA 204.93 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 192.935 205.7 193.305 ;
      VIA 204.93 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 187.515 205.72 187.845 ;
      VIA 204.93 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 187.495 205.7 187.865 ;
      VIA 204.93 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 182.075 205.72 182.405 ;
      VIA 204.93 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 182.055 205.7 182.425 ;
      VIA 204.93 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 176.635 205.72 176.965 ;
      VIA 204.93 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 176.615 205.7 176.985 ;
      VIA 204.93 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 171.195 205.72 171.525 ;
      VIA 204.93 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 171.175 205.7 171.545 ;
      VIA 204.93 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 165.755 205.72 166.085 ;
      VIA 204.93 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 165.735 205.7 166.105 ;
      VIA 204.93 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 160.315 205.72 160.645 ;
      VIA 204.93 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 160.295 205.7 160.665 ;
      VIA 204.93 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 154.875 205.72 155.205 ;
      VIA 204.93 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 154.855 205.7 155.225 ;
      VIA 204.93 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 149.435 205.72 149.765 ;
      VIA 204.93 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 149.415 205.7 149.785 ;
      VIA 204.93 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 143.995 205.72 144.325 ;
      VIA 204.93 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 143.975 205.7 144.345 ;
      VIA 204.93 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 138.555 205.72 138.885 ;
      VIA 204.93 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 138.535 205.7 138.905 ;
      VIA 204.93 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 133.115 205.72 133.445 ;
      VIA 204.93 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 133.095 205.7 133.465 ;
      VIA 204.93 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 127.675 205.72 128.005 ;
      VIA 204.93 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 127.655 205.7 128.025 ;
      VIA 204.93 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 122.235 205.72 122.565 ;
      VIA 204.93 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 122.215 205.7 122.585 ;
      VIA 204.93 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 116.795 205.72 117.125 ;
      VIA 204.93 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 116.775 205.7 117.145 ;
      VIA 204.93 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 111.355 205.72 111.685 ;
      VIA 204.93 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 111.335 205.7 111.705 ;
      VIA 204.93 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 105.915 205.72 106.245 ;
      VIA 204.93 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 105.895 205.7 106.265 ;
      VIA 204.93 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 100.475 205.72 100.805 ;
      VIA 204.93 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 100.455 205.7 100.825 ;
      VIA 204.93 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 95.035 205.72 95.365 ;
      VIA 204.93 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 95.015 205.7 95.385 ;
      VIA 204.93 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 89.595 205.72 89.925 ;
      VIA 204.93 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 89.575 205.7 89.945 ;
      VIA 204.93 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 84.155 205.72 84.485 ;
      VIA 204.93 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 84.135 205.7 84.505 ;
      VIA 204.93 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 78.715 205.72 79.045 ;
      VIA 204.93 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 78.695 205.7 79.065 ;
      VIA 204.93 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 73.275 205.72 73.605 ;
      VIA 204.93 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 73.255 205.7 73.625 ;
      VIA 204.93 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 67.835 205.72 68.165 ;
      VIA 204.93 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 67.815 205.7 68.185 ;
      VIA 204.93 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 62.395 205.72 62.725 ;
      VIA 204.93 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 62.375 205.7 62.745 ;
      VIA 204.93 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 56.955 205.72 57.285 ;
      VIA 204.93 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 56.935 205.7 57.305 ;
      VIA 204.93 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 51.515 205.72 51.845 ;
      VIA 204.93 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 51.495 205.7 51.865 ;
      VIA 204.93 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 46.075 205.72 46.405 ;
      VIA 204.93 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 46.055 205.7 46.425 ;
      VIA 204.93 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 40.635 205.72 40.965 ;
      VIA 204.93 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 40.615 205.7 40.985 ;
      VIA 204.93 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 35.195 205.72 35.525 ;
      VIA 204.93 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 35.175 205.7 35.545 ;
      VIA 204.93 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 29.755 205.72 30.085 ;
      VIA 204.93 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 29.735 205.7 30.105 ;
      VIA 204.93 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 24.315 205.72 24.645 ;
      VIA 204.93 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 24.295 205.7 24.665 ;
      VIA 204.93 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 18.875 205.72 19.205 ;
      VIA 204.93 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 18.855 205.7 19.225 ;
      VIA 204.93 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 13.435 205.72 13.765 ;
      VIA 204.93 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 13.415 205.7 13.785 ;
      VIA 204.93 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 7.995 205.72 8.325 ;
      VIA 204.93 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 7.975 205.7 8.345 ;
      VIA 204.93 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 2.555 205.72 2.885 ;
      VIA 204.93 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 2.535 205.7 2.905 ;
      VIA 204.93 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 415.995 178.58 416.325 ;
      VIA 177.79 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 415.975 178.56 416.345 ;
      VIA 177.79 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 410.555 178.58 410.885 ;
      VIA 177.79 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 410.535 178.56 410.905 ;
      VIA 177.79 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 405.115 178.58 405.445 ;
      VIA 177.79 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 405.095 178.56 405.465 ;
      VIA 177.79 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 399.675 178.58 400.005 ;
      VIA 177.79 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 399.655 178.56 400.025 ;
      VIA 177.79 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 394.235 178.58 394.565 ;
      VIA 177.79 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 394.215 178.56 394.585 ;
      VIA 177.79 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 388.795 178.58 389.125 ;
      VIA 177.79 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 388.775 178.56 389.145 ;
      VIA 177.79 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 383.355 178.58 383.685 ;
      VIA 177.79 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 383.335 178.56 383.705 ;
      VIA 177.79 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 377.915 178.58 378.245 ;
      VIA 177.79 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 377.895 178.56 378.265 ;
      VIA 177.79 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 372.475 178.58 372.805 ;
      VIA 177.79 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 372.455 178.56 372.825 ;
      VIA 177.79 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 367.035 178.58 367.365 ;
      VIA 177.79 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 367.015 178.56 367.385 ;
      VIA 177.79 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 361.595 178.58 361.925 ;
      VIA 177.79 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 361.575 178.56 361.945 ;
      VIA 177.79 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 356.155 178.58 356.485 ;
      VIA 177.79 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 356.135 178.56 356.505 ;
      VIA 177.79 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 350.715 178.58 351.045 ;
      VIA 177.79 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 350.695 178.56 351.065 ;
      VIA 177.79 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 345.275 178.58 345.605 ;
      VIA 177.79 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 345.255 178.56 345.625 ;
      VIA 177.79 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 339.835 178.58 340.165 ;
      VIA 177.79 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 339.815 178.56 340.185 ;
      VIA 177.79 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 334.395 178.58 334.725 ;
      VIA 177.79 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 334.375 178.56 334.745 ;
      VIA 177.79 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 328.955 178.58 329.285 ;
      VIA 177.79 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 328.935 178.56 329.305 ;
      VIA 177.79 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 323.515 178.58 323.845 ;
      VIA 177.79 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 323.495 178.56 323.865 ;
      VIA 177.79 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 318.075 178.58 318.405 ;
      VIA 177.79 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 318.055 178.56 318.425 ;
      VIA 177.79 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 312.635 178.58 312.965 ;
      VIA 177.79 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 312.615 178.56 312.985 ;
      VIA 177.79 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 307.195 178.58 307.525 ;
      VIA 177.79 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 307.175 178.56 307.545 ;
      VIA 177.79 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 301.755 178.58 302.085 ;
      VIA 177.79 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 301.735 178.56 302.105 ;
      VIA 177.79 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 296.315 178.58 296.645 ;
      VIA 177.79 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 296.295 178.56 296.665 ;
      VIA 177.79 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 290.875 178.58 291.205 ;
      VIA 177.79 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 290.855 178.56 291.225 ;
      VIA 177.79 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 285.435 178.58 285.765 ;
      VIA 177.79 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 285.415 178.56 285.785 ;
      VIA 177.79 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 279.995 178.58 280.325 ;
      VIA 177.79 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 279.975 178.56 280.345 ;
      VIA 177.79 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 274.555 178.58 274.885 ;
      VIA 177.79 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 274.535 178.56 274.905 ;
      VIA 177.79 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 269.115 178.58 269.445 ;
      VIA 177.79 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 269.095 178.56 269.465 ;
      VIA 177.79 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 263.675 178.58 264.005 ;
      VIA 177.79 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 263.655 178.56 264.025 ;
      VIA 177.79 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 258.235 178.58 258.565 ;
      VIA 177.79 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 258.215 178.56 258.585 ;
      VIA 177.79 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 252.795 178.58 253.125 ;
      VIA 177.79 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 252.775 178.56 253.145 ;
      VIA 177.79 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 247.355 178.58 247.685 ;
      VIA 177.79 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 247.335 178.56 247.705 ;
      VIA 177.79 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 241.915 178.58 242.245 ;
      VIA 177.79 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 241.895 178.56 242.265 ;
      VIA 177.79 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 236.475 178.58 236.805 ;
      VIA 177.79 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 236.455 178.56 236.825 ;
      VIA 177.79 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 231.035 178.58 231.365 ;
      VIA 177.79 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 231.015 178.56 231.385 ;
      VIA 177.79 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 225.595 178.58 225.925 ;
      VIA 177.79 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 225.575 178.56 225.945 ;
      VIA 177.79 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 220.155 178.58 220.485 ;
      VIA 177.79 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 220.135 178.56 220.505 ;
      VIA 177.79 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 214.715 178.58 215.045 ;
      VIA 177.79 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 214.695 178.56 215.065 ;
      VIA 177.79 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 209.275 178.58 209.605 ;
      VIA 177.79 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 209.255 178.56 209.625 ;
      VIA 177.79 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 203.835 178.58 204.165 ;
      VIA 177.79 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 203.815 178.56 204.185 ;
      VIA 177.79 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 198.395 178.58 198.725 ;
      VIA 177.79 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 198.375 178.56 198.745 ;
      VIA 177.79 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 192.955 178.58 193.285 ;
      VIA 177.79 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 192.935 178.56 193.305 ;
      VIA 177.79 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 187.515 178.58 187.845 ;
      VIA 177.79 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 187.495 178.56 187.865 ;
      VIA 177.79 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 182.075 178.58 182.405 ;
      VIA 177.79 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 182.055 178.56 182.425 ;
      VIA 177.79 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 176.635 178.58 176.965 ;
      VIA 177.79 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 176.615 178.56 176.985 ;
      VIA 177.79 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 171.195 178.58 171.525 ;
      VIA 177.79 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 171.175 178.56 171.545 ;
      VIA 177.79 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 165.755 178.58 166.085 ;
      VIA 177.79 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 165.735 178.56 166.105 ;
      VIA 177.79 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 160.315 178.58 160.645 ;
      VIA 177.79 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 160.295 178.56 160.665 ;
      VIA 177.79 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 154.875 178.58 155.205 ;
      VIA 177.79 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 154.855 178.56 155.225 ;
      VIA 177.79 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 149.435 178.58 149.765 ;
      VIA 177.79 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 149.415 178.56 149.785 ;
      VIA 177.79 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 143.995 178.58 144.325 ;
      VIA 177.79 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 143.975 178.56 144.345 ;
      VIA 177.79 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 138.555 178.58 138.885 ;
      VIA 177.79 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 138.535 178.56 138.905 ;
      VIA 177.79 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 133.115 178.58 133.445 ;
      VIA 177.79 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 133.095 178.56 133.465 ;
      VIA 177.79 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 127.675 178.58 128.005 ;
      VIA 177.79 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 127.655 178.56 128.025 ;
      VIA 177.79 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 122.235 178.58 122.565 ;
      VIA 177.79 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 122.215 178.56 122.585 ;
      VIA 177.79 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 116.795 178.58 117.125 ;
      VIA 177.79 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 116.775 178.56 117.145 ;
      VIA 177.79 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 111.355 178.58 111.685 ;
      VIA 177.79 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 111.335 178.56 111.705 ;
      VIA 177.79 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 105.915 178.58 106.245 ;
      VIA 177.79 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 105.895 178.56 106.265 ;
      VIA 177.79 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 100.475 178.58 100.805 ;
      VIA 177.79 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 100.455 178.56 100.825 ;
      VIA 177.79 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 95.035 178.58 95.365 ;
      VIA 177.79 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 95.015 178.56 95.385 ;
      VIA 177.79 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 89.595 178.58 89.925 ;
      VIA 177.79 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 89.575 178.56 89.945 ;
      VIA 177.79 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 84.155 178.58 84.485 ;
      VIA 177.79 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 84.135 178.56 84.505 ;
      VIA 177.79 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 78.715 178.58 79.045 ;
      VIA 177.79 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 78.695 178.56 79.065 ;
      VIA 177.79 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 73.275 178.58 73.605 ;
      VIA 177.79 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 73.255 178.56 73.625 ;
      VIA 177.79 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 67.835 178.58 68.165 ;
      VIA 177.79 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 67.815 178.56 68.185 ;
      VIA 177.79 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 62.395 178.58 62.725 ;
      VIA 177.79 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 62.375 178.56 62.745 ;
      VIA 177.79 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 56.955 178.58 57.285 ;
      VIA 177.79 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 56.935 178.56 57.305 ;
      VIA 177.79 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 51.515 178.58 51.845 ;
      VIA 177.79 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 51.495 178.56 51.865 ;
      VIA 177.79 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 46.075 178.58 46.405 ;
      VIA 177.79 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 46.055 178.56 46.425 ;
      VIA 177.79 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 40.635 178.58 40.965 ;
      VIA 177.79 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 40.615 178.56 40.985 ;
      VIA 177.79 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 35.195 178.58 35.525 ;
      VIA 177.79 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 35.175 178.56 35.545 ;
      VIA 177.79 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 29.755 178.58 30.085 ;
      VIA 177.79 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 29.735 178.56 30.105 ;
      VIA 177.79 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 24.315 178.58 24.645 ;
      VIA 177.79 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 24.295 178.56 24.665 ;
      VIA 177.79 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 18.875 178.58 19.205 ;
      VIA 177.79 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 18.855 178.56 19.225 ;
      VIA 177.79 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 13.435 178.58 13.765 ;
      VIA 177.79 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 13.415 178.56 13.785 ;
      VIA 177.79 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 7.995 178.58 8.325 ;
      VIA 177.79 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 7.975 178.56 8.345 ;
      VIA 177.79 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 2.555 178.58 2.885 ;
      VIA 177.79 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 2.535 178.56 2.905 ;
      VIA 177.79 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 415.995 151.44 416.325 ;
      VIA 150.65 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 415.975 151.42 416.345 ;
      VIA 150.65 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 410.555 151.44 410.885 ;
      VIA 150.65 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 410.535 151.42 410.905 ;
      VIA 150.65 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 405.115 151.44 405.445 ;
      VIA 150.65 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 405.095 151.42 405.465 ;
      VIA 150.65 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 399.675 151.44 400.005 ;
      VIA 150.65 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 399.655 151.42 400.025 ;
      VIA 150.65 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 394.235 151.44 394.565 ;
      VIA 150.65 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 394.215 151.42 394.585 ;
      VIA 150.65 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 388.795 151.44 389.125 ;
      VIA 150.65 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 388.775 151.42 389.145 ;
      VIA 150.65 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 383.355 151.44 383.685 ;
      VIA 150.65 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 383.335 151.42 383.705 ;
      VIA 150.65 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 377.915 151.44 378.245 ;
      VIA 150.65 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 377.895 151.42 378.265 ;
      VIA 150.65 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 372.475 151.44 372.805 ;
      VIA 150.65 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 372.455 151.42 372.825 ;
      VIA 150.65 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 367.035 151.44 367.365 ;
      VIA 150.65 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 367.015 151.42 367.385 ;
      VIA 150.65 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 361.595 151.44 361.925 ;
      VIA 150.65 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 361.575 151.42 361.945 ;
      VIA 150.65 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 356.155 151.44 356.485 ;
      VIA 150.65 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 356.135 151.42 356.505 ;
      VIA 150.65 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 350.715 151.44 351.045 ;
      VIA 150.65 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 350.695 151.42 351.065 ;
      VIA 150.65 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 345.275 151.44 345.605 ;
      VIA 150.65 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 345.255 151.42 345.625 ;
      VIA 150.65 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 339.835 151.44 340.165 ;
      VIA 150.65 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 339.815 151.42 340.185 ;
      VIA 150.65 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 334.395 151.44 334.725 ;
      VIA 150.65 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 334.375 151.42 334.745 ;
      VIA 150.65 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 328.955 151.44 329.285 ;
      VIA 150.65 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 328.935 151.42 329.305 ;
      VIA 150.65 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 323.515 151.44 323.845 ;
      VIA 150.65 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 323.495 151.42 323.865 ;
      VIA 150.65 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 318.075 151.44 318.405 ;
      VIA 150.65 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 318.055 151.42 318.425 ;
      VIA 150.65 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 312.635 151.44 312.965 ;
      VIA 150.65 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 312.615 151.42 312.985 ;
      VIA 150.65 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 307.195 151.44 307.525 ;
      VIA 150.65 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 307.175 151.42 307.545 ;
      VIA 150.65 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 301.755 151.44 302.085 ;
      VIA 150.65 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 301.735 151.42 302.105 ;
      VIA 150.65 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 296.315 151.44 296.645 ;
      VIA 150.65 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 296.295 151.42 296.665 ;
      VIA 150.65 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 290.875 151.44 291.205 ;
      VIA 150.65 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 290.855 151.42 291.225 ;
      VIA 150.65 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 285.435 151.44 285.765 ;
      VIA 150.65 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 285.415 151.42 285.785 ;
      VIA 150.65 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 279.995 151.44 280.325 ;
      VIA 150.65 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 279.975 151.42 280.345 ;
      VIA 150.65 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 274.555 151.44 274.885 ;
      VIA 150.65 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 274.535 151.42 274.905 ;
      VIA 150.65 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 269.115 151.44 269.445 ;
      VIA 150.65 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 269.095 151.42 269.465 ;
      VIA 150.65 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 263.675 151.44 264.005 ;
      VIA 150.65 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 263.655 151.42 264.025 ;
      VIA 150.65 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 258.235 151.44 258.565 ;
      VIA 150.65 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 258.215 151.42 258.585 ;
      VIA 150.65 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 252.795 151.44 253.125 ;
      VIA 150.65 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 252.775 151.42 253.145 ;
      VIA 150.65 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 247.355 151.44 247.685 ;
      VIA 150.65 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 247.335 151.42 247.705 ;
      VIA 150.65 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 241.915 151.44 242.245 ;
      VIA 150.65 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 241.895 151.42 242.265 ;
      VIA 150.65 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 236.475 151.44 236.805 ;
      VIA 150.65 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 236.455 151.42 236.825 ;
      VIA 150.65 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 231.035 151.44 231.365 ;
      VIA 150.65 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 231.015 151.42 231.385 ;
      VIA 150.65 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 225.595 151.44 225.925 ;
      VIA 150.65 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 225.575 151.42 225.945 ;
      VIA 150.65 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 220.155 151.44 220.485 ;
      VIA 150.65 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 220.135 151.42 220.505 ;
      VIA 150.65 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 214.715 151.44 215.045 ;
      VIA 150.65 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 214.695 151.42 215.065 ;
      VIA 150.65 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 209.275 151.44 209.605 ;
      VIA 150.65 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 209.255 151.42 209.625 ;
      VIA 150.65 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 203.835 151.44 204.165 ;
      VIA 150.65 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 203.815 151.42 204.185 ;
      VIA 150.65 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 198.395 151.44 198.725 ;
      VIA 150.65 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 198.375 151.42 198.745 ;
      VIA 150.65 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 192.955 151.44 193.285 ;
      VIA 150.65 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 192.935 151.42 193.305 ;
      VIA 150.65 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 187.515 151.44 187.845 ;
      VIA 150.65 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 187.495 151.42 187.865 ;
      VIA 150.65 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 182.075 151.44 182.405 ;
      VIA 150.65 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 182.055 151.42 182.425 ;
      VIA 150.65 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 176.635 151.44 176.965 ;
      VIA 150.65 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 176.615 151.42 176.985 ;
      VIA 150.65 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 171.195 151.44 171.525 ;
      VIA 150.65 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 171.175 151.42 171.545 ;
      VIA 150.65 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 165.755 151.44 166.085 ;
      VIA 150.65 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 165.735 151.42 166.105 ;
      VIA 150.65 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 160.315 151.44 160.645 ;
      VIA 150.65 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 160.295 151.42 160.665 ;
      VIA 150.65 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 154.875 151.44 155.205 ;
      VIA 150.65 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 154.855 151.42 155.225 ;
      VIA 150.65 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 149.435 151.44 149.765 ;
      VIA 150.65 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 149.415 151.42 149.785 ;
      VIA 150.65 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 143.995 151.44 144.325 ;
      VIA 150.65 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 143.975 151.42 144.345 ;
      VIA 150.65 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 138.555 151.44 138.885 ;
      VIA 150.65 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 138.535 151.42 138.905 ;
      VIA 150.65 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 133.115 151.44 133.445 ;
      VIA 150.65 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 133.095 151.42 133.465 ;
      VIA 150.65 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 127.675 151.44 128.005 ;
      VIA 150.65 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 127.655 151.42 128.025 ;
      VIA 150.65 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 122.235 151.44 122.565 ;
      VIA 150.65 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 122.215 151.42 122.585 ;
      VIA 150.65 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 116.795 151.44 117.125 ;
      VIA 150.65 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 116.775 151.42 117.145 ;
      VIA 150.65 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 111.355 151.44 111.685 ;
      VIA 150.65 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 111.335 151.42 111.705 ;
      VIA 150.65 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 105.915 151.44 106.245 ;
      VIA 150.65 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 105.895 151.42 106.265 ;
      VIA 150.65 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 100.475 151.44 100.805 ;
      VIA 150.65 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 100.455 151.42 100.825 ;
      VIA 150.65 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 95.035 151.44 95.365 ;
      VIA 150.65 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 95.015 151.42 95.385 ;
      VIA 150.65 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 89.595 151.44 89.925 ;
      VIA 150.65 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 89.575 151.42 89.945 ;
      VIA 150.65 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 84.155 151.44 84.485 ;
      VIA 150.65 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 84.135 151.42 84.505 ;
      VIA 150.65 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 78.715 151.44 79.045 ;
      VIA 150.65 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 78.695 151.42 79.065 ;
      VIA 150.65 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 73.275 151.44 73.605 ;
      VIA 150.65 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 73.255 151.42 73.625 ;
      VIA 150.65 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 67.835 151.44 68.165 ;
      VIA 150.65 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 67.815 151.42 68.185 ;
      VIA 150.65 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 62.395 151.44 62.725 ;
      VIA 150.65 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 62.375 151.42 62.745 ;
      VIA 150.65 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 56.955 151.44 57.285 ;
      VIA 150.65 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 56.935 151.42 57.305 ;
      VIA 150.65 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 51.515 151.44 51.845 ;
      VIA 150.65 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 51.495 151.42 51.865 ;
      VIA 150.65 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 46.075 151.44 46.405 ;
      VIA 150.65 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 46.055 151.42 46.425 ;
      VIA 150.65 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 40.635 151.44 40.965 ;
      VIA 150.65 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 40.615 151.42 40.985 ;
      VIA 150.65 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 35.195 151.44 35.525 ;
      VIA 150.65 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 35.175 151.42 35.545 ;
      VIA 150.65 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 29.755 151.44 30.085 ;
      VIA 150.65 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 29.735 151.42 30.105 ;
      VIA 150.65 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 24.315 151.44 24.645 ;
      VIA 150.65 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 24.295 151.42 24.665 ;
      VIA 150.65 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 18.875 151.44 19.205 ;
      VIA 150.65 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 18.855 151.42 19.225 ;
      VIA 150.65 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 13.435 151.44 13.765 ;
      VIA 150.65 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 13.415 151.42 13.785 ;
      VIA 150.65 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 7.995 151.44 8.325 ;
      VIA 150.65 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 7.975 151.42 8.345 ;
      VIA 150.65 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 2.555 151.44 2.885 ;
      VIA 150.65 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 2.535 151.42 2.905 ;
      VIA 150.65 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 415.995 124.3 416.325 ;
      VIA 123.51 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 415.975 124.28 416.345 ;
      VIA 123.51 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 410.555 124.3 410.885 ;
      VIA 123.51 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 410.535 124.28 410.905 ;
      VIA 123.51 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 405.115 124.3 405.445 ;
      VIA 123.51 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 405.095 124.28 405.465 ;
      VIA 123.51 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 399.675 124.3 400.005 ;
      VIA 123.51 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 399.655 124.28 400.025 ;
      VIA 123.51 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 394.235 124.3 394.565 ;
      VIA 123.51 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 394.215 124.28 394.585 ;
      VIA 123.51 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 388.795 124.3 389.125 ;
      VIA 123.51 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 388.775 124.28 389.145 ;
      VIA 123.51 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 383.355 124.3 383.685 ;
      VIA 123.51 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 383.335 124.28 383.705 ;
      VIA 123.51 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 377.915 124.3 378.245 ;
      VIA 123.51 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 377.895 124.28 378.265 ;
      VIA 123.51 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 372.475 124.3 372.805 ;
      VIA 123.51 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 372.455 124.28 372.825 ;
      VIA 123.51 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 367.035 124.3 367.365 ;
      VIA 123.51 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 367.015 124.28 367.385 ;
      VIA 123.51 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 361.595 124.3 361.925 ;
      VIA 123.51 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 361.575 124.28 361.945 ;
      VIA 123.51 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 356.155 124.3 356.485 ;
      VIA 123.51 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 356.135 124.28 356.505 ;
      VIA 123.51 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 350.715 124.3 351.045 ;
      VIA 123.51 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 350.695 124.28 351.065 ;
      VIA 123.51 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 345.275 124.3 345.605 ;
      VIA 123.51 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 345.255 124.28 345.625 ;
      VIA 123.51 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 339.835 124.3 340.165 ;
      VIA 123.51 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 339.815 124.28 340.185 ;
      VIA 123.51 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 334.395 124.3 334.725 ;
      VIA 123.51 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 334.375 124.28 334.745 ;
      VIA 123.51 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 328.955 124.3 329.285 ;
      VIA 123.51 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 328.935 124.28 329.305 ;
      VIA 123.51 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 323.515 124.3 323.845 ;
      VIA 123.51 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 323.495 124.28 323.865 ;
      VIA 123.51 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 318.075 124.3 318.405 ;
      VIA 123.51 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 318.055 124.28 318.425 ;
      VIA 123.51 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 312.635 124.3 312.965 ;
      VIA 123.51 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 312.615 124.28 312.985 ;
      VIA 123.51 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 307.195 124.3 307.525 ;
      VIA 123.51 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 307.175 124.28 307.545 ;
      VIA 123.51 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 301.755 124.3 302.085 ;
      VIA 123.51 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 301.735 124.28 302.105 ;
      VIA 123.51 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 296.315 124.3 296.645 ;
      VIA 123.51 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 296.295 124.28 296.665 ;
      VIA 123.51 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 290.875 124.3 291.205 ;
      VIA 123.51 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 290.855 124.28 291.225 ;
      VIA 123.51 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 285.435 124.3 285.765 ;
      VIA 123.51 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 285.415 124.28 285.785 ;
      VIA 123.51 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 279.995 124.3 280.325 ;
      VIA 123.51 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 279.975 124.28 280.345 ;
      VIA 123.51 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 274.555 124.3 274.885 ;
      VIA 123.51 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 274.535 124.28 274.905 ;
      VIA 123.51 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 269.115 124.3 269.445 ;
      VIA 123.51 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 269.095 124.28 269.465 ;
      VIA 123.51 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 263.675 124.3 264.005 ;
      VIA 123.51 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 263.655 124.28 264.025 ;
      VIA 123.51 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 258.235 124.3 258.565 ;
      VIA 123.51 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 258.215 124.28 258.585 ;
      VIA 123.51 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 252.795 124.3 253.125 ;
      VIA 123.51 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 252.775 124.28 253.145 ;
      VIA 123.51 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 247.355 124.3 247.685 ;
      VIA 123.51 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 247.335 124.28 247.705 ;
      VIA 123.51 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 241.915 124.3 242.245 ;
      VIA 123.51 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 241.895 124.28 242.265 ;
      VIA 123.51 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 236.475 124.3 236.805 ;
      VIA 123.51 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 236.455 124.28 236.825 ;
      VIA 123.51 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 231.035 124.3 231.365 ;
      VIA 123.51 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 231.015 124.28 231.385 ;
      VIA 123.51 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 225.595 124.3 225.925 ;
      VIA 123.51 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 225.575 124.28 225.945 ;
      VIA 123.51 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 220.155 124.3 220.485 ;
      VIA 123.51 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 220.135 124.28 220.505 ;
      VIA 123.51 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 214.715 124.3 215.045 ;
      VIA 123.51 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 214.695 124.28 215.065 ;
      VIA 123.51 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 209.275 124.3 209.605 ;
      VIA 123.51 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 209.255 124.28 209.625 ;
      VIA 123.51 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 203.835 124.3 204.165 ;
      VIA 123.51 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 203.815 124.28 204.185 ;
      VIA 123.51 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 198.395 124.3 198.725 ;
      VIA 123.51 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 198.375 124.28 198.745 ;
      VIA 123.51 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 192.955 124.3 193.285 ;
      VIA 123.51 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 192.935 124.28 193.305 ;
      VIA 123.51 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 187.515 124.3 187.845 ;
      VIA 123.51 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 187.495 124.28 187.865 ;
      VIA 123.51 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 182.075 124.3 182.405 ;
      VIA 123.51 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 182.055 124.28 182.425 ;
      VIA 123.51 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 176.635 124.3 176.965 ;
      VIA 123.51 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 176.615 124.28 176.985 ;
      VIA 123.51 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 171.195 124.3 171.525 ;
      VIA 123.51 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 171.175 124.28 171.545 ;
      VIA 123.51 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 165.755 124.3 166.085 ;
      VIA 123.51 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 165.735 124.28 166.105 ;
      VIA 123.51 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 160.315 124.3 160.645 ;
      VIA 123.51 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 160.295 124.28 160.665 ;
      VIA 123.51 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 154.875 124.3 155.205 ;
      VIA 123.51 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 154.855 124.28 155.225 ;
      VIA 123.51 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 149.435 124.3 149.765 ;
      VIA 123.51 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 149.415 124.28 149.785 ;
      VIA 123.51 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 143.995 124.3 144.325 ;
      VIA 123.51 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 143.975 124.28 144.345 ;
      VIA 123.51 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 138.555 124.3 138.885 ;
      VIA 123.51 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 138.535 124.28 138.905 ;
      VIA 123.51 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 133.115 124.3 133.445 ;
      VIA 123.51 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 133.095 124.28 133.465 ;
      VIA 123.51 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 127.675 124.3 128.005 ;
      VIA 123.51 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 127.655 124.28 128.025 ;
      VIA 123.51 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 122.235 124.3 122.565 ;
      VIA 123.51 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 122.215 124.28 122.585 ;
      VIA 123.51 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 116.795 124.3 117.125 ;
      VIA 123.51 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 116.775 124.28 117.145 ;
      VIA 123.51 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 111.355 124.3 111.685 ;
      VIA 123.51 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 111.335 124.28 111.705 ;
      VIA 123.51 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 105.915 124.3 106.245 ;
      VIA 123.51 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 105.895 124.28 106.265 ;
      VIA 123.51 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 100.475 124.3 100.805 ;
      VIA 123.51 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 100.455 124.28 100.825 ;
      VIA 123.51 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 95.035 124.3 95.365 ;
      VIA 123.51 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 95.015 124.28 95.385 ;
      VIA 123.51 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 89.595 124.3 89.925 ;
      VIA 123.51 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 89.575 124.28 89.945 ;
      VIA 123.51 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 84.155 124.3 84.485 ;
      VIA 123.51 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 84.135 124.28 84.505 ;
      VIA 123.51 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 78.715 124.3 79.045 ;
      VIA 123.51 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 78.695 124.28 79.065 ;
      VIA 123.51 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 73.275 124.3 73.605 ;
      VIA 123.51 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 73.255 124.28 73.625 ;
      VIA 123.51 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 67.835 124.3 68.165 ;
      VIA 123.51 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 67.815 124.28 68.185 ;
      VIA 123.51 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 62.395 124.3 62.725 ;
      VIA 123.51 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 62.375 124.28 62.745 ;
      VIA 123.51 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 56.955 124.3 57.285 ;
      VIA 123.51 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 56.935 124.28 57.305 ;
      VIA 123.51 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 51.515 124.3 51.845 ;
      VIA 123.51 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 51.495 124.28 51.865 ;
      VIA 123.51 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 46.075 124.3 46.405 ;
      VIA 123.51 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 46.055 124.28 46.425 ;
      VIA 123.51 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 40.635 124.3 40.965 ;
      VIA 123.51 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 40.615 124.28 40.985 ;
      VIA 123.51 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 35.195 124.3 35.525 ;
      VIA 123.51 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 35.175 124.28 35.545 ;
      VIA 123.51 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 29.755 124.3 30.085 ;
      VIA 123.51 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 29.735 124.28 30.105 ;
      VIA 123.51 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 24.315 124.3 24.645 ;
      VIA 123.51 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 24.295 124.28 24.665 ;
      VIA 123.51 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 18.875 124.3 19.205 ;
      VIA 123.51 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 18.855 124.28 19.225 ;
      VIA 123.51 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 13.435 124.3 13.765 ;
      VIA 123.51 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 13.415 124.28 13.785 ;
      VIA 123.51 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 7.995 124.3 8.325 ;
      VIA 123.51 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 7.975 124.28 8.345 ;
      VIA 123.51 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 2.555 124.3 2.885 ;
      VIA 123.51 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 2.535 124.28 2.905 ;
      VIA 123.51 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 415.995 97.16 416.325 ;
      VIA 96.37 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 415.975 97.14 416.345 ;
      VIA 96.37 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 410.555 97.16 410.885 ;
      VIA 96.37 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 410.535 97.14 410.905 ;
      VIA 96.37 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 405.115 97.16 405.445 ;
      VIA 96.37 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 405.095 97.14 405.465 ;
      VIA 96.37 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 399.675 97.16 400.005 ;
      VIA 96.37 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 399.655 97.14 400.025 ;
      VIA 96.37 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 394.235 97.16 394.565 ;
      VIA 96.37 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 394.215 97.14 394.585 ;
      VIA 96.37 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 388.795 97.16 389.125 ;
      VIA 96.37 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 388.775 97.14 389.145 ;
      VIA 96.37 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 383.355 97.16 383.685 ;
      VIA 96.37 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 383.335 97.14 383.705 ;
      VIA 96.37 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 377.915 97.16 378.245 ;
      VIA 96.37 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 377.895 97.14 378.265 ;
      VIA 96.37 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 372.475 97.16 372.805 ;
      VIA 96.37 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 372.455 97.14 372.825 ;
      VIA 96.37 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 367.035 97.16 367.365 ;
      VIA 96.37 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 367.015 97.14 367.385 ;
      VIA 96.37 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 361.595 97.16 361.925 ;
      VIA 96.37 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 361.575 97.14 361.945 ;
      VIA 96.37 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 356.155 97.16 356.485 ;
      VIA 96.37 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 356.135 97.14 356.505 ;
      VIA 96.37 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 350.715 97.16 351.045 ;
      VIA 96.37 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 350.695 97.14 351.065 ;
      VIA 96.37 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 345.275 97.16 345.605 ;
      VIA 96.37 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 345.255 97.14 345.625 ;
      VIA 96.37 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 339.835 97.16 340.165 ;
      VIA 96.37 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 339.815 97.14 340.185 ;
      VIA 96.37 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 334.395 97.16 334.725 ;
      VIA 96.37 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 334.375 97.14 334.745 ;
      VIA 96.37 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 328.955 97.16 329.285 ;
      VIA 96.37 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 328.935 97.14 329.305 ;
      VIA 96.37 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 323.515 97.16 323.845 ;
      VIA 96.37 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 323.495 97.14 323.865 ;
      VIA 96.37 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 318.075 97.16 318.405 ;
      VIA 96.37 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 318.055 97.14 318.425 ;
      VIA 96.37 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 312.635 97.16 312.965 ;
      VIA 96.37 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 312.615 97.14 312.985 ;
      VIA 96.37 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 307.195 97.16 307.525 ;
      VIA 96.37 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 307.175 97.14 307.545 ;
      VIA 96.37 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 301.755 97.16 302.085 ;
      VIA 96.37 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 301.735 97.14 302.105 ;
      VIA 96.37 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 296.315 97.16 296.645 ;
      VIA 96.37 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 296.295 97.14 296.665 ;
      VIA 96.37 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 290.875 97.16 291.205 ;
      VIA 96.37 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 290.855 97.14 291.225 ;
      VIA 96.37 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 285.435 97.16 285.765 ;
      VIA 96.37 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 285.415 97.14 285.785 ;
      VIA 96.37 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 279.995 97.16 280.325 ;
      VIA 96.37 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 279.975 97.14 280.345 ;
      VIA 96.37 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 274.555 97.16 274.885 ;
      VIA 96.37 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 274.535 97.14 274.905 ;
      VIA 96.37 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 269.115 97.16 269.445 ;
      VIA 96.37 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 269.095 97.14 269.465 ;
      VIA 96.37 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 263.675 97.16 264.005 ;
      VIA 96.37 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 263.655 97.14 264.025 ;
      VIA 96.37 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 258.235 97.16 258.565 ;
      VIA 96.37 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 258.215 97.14 258.585 ;
      VIA 96.37 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 252.795 97.16 253.125 ;
      VIA 96.37 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 252.775 97.14 253.145 ;
      VIA 96.37 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 247.355 97.16 247.685 ;
      VIA 96.37 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 247.335 97.14 247.705 ;
      VIA 96.37 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 241.915 97.16 242.245 ;
      VIA 96.37 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 241.895 97.14 242.265 ;
      VIA 96.37 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 236.475 97.16 236.805 ;
      VIA 96.37 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 236.455 97.14 236.825 ;
      VIA 96.37 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 231.035 97.16 231.365 ;
      VIA 96.37 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 231.015 97.14 231.385 ;
      VIA 96.37 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 225.595 97.16 225.925 ;
      VIA 96.37 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 225.575 97.14 225.945 ;
      VIA 96.37 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 220.155 97.16 220.485 ;
      VIA 96.37 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 220.135 97.14 220.505 ;
      VIA 96.37 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 214.715 97.16 215.045 ;
      VIA 96.37 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 214.695 97.14 215.065 ;
      VIA 96.37 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 209.275 97.16 209.605 ;
      VIA 96.37 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 209.255 97.14 209.625 ;
      VIA 96.37 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 203.835 97.16 204.165 ;
      VIA 96.37 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 203.815 97.14 204.185 ;
      VIA 96.37 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 198.395 97.16 198.725 ;
      VIA 96.37 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 198.375 97.14 198.745 ;
      VIA 96.37 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 192.955 97.16 193.285 ;
      VIA 96.37 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 192.935 97.14 193.305 ;
      VIA 96.37 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 187.515 97.16 187.845 ;
      VIA 96.37 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 187.495 97.14 187.865 ;
      VIA 96.37 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 182.075 97.16 182.405 ;
      VIA 96.37 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 182.055 97.14 182.425 ;
      VIA 96.37 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 176.635 97.16 176.965 ;
      VIA 96.37 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 176.615 97.14 176.985 ;
      VIA 96.37 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 171.195 97.16 171.525 ;
      VIA 96.37 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 171.175 97.14 171.545 ;
      VIA 96.37 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 165.755 97.16 166.085 ;
      VIA 96.37 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 165.735 97.14 166.105 ;
      VIA 96.37 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 160.315 97.16 160.645 ;
      VIA 96.37 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 160.295 97.14 160.665 ;
      VIA 96.37 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 154.875 97.16 155.205 ;
      VIA 96.37 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 154.855 97.14 155.225 ;
      VIA 96.37 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 149.435 97.16 149.765 ;
      VIA 96.37 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 149.415 97.14 149.785 ;
      VIA 96.37 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 143.995 97.16 144.325 ;
      VIA 96.37 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 143.975 97.14 144.345 ;
      VIA 96.37 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 138.555 97.16 138.885 ;
      VIA 96.37 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 138.535 97.14 138.905 ;
      VIA 96.37 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 133.115 97.16 133.445 ;
      VIA 96.37 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 133.095 97.14 133.465 ;
      VIA 96.37 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 127.675 97.16 128.005 ;
      VIA 96.37 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 127.655 97.14 128.025 ;
      VIA 96.37 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 122.235 97.16 122.565 ;
      VIA 96.37 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 122.215 97.14 122.585 ;
      VIA 96.37 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 116.795 97.16 117.125 ;
      VIA 96.37 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 116.775 97.14 117.145 ;
      VIA 96.37 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 111.355 97.16 111.685 ;
      VIA 96.37 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 111.335 97.14 111.705 ;
      VIA 96.37 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 105.915 97.16 106.245 ;
      VIA 96.37 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 105.895 97.14 106.265 ;
      VIA 96.37 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 100.475 97.16 100.805 ;
      VIA 96.37 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 100.455 97.14 100.825 ;
      VIA 96.37 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 95.035 97.16 95.365 ;
      VIA 96.37 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 95.015 97.14 95.385 ;
      VIA 96.37 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 89.595 97.16 89.925 ;
      VIA 96.37 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 89.575 97.14 89.945 ;
      VIA 96.37 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 84.155 97.16 84.485 ;
      VIA 96.37 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 84.135 97.14 84.505 ;
      VIA 96.37 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 78.715 97.16 79.045 ;
      VIA 96.37 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 78.695 97.14 79.065 ;
      VIA 96.37 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 73.275 97.16 73.605 ;
      VIA 96.37 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 73.255 97.14 73.625 ;
      VIA 96.37 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 67.835 97.16 68.165 ;
      VIA 96.37 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 67.815 97.14 68.185 ;
      VIA 96.37 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 62.395 97.16 62.725 ;
      VIA 96.37 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 62.375 97.14 62.745 ;
      VIA 96.37 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 56.955 97.16 57.285 ;
      VIA 96.37 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 56.935 97.14 57.305 ;
      VIA 96.37 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 51.515 97.16 51.845 ;
      VIA 96.37 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 51.495 97.14 51.865 ;
      VIA 96.37 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 46.075 97.16 46.405 ;
      VIA 96.37 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 46.055 97.14 46.425 ;
      VIA 96.37 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 40.635 97.16 40.965 ;
      VIA 96.37 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 40.615 97.14 40.985 ;
      VIA 96.37 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 35.195 97.16 35.525 ;
      VIA 96.37 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 35.175 97.14 35.545 ;
      VIA 96.37 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 29.755 97.16 30.085 ;
      VIA 96.37 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 29.735 97.14 30.105 ;
      VIA 96.37 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 24.315 97.16 24.645 ;
      VIA 96.37 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 24.295 97.14 24.665 ;
      VIA 96.37 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 18.875 97.16 19.205 ;
      VIA 96.37 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 18.855 97.14 19.225 ;
      VIA 96.37 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 13.435 97.16 13.765 ;
      VIA 96.37 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 13.415 97.14 13.785 ;
      VIA 96.37 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 7.995 97.16 8.325 ;
      VIA 96.37 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 7.975 97.14 8.345 ;
      VIA 96.37 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 2.555 97.16 2.885 ;
      VIA 96.37 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 2.535 97.14 2.905 ;
      VIA 96.37 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 415.995 70.02 416.325 ;
      VIA 69.23 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 415.975 70 416.345 ;
      VIA 69.23 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 410.555 70.02 410.885 ;
      VIA 69.23 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 410.535 70 410.905 ;
      VIA 69.23 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 405.115 70.02 405.445 ;
      VIA 69.23 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 405.095 70 405.465 ;
      VIA 69.23 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 399.675 70.02 400.005 ;
      VIA 69.23 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 399.655 70 400.025 ;
      VIA 69.23 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 394.235 70.02 394.565 ;
      VIA 69.23 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 394.215 70 394.585 ;
      VIA 69.23 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 388.795 70.02 389.125 ;
      VIA 69.23 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 388.775 70 389.145 ;
      VIA 69.23 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 383.355 70.02 383.685 ;
      VIA 69.23 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 383.335 70 383.705 ;
      VIA 69.23 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 377.915 70.02 378.245 ;
      VIA 69.23 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 377.895 70 378.265 ;
      VIA 69.23 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 372.475 70.02 372.805 ;
      VIA 69.23 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 372.455 70 372.825 ;
      VIA 69.23 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 367.035 70.02 367.365 ;
      VIA 69.23 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 367.015 70 367.385 ;
      VIA 69.23 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 361.595 70.02 361.925 ;
      VIA 69.23 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 361.575 70 361.945 ;
      VIA 69.23 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 356.155 70.02 356.485 ;
      VIA 69.23 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 356.135 70 356.505 ;
      VIA 69.23 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 350.715 70.02 351.045 ;
      VIA 69.23 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 350.695 70 351.065 ;
      VIA 69.23 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 345.275 70.02 345.605 ;
      VIA 69.23 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 345.255 70 345.625 ;
      VIA 69.23 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 339.835 70.02 340.165 ;
      VIA 69.23 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 339.815 70 340.185 ;
      VIA 69.23 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 334.395 70.02 334.725 ;
      VIA 69.23 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 334.375 70 334.745 ;
      VIA 69.23 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 328.955 70.02 329.285 ;
      VIA 69.23 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 328.935 70 329.305 ;
      VIA 69.23 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 323.515 70.02 323.845 ;
      VIA 69.23 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 323.495 70 323.865 ;
      VIA 69.23 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 318.075 70.02 318.405 ;
      VIA 69.23 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 318.055 70 318.425 ;
      VIA 69.23 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 312.635 70.02 312.965 ;
      VIA 69.23 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 312.615 70 312.985 ;
      VIA 69.23 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 307.195 70.02 307.525 ;
      VIA 69.23 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 307.175 70 307.545 ;
      VIA 69.23 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 301.755 70.02 302.085 ;
      VIA 69.23 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 301.735 70 302.105 ;
      VIA 69.23 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 296.315 70.02 296.645 ;
      VIA 69.23 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 296.295 70 296.665 ;
      VIA 69.23 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 290.875 70.02 291.205 ;
      VIA 69.23 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 290.855 70 291.225 ;
      VIA 69.23 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 285.435 70.02 285.765 ;
      VIA 69.23 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 285.415 70 285.785 ;
      VIA 69.23 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 279.995 70.02 280.325 ;
      VIA 69.23 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 279.975 70 280.345 ;
      VIA 69.23 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 274.555 70.02 274.885 ;
      VIA 69.23 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 274.535 70 274.905 ;
      VIA 69.23 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 269.115 70.02 269.445 ;
      VIA 69.23 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 269.095 70 269.465 ;
      VIA 69.23 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 263.675 70.02 264.005 ;
      VIA 69.23 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 263.655 70 264.025 ;
      VIA 69.23 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 258.235 70.02 258.565 ;
      VIA 69.23 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 258.215 70 258.585 ;
      VIA 69.23 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 252.795 70.02 253.125 ;
      VIA 69.23 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 252.775 70 253.145 ;
      VIA 69.23 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 247.355 70.02 247.685 ;
      VIA 69.23 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 247.335 70 247.705 ;
      VIA 69.23 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 241.915 70.02 242.245 ;
      VIA 69.23 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 241.895 70 242.265 ;
      VIA 69.23 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 236.475 70.02 236.805 ;
      VIA 69.23 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 236.455 70 236.825 ;
      VIA 69.23 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 231.035 70.02 231.365 ;
      VIA 69.23 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 231.015 70 231.385 ;
      VIA 69.23 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 225.595 70.02 225.925 ;
      VIA 69.23 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 225.575 70 225.945 ;
      VIA 69.23 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 220.155 70.02 220.485 ;
      VIA 69.23 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 220.135 70 220.505 ;
      VIA 69.23 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 214.715 70.02 215.045 ;
      VIA 69.23 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 214.695 70 215.065 ;
      VIA 69.23 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 209.275 70.02 209.605 ;
      VIA 69.23 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 209.255 70 209.625 ;
      VIA 69.23 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 203.835 70.02 204.165 ;
      VIA 69.23 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 203.815 70 204.185 ;
      VIA 69.23 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 198.395 70.02 198.725 ;
      VIA 69.23 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 198.375 70 198.745 ;
      VIA 69.23 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 192.955 70.02 193.285 ;
      VIA 69.23 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 192.935 70 193.305 ;
      VIA 69.23 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 187.515 70.02 187.845 ;
      VIA 69.23 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 187.495 70 187.865 ;
      VIA 69.23 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 182.075 70.02 182.405 ;
      VIA 69.23 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 182.055 70 182.425 ;
      VIA 69.23 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 176.635 70.02 176.965 ;
      VIA 69.23 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 176.615 70 176.985 ;
      VIA 69.23 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 171.195 70.02 171.525 ;
      VIA 69.23 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 171.175 70 171.545 ;
      VIA 69.23 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 165.755 70.02 166.085 ;
      VIA 69.23 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 165.735 70 166.105 ;
      VIA 69.23 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 160.315 70.02 160.645 ;
      VIA 69.23 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 160.295 70 160.665 ;
      VIA 69.23 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 154.875 70.02 155.205 ;
      VIA 69.23 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 154.855 70 155.225 ;
      VIA 69.23 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 149.435 70.02 149.765 ;
      VIA 69.23 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 149.415 70 149.785 ;
      VIA 69.23 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 143.995 70.02 144.325 ;
      VIA 69.23 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 143.975 70 144.345 ;
      VIA 69.23 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 138.555 70.02 138.885 ;
      VIA 69.23 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 138.535 70 138.905 ;
      VIA 69.23 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 133.115 70.02 133.445 ;
      VIA 69.23 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 133.095 70 133.465 ;
      VIA 69.23 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 127.675 70.02 128.005 ;
      VIA 69.23 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 127.655 70 128.025 ;
      VIA 69.23 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 122.235 70.02 122.565 ;
      VIA 69.23 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 122.215 70 122.585 ;
      VIA 69.23 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 116.795 70.02 117.125 ;
      VIA 69.23 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 116.775 70 117.145 ;
      VIA 69.23 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 111.355 70.02 111.685 ;
      VIA 69.23 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 111.335 70 111.705 ;
      VIA 69.23 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 105.915 70.02 106.245 ;
      VIA 69.23 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 105.895 70 106.265 ;
      VIA 69.23 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 100.475 70.02 100.805 ;
      VIA 69.23 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 100.455 70 100.825 ;
      VIA 69.23 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 95.035 70.02 95.365 ;
      VIA 69.23 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 95.015 70 95.385 ;
      VIA 69.23 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 89.595 70.02 89.925 ;
      VIA 69.23 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 89.575 70 89.945 ;
      VIA 69.23 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 84.155 70.02 84.485 ;
      VIA 69.23 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 84.135 70 84.505 ;
      VIA 69.23 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 78.715 70.02 79.045 ;
      VIA 69.23 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 78.695 70 79.065 ;
      VIA 69.23 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 73.275 70.02 73.605 ;
      VIA 69.23 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 73.255 70 73.625 ;
      VIA 69.23 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 67.835 70.02 68.165 ;
      VIA 69.23 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 67.815 70 68.185 ;
      VIA 69.23 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 62.395 70.02 62.725 ;
      VIA 69.23 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 62.375 70 62.745 ;
      VIA 69.23 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 56.955 70.02 57.285 ;
      VIA 69.23 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 56.935 70 57.305 ;
      VIA 69.23 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 51.515 70.02 51.845 ;
      VIA 69.23 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 51.495 70 51.865 ;
      VIA 69.23 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 46.075 70.02 46.405 ;
      VIA 69.23 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 46.055 70 46.425 ;
      VIA 69.23 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 40.635 70.02 40.965 ;
      VIA 69.23 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 40.615 70 40.985 ;
      VIA 69.23 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 35.195 70.02 35.525 ;
      VIA 69.23 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 35.175 70 35.545 ;
      VIA 69.23 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 29.755 70.02 30.085 ;
      VIA 69.23 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 29.735 70 30.105 ;
      VIA 69.23 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 24.315 70.02 24.645 ;
      VIA 69.23 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 24.295 70 24.665 ;
      VIA 69.23 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 18.875 70.02 19.205 ;
      VIA 69.23 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 18.855 70 19.225 ;
      VIA 69.23 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 13.435 70.02 13.765 ;
      VIA 69.23 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 13.415 70 13.785 ;
      VIA 69.23 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 7.995 70.02 8.325 ;
      VIA 69.23 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 7.975 70 8.345 ;
      VIA 69.23 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 2.555 70.02 2.885 ;
      VIA 69.23 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 2.535 70 2.905 ;
      VIA 69.23 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 415.995 42.88 416.325 ;
      VIA 42.09 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 415.975 42.86 416.345 ;
      VIA 42.09 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 410.555 42.88 410.885 ;
      VIA 42.09 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 410.535 42.86 410.905 ;
      VIA 42.09 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 405.115 42.88 405.445 ;
      VIA 42.09 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 405.095 42.86 405.465 ;
      VIA 42.09 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 399.675 42.88 400.005 ;
      VIA 42.09 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 399.655 42.86 400.025 ;
      VIA 42.09 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 394.235 42.88 394.565 ;
      VIA 42.09 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 394.215 42.86 394.585 ;
      VIA 42.09 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 388.795 42.88 389.125 ;
      VIA 42.09 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 388.775 42.86 389.145 ;
      VIA 42.09 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 383.355 42.88 383.685 ;
      VIA 42.09 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 383.335 42.86 383.705 ;
      VIA 42.09 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 377.915 42.88 378.245 ;
      VIA 42.09 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 377.895 42.86 378.265 ;
      VIA 42.09 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 372.475 42.88 372.805 ;
      VIA 42.09 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 372.455 42.86 372.825 ;
      VIA 42.09 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 367.035 42.88 367.365 ;
      VIA 42.09 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 367.015 42.86 367.385 ;
      VIA 42.09 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 361.595 42.88 361.925 ;
      VIA 42.09 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 361.575 42.86 361.945 ;
      VIA 42.09 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 356.155 42.88 356.485 ;
      VIA 42.09 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 356.135 42.86 356.505 ;
      VIA 42.09 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 350.715 42.88 351.045 ;
      VIA 42.09 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 350.695 42.86 351.065 ;
      VIA 42.09 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 345.275 42.88 345.605 ;
      VIA 42.09 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 345.255 42.86 345.625 ;
      VIA 42.09 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 339.835 42.88 340.165 ;
      VIA 42.09 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 339.815 42.86 340.185 ;
      VIA 42.09 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 334.395 42.88 334.725 ;
      VIA 42.09 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 334.375 42.86 334.745 ;
      VIA 42.09 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 328.955 42.88 329.285 ;
      VIA 42.09 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 328.935 42.86 329.305 ;
      VIA 42.09 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 323.515 42.88 323.845 ;
      VIA 42.09 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 323.495 42.86 323.865 ;
      VIA 42.09 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 318.075 42.88 318.405 ;
      VIA 42.09 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 318.055 42.86 318.425 ;
      VIA 42.09 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 312.635 42.88 312.965 ;
      VIA 42.09 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 312.615 42.86 312.985 ;
      VIA 42.09 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 307.195 42.88 307.525 ;
      VIA 42.09 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 307.175 42.86 307.545 ;
      VIA 42.09 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 301.755 42.88 302.085 ;
      VIA 42.09 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 301.735 42.86 302.105 ;
      VIA 42.09 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 296.315 42.88 296.645 ;
      VIA 42.09 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 296.295 42.86 296.665 ;
      VIA 42.09 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 290.875 42.88 291.205 ;
      VIA 42.09 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 290.855 42.86 291.225 ;
      VIA 42.09 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 285.435 42.88 285.765 ;
      VIA 42.09 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 285.415 42.86 285.785 ;
      VIA 42.09 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 279.995 42.88 280.325 ;
      VIA 42.09 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 279.975 42.86 280.345 ;
      VIA 42.09 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 274.555 42.88 274.885 ;
      VIA 42.09 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 274.535 42.86 274.905 ;
      VIA 42.09 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 269.115 42.88 269.445 ;
      VIA 42.09 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 269.095 42.86 269.465 ;
      VIA 42.09 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 263.675 42.88 264.005 ;
      VIA 42.09 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 263.655 42.86 264.025 ;
      VIA 42.09 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 258.235 42.88 258.565 ;
      VIA 42.09 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 258.215 42.86 258.585 ;
      VIA 42.09 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 252.795 42.88 253.125 ;
      VIA 42.09 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 252.775 42.86 253.145 ;
      VIA 42.09 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 247.355 42.88 247.685 ;
      VIA 42.09 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 247.335 42.86 247.705 ;
      VIA 42.09 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 241.915 42.88 242.245 ;
      VIA 42.09 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 241.895 42.86 242.265 ;
      VIA 42.09 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 236.475 42.88 236.805 ;
      VIA 42.09 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 236.455 42.86 236.825 ;
      VIA 42.09 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 231.035 42.88 231.365 ;
      VIA 42.09 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 231.015 42.86 231.385 ;
      VIA 42.09 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 225.595 42.88 225.925 ;
      VIA 42.09 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 225.575 42.86 225.945 ;
      VIA 42.09 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 220.155 42.88 220.485 ;
      VIA 42.09 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 220.135 42.86 220.505 ;
      VIA 42.09 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 214.715 42.88 215.045 ;
      VIA 42.09 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 214.695 42.86 215.065 ;
      VIA 42.09 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 209.275 42.88 209.605 ;
      VIA 42.09 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 209.255 42.86 209.625 ;
      VIA 42.09 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 203.835 42.88 204.165 ;
      VIA 42.09 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 203.815 42.86 204.185 ;
      VIA 42.09 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 198.395 42.88 198.725 ;
      VIA 42.09 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 198.375 42.86 198.745 ;
      VIA 42.09 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 192.955 42.88 193.285 ;
      VIA 42.09 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 192.935 42.86 193.305 ;
      VIA 42.09 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 187.515 42.88 187.845 ;
      VIA 42.09 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 187.495 42.86 187.865 ;
      VIA 42.09 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 182.075 42.88 182.405 ;
      VIA 42.09 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 182.055 42.86 182.425 ;
      VIA 42.09 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 176.635 42.88 176.965 ;
      VIA 42.09 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 176.615 42.86 176.985 ;
      VIA 42.09 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 171.195 42.88 171.525 ;
      VIA 42.09 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 171.175 42.86 171.545 ;
      VIA 42.09 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 165.755 42.88 166.085 ;
      VIA 42.09 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 165.735 42.86 166.105 ;
      VIA 42.09 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 160.315 42.88 160.645 ;
      VIA 42.09 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 160.295 42.86 160.665 ;
      VIA 42.09 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 154.875 42.88 155.205 ;
      VIA 42.09 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 154.855 42.86 155.225 ;
      VIA 42.09 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 149.435 42.88 149.765 ;
      VIA 42.09 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 149.415 42.86 149.785 ;
      VIA 42.09 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 143.995 42.88 144.325 ;
      VIA 42.09 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 143.975 42.86 144.345 ;
      VIA 42.09 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 138.555 42.88 138.885 ;
      VIA 42.09 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 138.535 42.86 138.905 ;
      VIA 42.09 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 133.115 42.88 133.445 ;
      VIA 42.09 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 133.095 42.86 133.465 ;
      VIA 42.09 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 127.675 42.88 128.005 ;
      VIA 42.09 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 127.655 42.86 128.025 ;
      VIA 42.09 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 122.235 42.88 122.565 ;
      VIA 42.09 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 122.215 42.86 122.585 ;
      VIA 42.09 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 116.795 42.88 117.125 ;
      VIA 42.09 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 116.775 42.86 117.145 ;
      VIA 42.09 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 111.355 42.88 111.685 ;
      VIA 42.09 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 111.335 42.86 111.705 ;
      VIA 42.09 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 105.915 42.88 106.245 ;
      VIA 42.09 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 105.895 42.86 106.265 ;
      VIA 42.09 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 100.475 42.88 100.805 ;
      VIA 42.09 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 100.455 42.86 100.825 ;
      VIA 42.09 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 95.035 42.88 95.365 ;
      VIA 42.09 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 95.015 42.86 95.385 ;
      VIA 42.09 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 89.595 42.88 89.925 ;
      VIA 42.09 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 89.575 42.86 89.945 ;
      VIA 42.09 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 84.155 42.88 84.485 ;
      VIA 42.09 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 84.135 42.86 84.505 ;
      VIA 42.09 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 78.715 42.88 79.045 ;
      VIA 42.09 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 78.695 42.86 79.065 ;
      VIA 42.09 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 73.275 42.88 73.605 ;
      VIA 42.09 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 73.255 42.86 73.625 ;
      VIA 42.09 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 67.835 42.88 68.165 ;
      VIA 42.09 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 67.815 42.86 68.185 ;
      VIA 42.09 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 62.395 42.88 62.725 ;
      VIA 42.09 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 62.375 42.86 62.745 ;
      VIA 42.09 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 56.955 42.88 57.285 ;
      VIA 42.09 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 56.935 42.86 57.305 ;
      VIA 42.09 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 51.515 42.88 51.845 ;
      VIA 42.09 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 51.495 42.86 51.865 ;
      VIA 42.09 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 46.075 42.88 46.405 ;
      VIA 42.09 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 46.055 42.86 46.425 ;
      VIA 42.09 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 40.635 42.88 40.965 ;
      VIA 42.09 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 40.615 42.86 40.985 ;
      VIA 42.09 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 35.195 42.88 35.525 ;
      VIA 42.09 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 35.175 42.86 35.545 ;
      VIA 42.09 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 29.755 42.88 30.085 ;
      VIA 42.09 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 29.735 42.86 30.105 ;
      VIA 42.09 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 24.315 42.88 24.645 ;
      VIA 42.09 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 24.295 42.86 24.665 ;
      VIA 42.09 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 18.875 42.88 19.205 ;
      VIA 42.09 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 18.855 42.86 19.225 ;
      VIA 42.09 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 13.435 42.88 13.765 ;
      VIA 42.09 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 13.415 42.86 13.785 ;
      VIA 42.09 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 7.995 42.88 8.325 ;
      VIA 42.09 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 7.975 42.86 8.345 ;
      VIA 42.09 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 2.555 42.88 2.885 ;
      VIA 42.09 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 2.535 42.86 2.905 ;
      VIA 42.09 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 415.995 15.74 416.325 ;
      VIA 14.95 416.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 415.975 15.72 416.345 ;
      VIA 14.95 416.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 416.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 410.555 15.74 410.885 ;
      VIA 14.95 410.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 410.535 15.72 410.905 ;
      VIA 14.95 410.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 410.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 405.115 15.74 405.445 ;
      VIA 14.95 405.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 405.095 15.72 405.465 ;
      VIA 14.95 405.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 405.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 399.675 15.74 400.005 ;
      VIA 14.95 399.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 399.655 15.72 400.025 ;
      VIA 14.95 399.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 399.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 394.235 15.74 394.565 ;
      VIA 14.95 394.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 394.215 15.72 394.585 ;
      VIA 14.95 394.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 394.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 388.795 15.74 389.125 ;
      VIA 14.95 388.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 388.775 15.72 389.145 ;
      VIA 14.95 388.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 388.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 383.355 15.74 383.685 ;
      VIA 14.95 383.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 383.335 15.72 383.705 ;
      VIA 14.95 383.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 383.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 377.915 15.74 378.245 ;
      VIA 14.95 378.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 377.895 15.72 378.265 ;
      VIA 14.95 378.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 378.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 372.475 15.74 372.805 ;
      VIA 14.95 372.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 372.455 15.72 372.825 ;
      VIA 14.95 372.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 372.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 367.035 15.74 367.365 ;
      VIA 14.95 367.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 367.015 15.72 367.385 ;
      VIA 14.95 367.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 367.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 361.595 15.74 361.925 ;
      VIA 14.95 361.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 361.575 15.72 361.945 ;
      VIA 14.95 361.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 361.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 356.155 15.74 356.485 ;
      VIA 14.95 356.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 356.135 15.72 356.505 ;
      VIA 14.95 356.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 356.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 350.715 15.74 351.045 ;
      VIA 14.95 350.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 350.695 15.72 351.065 ;
      VIA 14.95 350.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 350.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 345.275 15.74 345.605 ;
      VIA 14.95 345.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 345.255 15.72 345.625 ;
      VIA 14.95 345.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 345.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 339.835 15.74 340.165 ;
      VIA 14.95 340 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 339.815 15.72 340.185 ;
      VIA 14.95 340 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 340 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 334.395 15.74 334.725 ;
      VIA 14.95 334.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 334.375 15.72 334.745 ;
      VIA 14.95 334.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 334.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 328.955 15.74 329.285 ;
      VIA 14.95 329.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 328.935 15.72 329.305 ;
      VIA 14.95 329.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 329.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 323.515 15.74 323.845 ;
      VIA 14.95 323.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 323.495 15.72 323.865 ;
      VIA 14.95 323.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 323.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 318.075 15.74 318.405 ;
      VIA 14.95 318.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 318.055 15.72 318.425 ;
      VIA 14.95 318.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 318.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 312.635 15.74 312.965 ;
      VIA 14.95 312.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 312.615 15.72 312.985 ;
      VIA 14.95 312.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 312.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 307.195 15.74 307.525 ;
      VIA 14.95 307.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 307.175 15.72 307.545 ;
      VIA 14.95 307.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 307.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 301.755 15.74 302.085 ;
      VIA 14.95 301.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 301.735 15.72 302.105 ;
      VIA 14.95 301.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 301.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 296.315 15.74 296.645 ;
      VIA 14.95 296.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 296.295 15.72 296.665 ;
      VIA 14.95 296.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 296.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 290.875 15.74 291.205 ;
      VIA 14.95 291.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 290.855 15.72 291.225 ;
      VIA 14.95 291.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 291.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 285.435 15.74 285.765 ;
      VIA 14.95 285.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 285.415 15.72 285.785 ;
      VIA 14.95 285.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 285.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 279.995 15.74 280.325 ;
      VIA 14.95 280.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 279.975 15.72 280.345 ;
      VIA 14.95 280.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 280.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 274.555 15.74 274.885 ;
      VIA 14.95 274.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 274.535 15.72 274.905 ;
      VIA 14.95 274.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 274.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 269.115 15.74 269.445 ;
      VIA 14.95 269.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 269.095 15.72 269.465 ;
      VIA 14.95 269.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 269.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 263.675 15.74 264.005 ;
      VIA 14.95 263.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 263.655 15.72 264.025 ;
      VIA 14.95 263.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 263.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 258.235 15.74 258.565 ;
      VIA 14.95 258.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 258.215 15.72 258.585 ;
      VIA 14.95 258.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 258.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 252.795 15.74 253.125 ;
      VIA 14.95 252.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 252.775 15.72 253.145 ;
      VIA 14.95 252.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 252.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 247.355 15.74 247.685 ;
      VIA 14.95 247.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 247.335 15.72 247.705 ;
      VIA 14.95 247.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 247.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 241.915 15.74 242.245 ;
      VIA 14.95 242.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 241.895 15.72 242.265 ;
      VIA 14.95 242.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 242.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 236.475 15.74 236.805 ;
      VIA 14.95 236.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 236.455 15.72 236.825 ;
      VIA 14.95 236.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 236.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 231.035 15.74 231.365 ;
      VIA 14.95 231.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 231.015 15.72 231.385 ;
      VIA 14.95 231.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 231.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 225.595 15.74 225.925 ;
      VIA 14.95 225.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 225.575 15.72 225.945 ;
      VIA 14.95 225.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 225.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 220.155 15.74 220.485 ;
      VIA 14.95 220.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 220.135 15.72 220.505 ;
      VIA 14.95 220.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 220.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 214.715 15.74 215.045 ;
      VIA 14.95 214.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 214.695 15.72 215.065 ;
      VIA 14.95 214.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 214.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 209.275 15.74 209.605 ;
      VIA 14.95 209.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 209.255 15.72 209.625 ;
      VIA 14.95 209.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 209.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 203.835 15.74 204.165 ;
      VIA 14.95 204 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 203.815 15.72 204.185 ;
      VIA 14.95 204 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 204 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 198.395 15.74 198.725 ;
      VIA 14.95 198.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 198.375 15.72 198.745 ;
      VIA 14.95 198.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 198.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 192.955 15.74 193.285 ;
      VIA 14.95 193.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 192.935 15.72 193.305 ;
      VIA 14.95 193.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 193.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 187.515 15.74 187.845 ;
      VIA 14.95 187.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 187.495 15.72 187.865 ;
      VIA 14.95 187.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 187.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 182.075 15.74 182.405 ;
      VIA 14.95 182.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 182.055 15.72 182.425 ;
      VIA 14.95 182.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 182.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 176.635 15.74 176.965 ;
      VIA 14.95 176.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 176.615 15.72 176.985 ;
      VIA 14.95 176.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 176.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 171.195 15.74 171.525 ;
      VIA 14.95 171.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 171.175 15.72 171.545 ;
      VIA 14.95 171.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 171.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 165.755 15.74 166.085 ;
      VIA 14.95 165.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 165.735 15.72 166.105 ;
      VIA 14.95 165.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 165.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 160.315 15.74 160.645 ;
      VIA 14.95 160.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 160.295 15.72 160.665 ;
      VIA 14.95 160.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 160.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 154.875 15.74 155.205 ;
      VIA 14.95 155.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 154.855 15.72 155.225 ;
      VIA 14.95 155.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 155.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 149.435 15.74 149.765 ;
      VIA 14.95 149.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 149.415 15.72 149.785 ;
      VIA 14.95 149.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 149.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 143.995 15.74 144.325 ;
      VIA 14.95 144.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 143.975 15.72 144.345 ;
      VIA 14.95 144.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 144.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 138.555 15.74 138.885 ;
      VIA 14.95 138.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 138.535 15.72 138.905 ;
      VIA 14.95 138.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 138.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 133.115 15.74 133.445 ;
      VIA 14.95 133.28 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 133.095 15.72 133.465 ;
      VIA 14.95 133.28 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 133.28 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 127.675 15.74 128.005 ;
      VIA 14.95 127.84 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 127.655 15.72 128.025 ;
      VIA 14.95 127.84 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 127.84 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 122.235 15.74 122.565 ;
      VIA 14.95 122.4 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 122.215 15.72 122.585 ;
      VIA 14.95 122.4 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 122.4 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 116.795 15.74 117.125 ;
      VIA 14.95 116.96 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 116.775 15.72 117.145 ;
      VIA 14.95 116.96 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 116.96 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 111.355 15.74 111.685 ;
      VIA 14.95 111.52 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 111.335 15.72 111.705 ;
      VIA 14.95 111.52 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 111.52 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 105.915 15.74 106.245 ;
      VIA 14.95 106.08 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 105.895 15.72 106.265 ;
      VIA 14.95 106.08 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 106.08 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 100.475 15.74 100.805 ;
      VIA 14.95 100.64 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 100.455 15.72 100.825 ;
      VIA 14.95 100.64 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 100.64 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 95.035 15.74 95.365 ;
      VIA 14.95 95.2 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 95.015 15.72 95.385 ;
      VIA 14.95 95.2 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 95.2 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 89.595 15.74 89.925 ;
      VIA 14.95 89.76 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 89.575 15.72 89.945 ;
      VIA 14.95 89.76 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 89.76 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 84.155 15.74 84.485 ;
      VIA 14.95 84.32 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 84.135 15.72 84.505 ;
      VIA 14.95 84.32 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 84.32 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 78.715 15.74 79.045 ;
      VIA 14.95 78.88 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 78.695 15.72 79.065 ;
      VIA 14.95 78.88 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 78.88 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 73.275 15.74 73.605 ;
      VIA 14.95 73.44 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 73.255 15.72 73.625 ;
      VIA 14.95 73.44 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 73.44 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 67.835 15.74 68.165 ;
      VIA 14.95 68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 67.815 15.72 68.185 ;
      VIA 14.95 68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 62.395 15.74 62.725 ;
      VIA 14.95 62.56 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 62.375 15.72 62.745 ;
      VIA 14.95 62.56 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 62.56 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 56.955 15.74 57.285 ;
      VIA 14.95 57.12 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 56.935 15.72 57.305 ;
      VIA 14.95 57.12 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 57.12 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 51.515 15.74 51.845 ;
      VIA 14.95 51.68 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 51.495 15.72 51.865 ;
      VIA 14.95 51.68 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 51.68 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 46.075 15.74 46.405 ;
      VIA 14.95 46.24 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 46.055 15.72 46.425 ;
      VIA 14.95 46.24 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 46.24 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 40.635 15.74 40.965 ;
      VIA 14.95 40.8 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 40.615 15.72 40.985 ;
      VIA 14.95 40.8 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 40.8 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 35.195 15.74 35.525 ;
      VIA 14.95 35.36 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 35.175 15.72 35.545 ;
      VIA 14.95 35.36 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 35.36 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 29.755 15.74 30.085 ;
      VIA 14.95 29.92 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 29.735 15.72 30.105 ;
      VIA 14.95 29.92 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 29.92 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 24.315 15.74 24.645 ;
      VIA 14.95 24.48 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 24.295 15.72 24.665 ;
      VIA 14.95 24.48 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 24.48 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 18.875 15.74 19.205 ;
      VIA 14.95 19.04 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 18.855 15.72 19.225 ;
      VIA 14.95 19.04 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 19.04 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 13.435 15.74 13.765 ;
      VIA 14.95 13.6 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 13.415 15.72 13.785 ;
      VIA 14.95 13.6 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 13.6 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 7.995 15.74 8.325 ;
      VIA 14.95 8.16 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 7.975 15.72 8.345 ;
      VIA 14.95 8.16 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 8.16 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 2.555 15.74 2.885 ;
      VIA 14.95 2.72 ibex_register_file_ff_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 2.535 15.72 2.905 ;
      VIA 14.95 2.72 ibex_register_file_ff_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 2.72 ibex_register_file_ff_via2_3_1600_480_1_5_320_320 ;
    END
  END VSS
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 412.27 0.8 412.57 ;
    END
  END clk_i
  PIN dummy_instr_id_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  4.3 0 4.44 0.485 ;
    END
  END dummy_instr_id_i
  PIN raddr_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  215.44 0 215.58 0.485 ;
    END
  END raddr_a_i[0]
  PIN raddr_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  219.58 0 219.72 0.485 ;
    END
  END raddr_a_i[1]
  PIN raddr_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 171.55 421.97 171.85 ;
    END
  END raddr_a_i[2]
  PIN raddr_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  211.3 0 211.44 0.485 ;
    END
  END raddr_a_i[3]
  PIN raddr_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  277.54 0 277.68 0.485 ;
    END
  END raddr_a_i[4]
  PIN raddr_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  182.32 0 182.46 0.485 ;
    END
  END raddr_b_i[0]
  PIN raddr_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 175.63 421.97 175.93 ;
    END
  END raddr_b_i[1]
  PIN raddr_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  215.44 421.485 215.58 421.97 ;
    END
  END raddr_b_i[2]
  PIN raddr_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 179.71 421.97 180.01 ;
    END
  END raddr_b_i[3]
  PIN raddr_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 187.87 421.97 188.17 ;
    END
  END raddr_b_i[4]
  PIN rdata_a_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 134.83 421.97 135.13 ;
    END
  END rdata_a_o[0]
  PIN rdata_a_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 155.23 421.97 155.53 ;
    END
  END rdata_a_o[10]
  PIN rdata_a_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 151.15 421.97 151.45 ;
    END
  END rdata_a_o[11]
  PIN rdata_a_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 147.07 421.97 147.37 ;
    END
  END rdata_a_o[12]
  PIN rdata_a_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 208.27 421.97 208.57 ;
    END
  END rdata_a_o[13]
  PIN rdata_a_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 244.99 421.97 245.29 ;
    END
  END rdata_a_o[14]
  PIN rdata_a_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 277.63 421.97 277.93 ;
    END
  END rdata_a_o[15]
  PIN rdata_a_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 318.43 421.97 318.73 ;
    END
  END rdata_a_o[16]
  PIN rdata_a_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 322.51 421.97 322.81 ;
    END
  END rdata_a_o[17]
  PIN rdata_a_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  289.96 421.485 290.1 421.97 ;
    END
  END rdata_a_o[18]
  PIN rdata_a_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  252.7 421.485 252.84 421.97 ;
    END
  END rdata_a_o[19]
  PIN rdata_a_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 249.07 421.97 249.37 ;
    END
  END rdata_a_o[1]
  PIN rdata_a_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  203.02 421.485 203.16 421.97 ;
    END
  END rdata_a_o[20]
  PIN rdata_a_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  207.16 421.485 207.3 421.97 ;
    END
  END rdata_a_o[21]
  PIN rdata_a_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.04 421.485 174.18 421.97 ;
    END
  END rdata_a_o[22]
  PIN rdata_a_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140.92 421.485 141.06 421.97 ;
    END
  END rdata_a_o[23]
  PIN rdata_a_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 326.59 0.8 326.89 ;
    END
  END rdata_a_o[24]
  PIN rdata_a_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 322.51 0.8 322.81 ;
    END
  END rdata_a_o[25]
  PIN rdata_a_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 302.11 0.8 302.41 ;
    END
  END rdata_a_o[26]
  PIN rdata_a_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 261.31 0.8 261.61 ;
    END
  END rdata_a_o[27]
  PIN rdata_a_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 228.67 0.8 228.97 ;
    END
  END rdata_a_o[28]
  PIN rdata_a_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 200.11 0.8 200.41 ;
    END
  END rdata_a_o[29]
  PIN rdata_a_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 167.47 0.8 167.77 ;
    END
  END rdata_a_o[2]
  PIN rdata_a_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 187.87 0.8 188.17 ;
    END
  END rdata_a_o[30]
  PIN rdata_a_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  178.18 0 178.32 0.485 ;
    END
  END rdata_a_o[31]
  PIN rdata_a_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 130.75 0.8 131.05 ;
    END
  END rdata_a_o[3]
  PIN rdata_a_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 98.11 0.8 98.41 ;
    END
  END rdata_a_o[4]
  PIN rdata_a_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  116.08 0 116.22 0.485 ;
    END
  END rdata_a_o[5]
  PIN rdata_a_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  161.62 0 161.76 0.485 ;
    END
  END rdata_a_o[6]
  PIN rdata_a_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  203.02 0 203.16 0.485 ;
    END
  END rdata_a_o[7]
  PIN rdata_a_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  248.56 0 248.7 0.485 ;
    END
  END rdata_a_o[8]
  PIN rdata_a_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  289.96 0 290.1 0.485 ;
    END
  END rdata_a_o[9]
  PIN rdata_b_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 163.39 421.97 163.69 ;
    END
  END rdata_b_o[0]
  PIN rdata_b_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 138.91 421.97 139.21 ;
    END
  END rdata_b_o[10]
  PIN rdata_b_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 142.99 421.97 143.29 ;
    END
  END rdata_b_o[11]
  PIN rdata_b_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 159.31 421.97 159.61 ;
    END
  END rdata_b_o[12]
  PIN rdata_b_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 204.19 421.97 204.49 ;
    END
  END rdata_b_o[13]
  PIN rdata_b_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 236.83 421.97 237.13 ;
    END
  END rdata_b_o[14]
  PIN rdata_b_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 273.55 421.97 273.85 ;
    END
  END rdata_b_o[15]
  PIN rdata_b_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 293.95 421.97 294.25 ;
    END
  END rdata_b_o[16]
  PIN rdata_b_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  306.52 421.485 306.66 421.97 ;
    END
  END rdata_b_o[17]
  PIN rdata_b_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  281.68 421.485 281.82 421.97 ;
    END
  END rdata_b_o[18]
  PIN rdata_b_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  248.56 421.485 248.7 421.97 ;
    END
  END rdata_b_o[19]
  PIN rdata_b_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 240.91 421.97 241.21 ;
    END
  END rdata_b_o[1]
  PIN rdata_b_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  219.58 421.485 219.72 421.97 ;
    END
  END rdata_b_o[20]
  PIN rdata_b_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  211.3 421.485 211.44 421.97 ;
    END
  END rdata_b_o[21]
  PIN rdata_b_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  178.18 421.485 178.32 421.97 ;
    END
  END rdata_b_o[22]
  PIN rdata_b_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  145.06 421.485 145.2 421.97 ;
    END
  END rdata_b_o[23]
  PIN rdata_b_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  107.8 421.485 107.94 421.97 ;
    END
  END rdata_b_o[24]
  PIN rdata_b_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  111.94 421.485 112.08 421.97 ;
    END
  END rdata_b_o[25]
  PIN rdata_b_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 273.55 0.8 273.85 ;
    END
  END rdata_b_o[26]
  PIN rdata_b_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 257.23 0.8 257.53 ;
    END
  END rdata_b_o[27]
  PIN rdata_b_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 224.59 0.8 224.89 ;
    END
  END rdata_b_o[28]
  PIN rdata_b_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 196.03 0.8 196.33 ;
    END
  END rdata_b_o[29]
  PIN rdata_b_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 171.55 0.8 171.85 ;
    END
  END rdata_b_o[2]
  PIN rdata_b_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  190.6 0 190.74 0.485 ;
    END
  END rdata_b_o[30]
  PIN rdata_b_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  194.74 0 194.88 0.485 ;
    END
  END rdata_b_o[31]
  PIN rdata_b_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 134.83 0.8 135.13 ;
    END
  END rdata_b_o[3]
  PIN rdata_b_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.66 0 103.8 0.485 ;
    END
  END rdata_b_o[4]
  PIN rdata_b_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  111.94 0 112.08 0.485 ;
    END
  END rdata_b_o[5]
  PIN rdata_b_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  169.9 0 170.04 0.485 ;
    END
  END rdata_b_o[6]
  PIN rdata_b_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  198.88 0 199.02 0.485 ;
    END
  END rdata_b_o[7]
  PIN rdata_b_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  240.28 0 240.42 0.485 ;
    END
  END rdata_b_o[8]
  PIN rdata_b_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  265.12 0 265.26 0.485 ;
    END
  END rdata_b_o[9]
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 16.51 421.97 16.81 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  8.44 0 8.58 0.485 ;
    END
  END test_en_i
  PIN waddr_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 224.59 421.97 224.89 ;
    END
  END waddr_a_i[0]
  PIN waddr_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 216.43 421.97 216.73 ;
    END
  END waddr_a_i[1]
  PIN waddr_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 191.95 421.97 192.25 ;
    END
  END waddr_a_i[2]
  PIN waddr_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 183.79 421.97 184.09 ;
    END
  END waddr_a_i[3]
  PIN waddr_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 200.11 421.97 200.41 ;
    END
  END waddr_a_i[4]
  PIN wdata_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  269.26 0 269.4 0.485 ;
    END
  END wdata_a_i[0]
  PIN wdata_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  302.38 0 302.52 0.485 ;
    END
  END wdata_a_i[10]
  PIN wdata_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 106.27 421.97 106.57 ;
    END
  END wdata_a_i[11]
  PIN wdata_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 130.75 421.97 131.05 ;
    END
  END wdata_a_i[12]
  PIN wdata_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 220.51 421.97 220.81 ;
    END
  END wdata_a_i[13]
  PIN wdata_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 232.75 421.97 233.05 ;
    END
  END wdata_a_i[14]
  PIN wdata_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 298.03 421.97 298.33 ;
    END
  END wdata_a_i[15]
  PIN wdata_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 334.75 421.97 335.05 ;
    END
  END wdata_a_i[16]
  PIN wdata_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  314.8 421.485 314.94 421.97 ;
    END
  END wdata_a_i[17]
  PIN wdata_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  277.54 421.485 277.68 421.97 ;
    END
  END wdata_a_i[18]
  PIN wdata_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  244.42 421.485 244.56 421.97 ;
    END
  END wdata_a_i[19]
  PIN wdata_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 212.35 421.97 212.65 ;
    END
  END wdata_a_i[1]
  PIN wdata_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  198.88 421.485 199.02 421.97 ;
    END
  END wdata_a_i[20]
  PIN wdata_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  194.74 421.485 194.88 421.97 ;
    END
  END wdata_a_i[21]
  PIN wdata_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  161.62 421.485 161.76 421.97 ;
    END
  END wdata_a_i[22]
  PIN wdata_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  124.36 421.485 124.5 421.97 ;
    END
  END wdata_a_i[23]
  PIN wdata_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.4 421.485 66.54 421.97 ;
    END
  END wdata_a_i[24]
  PIN wdata_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 371.47 0.8 371.77 ;
    END
  END wdata_a_i[25]
  PIN wdata_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 314.35 0.8 314.65 ;
    END
  END wdata_a_i[26]
  PIN wdata_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 253.15 0.8 253.45 ;
    END
  END wdata_a_i[27]
  PIN wdata_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 220.51 0.8 220.81 ;
    END
  END wdata_a_i[28]
  PIN wdata_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 216.43 0.8 216.73 ;
    END
  END wdata_a_i[29]
  PIN wdata_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 163.39 0.8 163.69 ;
    END
  END wdata_a_i[2]
  PIN wdata_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 236.83 0.8 237.13 ;
    END
  END wdata_a_i[30]
  PIN wdata_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 204.19 0.8 204.49 ;
    END
  END wdata_a_i[31]
  PIN wdata_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 122.59 0.8 122.89 ;
    END
  END wdata_a_i[3]
  PIN wdata_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 77.71 0.8 78.01 ;
    END
  END wdata_a_i[4]
  PIN wdata_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.52 0 99.66 0.485 ;
    END
  END wdata_a_i[5]
  PIN wdata_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  136.78 0 136.92 0.485 ;
    END
  END wdata_a_i[6]
  PIN wdata_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.04 0 174.18 0.485 ;
    END
  END wdata_a_i[7]
  PIN wdata_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  227.86 0 228 0.485 ;
    END
  END wdata_a_i[8]
  PIN wdata_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  273.4 0 273.54 0.485 ;
    END
  END wdata_a_i[9]
  PIN we_a_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  421.17 196.03 421.97 196.33 ;
    END
  END we_a_i
  OBS
    LAYER nwell ;
     RECT  0 0 421.97 421.97 ;
    LAYER pwell ;
     RECT  0 0 421.97 421.97 ;
    LAYER li1 ;
     RECT  0 0 421.97 421.97 ;
    LAYER met1 ;
     RECT  0 0 421.97 421.97 ;
    LAYER met2 ;
     RECT  0 0 421.97 421.97 ;
    LAYER met3 ;
     RECT  0 0 421.97 421.97 ;
    LAYER met4 ;
     RECT  0 0 421.97 421.97 ;
    LAYER met5 ;
     RECT  0 0 421.97 421.97 ;
  END
END ibex_register_file_ff
END LIBRARY
