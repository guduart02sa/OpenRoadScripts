module riscv_top (clk,
    memwrite,
    ready,
    reset,
    suspend,
    valid,
    valid_reg,
    dataadr,
    instr,
    pc,
    writedata);
 input clk;
 output memwrite;
 output ready;
 input reset;
 output suspend;
 input valid;
 input valid_reg;
 output [31:0] dataadr;
 input [31:0] instr;
 output [31:0] pc;
 output [31:0] writedata;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire clk_regs;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire \dmem.ce_mem[0] ;
 wire \dmem.ce_mem[1] ;
 wire \dmem.ce_mem[2] ;
 wire \dmem.ce_mem[3] ;
 wire \dmem.inter_dmem0[0] ;
 wire \dmem.inter_dmem0[10] ;
 wire \dmem.inter_dmem0[11] ;
 wire \dmem.inter_dmem0[12] ;
 wire \dmem.inter_dmem0[13] ;
 wire \dmem.inter_dmem0[14] ;
 wire \dmem.inter_dmem0[15] ;
 wire \dmem.inter_dmem0[16] ;
 wire \dmem.inter_dmem0[17] ;
 wire \dmem.inter_dmem0[18] ;
 wire \dmem.inter_dmem0[19] ;
 wire \dmem.inter_dmem0[1] ;
 wire \dmem.inter_dmem0[20] ;
 wire \dmem.inter_dmem0[21] ;
 wire \dmem.inter_dmem0[22] ;
 wire \dmem.inter_dmem0[23] ;
 wire \dmem.inter_dmem0[24] ;
 wire \dmem.inter_dmem0[25] ;
 wire \dmem.inter_dmem0[26] ;
 wire \dmem.inter_dmem0[27] ;
 wire \dmem.inter_dmem0[28] ;
 wire \dmem.inter_dmem0[29] ;
 wire \dmem.inter_dmem0[2] ;
 wire \dmem.inter_dmem0[30] ;
 wire \dmem.inter_dmem0[31] ;
 wire \dmem.inter_dmem0[3] ;
 wire \dmem.inter_dmem0[4] ;
 wire \dmem.inter_dmem0[5] ;
 wire \dmem.inter_dmem0[6] ;
 wire \dmem.inter_dmem0[7] ;
 wire \dmem.inter_dmem0[8] ;
 wire \dmem.inter_dmem0[9] ;
 wire \dmem.inter_dmem1[0] ;
 wire \dmem.inter_dmem1[10] ;
 wire \dmem.inter_dmem1[11] ;
 wire \dmem.inter_dmem1[12] ;
 wire \dmem.inter_dmem1[13] ;
 wire \dmem.inter_dmem1[14] ;
 wire \dmem.inter_dmem1[15] ;
 wire \dmem.inter_dmem1[16] ;
 wire \dmem.inter_dmem1[17] ;
 wire \dmem.inter_dmem1[18] ;
 wire \dmem.inter_dmem1[19] ;
 wire \dmem.inter_dmem1[1] ;
 wire \dmem.inter_dmem1[20] ;
 wire \dmem.inter_dmem1[21] ;
 wire \dmem.inter_dmem1[22] ;
 wire \dmem.inter_dmem1[23] ;
 wire \dmem.inter_dmem1[24] ;
 wire \dmem.inter_dmem1[25] ;
 wire \dmem.inter_dmem1[26] ;
 wire \dmem.inter_dmem1[27] ;
 wire \dmem.inter_dmem1[28] ;
 wire \dmem.inter_dmem1[29] ;
 wire \dmem.inter_dmem1[2] ;
 wire \dmem.inter_dmem1[30] ;
 wire \dmem.inter_dmem1[31] ;
 wire \dmem.inter_dmem1[3] ;
 wire \dmem.inter_dmem1[4] ;
 wire \dmem.inter_dmem1[5] ;
 wire \dmem.inter_dmem1[6] ;
 wire \dmem.inter_dmem1[7] ;
 wire \dmem.inter_dmem1[8] ;
 wire \dmem.inter_dmem1[9] ;
 wire \dmem.inter_dmem2[0] ;
 wire \dmem.inter_dmem2[10] ;
 wire \dmem.inter_dmem2[11] ;
 wire \dmem.inter_dmem2[12] ;
 wire \dmem.inter_dmem2[13] ;
 wire \dmem.inter_dmem2[14] ;
 wire \dmem.inter_dmem2[15] ;
 wire \dmem.inter_dmem2[16] ;
 wire \dmem.inter_dmem2[17] ;
 wire \dmem.inter_dmem2[18] ;
 wire \dmem.inter_dmem2[19] ;
 wire \dmem.inter_dmem2[1] ;
 wire \dmem.inter_dmem2[20] ;
 wire \dmem.inter_dmem2[21] ;
 wire \dmem.inter_dmem2[22] ;
 wire \dmem.inter_dmem2[23] ;
 wire \dmem.inter_dmem2[24] ;
 wire \dmem.inter_dmem2[25] ;
 wire \dmem.inter_dmem2[26] ;
 wire \dmem.inter_dmem2[27] ;
 wire \dmem.inter_dmem2[28] ;
 wire \dmem.inter_dmem2[29] ;
 wire \dmem.inter_dmem2[2] ;
 wire \dmem.inter_dmem2[30] ;
 wire \dmem.inter_dmem2[31] ;
 wire \dmem.inter_dmem2[3] ;
 wire \dmem.inter_dmem2[4] ;
 wire \dmem.inter_dmem2[5] ;
 wire \dmem.inter_dmem2[6] ;
 wire \dmem.inter_dmem2[7] ;
 wire \dmem.inter_dmem2[8] ;
 wire \dmem.inter_dmem2[9] ;
 wire \dmem.inter_dmem3[0] ;
 wire \dmem.inter_dmem3[10] ;
 wire \dmem.inter_dmem3[11] ;
 wire \dmem.inter_dmem3[12] ;
 wire \dmem.inter_dmem3[13] ;
 wire \dmem.inter_dmem3[14] ;
 wire \dmem.inter_dmem3[15] ;
 wire \dmem.inter_dmem3[16] ;
 wire \dmem.inter_dmem3[17] ;
 wire \dmem.inter_dmem3[18] ;
 wire \dmem.inter_dmem3[19] ;
 wire \dmem.inter_dmem3[1] ;
 wire \dmem.inter_dmem3[20] ;
 wire \dmem.inter_dmem3[21] ;
 wire \dmem.inter_dmem3[22] ;
 wire \dmem.inter_dmem3[23] ;
 wire \dmem.inter_dmem3[24] ;
 wire \dmem.inter_dmem3[25] ;
 wire \dmem.inter_dmem3[26] ;
 wire \dmem.inter_dmem3[27] ;
 wire \dmem.inter_dmem3[28] ;
 wire \dmem.inter_dmem3[29] ;
 wire \dmem.inter_dmem3[2] ;
 wire \dmem.inter_dmem3[30] ;
 wire \dmem.inter_dmem3[31] ;
 wire \dmem.inter_dmem3[3] ;
 wire \dmem.inter_dmem3[4] ;
 wire \dmem.inter_dmem3[5] ;
 wire \dmem.inter_dmem3[6] ;
 wire \dmem.inter_dmem3[7] ;
 wire \dmem.inter_dmem3[8] ;
 wire \dmem.inter_dmem3[9] ;
 wire \dmem.we_mem[0] ;
 wire \dmem.we_mem[1] ;
 wire \dmem.we_mem[2] ;
 wire \dmem.we_mem[3] ;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire \riscv.dp.ISRmux.d0[10] ;
 wire \riscv.dp.ISRmux.d0[11] ;
 wire \riscv.dp.ISRmux.d0[12] ;
 wire \riscv.dp.ISRmux.d0[13] ;
 wire \riscv.dp.ISRmux.d0[14] ;
 wire \riscv.dp.ISRmux.d0[15] ;
 wire \riscv.dp.ISRmux.d0[16] ;
 wire \riscv.dp.ISRmux.d0[17] ;
 wire \riscv.dp.ISRmux.d0[18] ;
 wire \riscv.dp.ISRmux.d0[19] ;
 wire \riscv.dp.ISRmux.d0[20] ;
 wire \riscv.dp.ISRmux.d0[21] ;
 wire \riscv.dp.ISRmux.d0[22] ;
 wire \riscv.dp.ISRmux.d0[23] ;
 wire \riscv.dp.ISRmux.d0[24] ;
 wire \riscv.dp.ISRmux.d0[25] ;
 wire \riscv.dp.ISRmux.d0[26] ;
 wire \riscv.dp.ISRmux.d0[27] ;
 wire \riscv.dp.ISRmux.d0[28] ;
 wire \riscv.dp.ISRmux.d0[29] ;
 wire \riscv.dp.ISRmux.d0[2] ;
 wire \riscv.dp.ISRmux.d0[30] ;
 wire \riscv.dp.ISRmux.d0[31] ;
 wire \riscv.dp.ISRmux.d0[3] ;
 wire \riscv.dp.ISRmux.d0[4] ;
 wire \riscv.dp.ISRmux.d0[5] ;
 wire \riscv.dp.ISRmux.d0[6] ;
 wire \riscv.dp.ISRmux.d0[7] ;
 wire \riscv.dp.ISRmux.d0[8] ;
 wire \riscv.dp.ISRmux.d0[9] ;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_2_0_0_clk_regs;
 wire clknet_2_1_0_clk_regs;
 wire clknet_2_2_0_clk_regs;
 wire clknet_2_3_0_clk_regs;

 INVx3_ASAP7_75t_R _10170_ (.A(_01159_),
    .Y(_03372_));
 BUFx12f_ASAP7_75t_R _10171_ (.A(_03372_),
    .Y(_03373_));
 BUFx12f_ASAP7_75t_R _10172_ (.A(_03373_),
    .Y(_03374_));
 BUFx16f_ASAP7_75t_R _10173_ (.A(_03374_),
    .Y(_03375_));
 BUFx16f_ASAP7_75t_R _10174_ (.A(_03375_),
    .Y(_03376_));
 BUFx12f_ASAP7_75t_R _10175_ (.A(_03376_),
    .Y(_03377_));
 BUFx10_ASAP7_75t_R _10176_ (.A(_03377_),
    .Y(_03378_));
 BUFx10_ASAP7_75t_R _10177_ (.A(_03378_),
    .Y(_03379_));
 BUFx6f_ASAP7_75t_R _10178_ (.A(_03379_),
    .Y(_03380_));
 BUFx6f_ASAP7_75t_R _10179_ (.A(_03380_),
    .Y(_03381_));
 BUFx12_ASAP7_75t_R _10180_ (.A(_03381_),
    .Y(_03382_));
 BUFx6f_ASAP7_75t_R _10181_ (.A(_03382_),
    .Y(net89));
 NAND2x1_ASAP7_75t_R _10182_ (.A(net15),
    .B(_03373_),
    .Y(_03383_));
 BUFx4f_ASAP7_75t_R _10183_ (.A(_03383_),
    .Y(_03384_));
 INVx3_ASAP7_75t_R _10184_ (.A(net13),
    .Y(_03385_));
 BUFx6f_ASAP7_75t_R _10185_ (.A(_03385_),
    .Y(_03386_));
 BUFx4f_ASAP7_75t_R _10186_ (.A(net13),
    .Y(_03387_));
 BUFx4f_ASAP7_75t_R _10187_ (.A(_03387_),
    .Y(_03388_));
 AND2x2_ASAP7_75t_R _10188_ (.A(_03388_),
    .B(_00027_),
    .Y(_03389_));
 AO21x1_ASAP7_75t_R _10189_ (.A1(_03386_),
    .A2(_00025_),
    .B(_03389_),
    .Y(_03390_));
 BUFx6f_ASAP7_75t_R _10190_ (.A(net13),
    .Y(_03391_));
 BUFx4f_ASAP7_75t_R _10191_ (.A(_03391_),
    .Y(_03392_));
 BUFx12_ASAP7_75t_R _10192_ (.A(_03372_),
    .Y(_03393_));
 BUFx16f_ASAP7_75t_R _10193_ (.A(_03393_),
    .Y(_03394_));
 BUFx12_ASAP7_75t_R _10194_ (.A(_03394_),
    .Y(_03395_));
 BUFx4f_ASAP7_75t_R _10195_ (.A(net15),
    .Y(_03396_));
 AO21x1_ASAP7_75t_R _10196_ (.A1(_03385_),
    .A2(_00009_),
    .B(_03396_),
    .Y(_03397_));
 AO22x1_ASAP7_75t_R _10197_ (.A1(_03392_),
    .A2(_00011_),
    .B1(_03395_),
    .B2(_03397_),
    .Y(_03398_));
 BUFx6f_ASAP7_75t_R _10198_ (.A(net12),
    .Y(_03399_));
 BUFx6f_ASAP7_75t_R _10199_ (.A(_03399_),
    .Y(_03400_));
 OA211x2_ASAP7_75t_R _10200_ (.A1(_03384_),
    .A2(_03390_),
    .B(_03398_),
    .C(_03400_),
    .Y(_03401_));
 BUFx12f_ASAP7_75t_R _10201_ (.A(_03373_),
    .Y(_03402_));
 AND3x1_ASAP7_75t_R _10202_ (.A(_03396_),
    .B(_00024_),
    .C(_03402_),
    .Y(_03403_));
 AO21x1_ASAP7_75t_R _10203_ (.A1(_00008_),
    .A2(_03384_),
    .B(_03403_),
    .Y(_03404_));
 NOR2x2_ASAP7_75t_R _10204_ (.A(_03399_),
    .B(_03391_),
    .Y(_03405_));
 INVx1_ASAP7_75t_R _10205_ (.A(net12),
    .Y(_03406_));
 BUFx4f_ASAP7_75t_R _10206_ (.A(_03406_),
    .Y(_03407_));
 AND2x2_ASAP7_75t_R _10207_ (.A(_03407_),
    .B(_03392_),
    .Y(_03408_));
 AND3x1_ASAP7_75t_R _10208_ (.A(_03396_),
    .B(_00026_),
    .C(_03402_),
    .Y(_03409_));
 AO21x1_ASAP7_75t_R _10209_ (.A1(_00010_),
    .A2(_03384_),
    .B(_03409_),
    .Y(_03410_));
 BUFx6f_ASAP7_75t_R _10210_ (.A(instr[22]),
    .Y(_03411_));
 BUFx6f_ASAP7_75t_R _10211_ (.A(_03411_),
    .Y(_03412_));
 CKINVDCx10_ASAP7_75t_R _10212_ (.A(net14),
    .Y(_03413_));
 BUFx10_ASAP7_75t_R _10213_ (.A(_01159_),
    .Y(_03414_));
 BUFx12_ASAP7_75t_R _10214_ (.A(_03414_),
    .Y(_03415_));
 OR3x1_ASAP7_75t_R _10215_ (.A(_03412_),
    .B(_03413_),
    .C(_03415_),
    .Y(_03416_));
 AO221x1_ASAP7_75t_R _10216_ (.A1(_03404_),
    .A2(_03405_),
    .B1(_03408_),
    .B2(_03410_),
    .C(_03416_),
    .Y(_03417_));
 INVx5_ASAP7_75t_R _10217_ (.A(_03411_),
    .Y(_03418_));
 BUFx10_ASAP7_75t_R _10218_ (.A(_03415_),
    .Y(_03419_));
 OR3x4_ASAP7_75t_R _10219_ (.A(_03418_),
    .B(_03413_),
    .C(_03419_),
    .Y(_03420_));
 BUFx4f_ASAP7_75t_R _10220_ (.A(_03406_),
    .Y(_03421_));
 BUFx4f_ASAP7_75t_R _10221_ (.A(_03421_),
    .Y(_03422_));
 BUFx4f_ASAP7_75t_R _10222_ (.A(_03422_),
    .Y(_03423_));
 BUFx4f_ASAP7_75t_R _10223_ (.A(_03385_),
    .Y(_03424_));
 AND3x1_ASAP7_75t_R _10224_ (.A(_03424_),
    .B(_00013_),
    .C(_03395_),
    .Y(_03425_));
 BUFx4f_ASAP7_75t_R _10225_ (.A(_03388_),
    .Y(_03426_));
 AO21x1_ASAP7_75t_R _10226_ (.A1(_03426_),
    .A2(_00015_),
    .B(_03396_),
    .Y(_03427_));
 AND3x1_ASAP7_75t_R _10227_ (.A(_03424_),
    .B(_00029_),
    .C(_03395_),
    .Y(_03428_));
 INVx2_ASAP7_75t_R _10228_ (.A(net15),
    .Y(_03429_));
 AO21x1_ASAP7_75t_R _10229_ (.A1(_03426_),
    .A2(_00031_),
    .B(_03429_),
    .Y(_03430_));
 OAI22x1_ASAP7_75t_R _10230_ (.A1(_03425_),
    .A2(_03427_),
    .B1(_03428_),
    .B2(_03430_),
    .Y(_03431_));
 BUFx4f_ASAP7_75t_R _10231_ (.A(_03387_),
    .Y(_03432_));
 INVx1_ASAP7_75t_R _10232_ (.A(_00012_),
    .Y(_03433_));
 NAND2x1_ASAP7_75t_R _10233_ (.A(_03391_),
    .B(_00014_),
    .Y(_03434_));
 OA211x2_ASAP7_75t_R _10234_ (.A1(_03432_),
    .A2(_03433_),
    .B(_03429_),
    .C(_03434_),
    .Y(_03435_));
 INVx2_ASAP7_75t_R _10235_ (.A(_00028_),
    .Y(_03436_));
 NAND2x1_ASAP7_75t_R _10236_ (.A(_03391_),
    .B(_00030_),
    .Y(_03437_));
 OA211x2_ASAP7_75t_R _10237_ (.A1(_03432_),
    .A2(_03436_),
    .B(_03437_),
    .C(_03396_),
    .Y(_03438_));
 OR3x1_ASAP7_75t_R _10238_ (.A(_03400_),
    .B(_03435_),
    .C(_03438_),
    .Y(_03439_));
 OAI21x1_ASAP7_75t_R _10239_ (.A1(_03423_),
    .A2(_03431_),
    .B(_03439_),
    .Y(_03440_));
 OA22x2_ASAP7_75t_R _10240_ (.A1(_03401_),
    .A2(_03417_),
    .B1(_03420_),
    .B2(_03440_),
    .Y(_03441_));
 BUFx6f_ASAP7_75t_R _10241_ (.A(net14),
    .Y(_03442_));
 BUFx12f_ASAP7_75t_R _10242_ (.A(_03394_),
    .Y(_03443_));
 NAND2x2_ASAP7_75t_R _10243_ (.A(_03442_),
    .B(_03443_),
    .Y(_03444_));
 OR5x2_ASAP7_75t_R _10244_ (.A(net12),
    .B(_03387_),
    .C(_03411_),
    .D(net14),
    .E(net15),
    .Y(_03445_));
 AND2x2_ASAP7_75t_R _10245_ (.A(_03374_),
    .B(_03445_),
    .Y(_03446_));
 BUFx16f_ASAP7_75t_R _10246_ (.A(_03446_),
    .Y(_03447_));
 NAND2x2_ASAP7_75t_R _10247_ (.A(_03444_),
    .B(_03447_),
    .Y(_03448_));
 NAND2x2_ASAP7_75t_R _10248_ (.A(_03411_),
    .B(_03394_),
    .Y(_03449_));
 AND3x1_ASAP7_75t_R _10249_ (.A(_03399_),
    .B(_00005_),
    .C(_03394_),
    .Y(_03450_));
 AO21x1_ASAP7_75t_R _10250_ (.A1(_03421_),
    .A2(_00004_),
    .B(_03391_),
    .Y(_03451_));
 AND2x2_ASAP7_75t_R _10251_ (.A(net12),
    .B(_00007_),
    .Y(_03452_));
 AO21x1_ASAP7_75t_R _10252_ (.A1(_03421_),
    .A2(_00006_),
    .B(_03452_),
    .Y(_03453_));
 OA22x2_ASAP7_75t_R _10253_ (.A1(_03450_),
    .A2(_03451_),
    .B1(_03453_),
    .B2(_03424_),
    .Y(_03454_));
 AND2x2_ASAP7_75t_R _10254_ (.A(_03387_),
    .B(_00003_),
    .Y(_03455_));
 AO21x1_ASAP7_75t_R _10255_ (.A1(_00001_),
    .A2(_03385_),
    .B(_03455_),
    .Y(_03456_));
 NAND2x1_ASAP7_75t_R _10256_ (.A(_03399_),
    .B(_03418_),
    .Y(_03457_));
 AND2x2_ASAP7_75t_R _10257_ (.A(net13),
    .B(_00002_),
    .Y(_03458_));
 OR3x1_ASAP7_75t_R _10258_ (.A(net12),
    .B(_03411_),
    .C(_03458_),
    .Y(_03459_));
 OA211x2_ASAP7_75t_R _10259_ (.A1(_03456_),
    .A2(_03457_),
    .B(_03459_),
    .C(_03374_),
    .Y(_03460_));
 OA21x2_ASAP7_75t_R _10260_ (.A1(_03415_),
    .A2(_03405_),
    .B(_00000_),
    .Y(_03461_));
 OA222x2_ASAP7_75t_R _10261_ (.A1(_03429_),
    .A2(_03419_),
    .B1(_03449_),
    .B2(_03454_),
    .C1(_03460_),
    .C2(_03461_),
    .Y(_03462_));
 AND3x1_ASAP7_75t_R _10262_ (.A(_03424_),
    .B(_00017_),
    .C(_03374_),
    .Y(_03463_));
 AO21x1_ASAP7_75t_R _10263_ (.A1(_03432_),
    .A2(_00019_),
    .B(_03407_),
    .Y(_03464_));
 AND2x2_ASAP7_75t_R _10264_ (.A(_03391_),
    .B(_00018_),
    .Y(_03465_));
 AO21x1_ASAP7_75t_R _10265_ (.A1(_03424_),
    .A2(_00016_),
    .B(_03465_),
    .Y(_03466_));
 OAI22x1_ASAP7_75t_R _10266_ (.A1(_03463_),
    .A2(_03464_),
    .B1(_03466_),
    .B2(_03400_),
    .Y(_03467_));
 INVx2_ASAP7_75t_R _10267_ (.A(_00020_),
    .Y(_03468_));
 NAND2x1_ASAP7_75t_R _10268_ (.A(_03387_),
    .B(_00022_),
    .Y(_03469_));
 OA211x2_ASAP7_75t_R _10269_ (.A1(_03388_),
    .A2(_03468_),
    .B(_03469_),
    .C(_03421_),
    .Y(_03470_));
 INVx2_ASAP7_75t_R _10270_ (.A(_00021_),
    .Y(_03471_));
 NAND2x1_ASAP7_75t_R _10271_ (.A(_03387_),
    .B(_00023_),
    .Y(_03472_));
 OA211x2_ASAP7_75t_R _10272_ (.A1(_03388_),
    .A2(_03471_),
    .B(_03472_),
    .C(_03399_),
    .Y(_03473_));
 AND2x6_ASAP7_75t_R _10273_ (.A(_03411_),
    .B(_03394_),
    .Y(_03474_));
 OA21x2_ASAP7_75t_R _10274_ (.A1(_03470_),
    .A2(_03473_),
    .B(_03474_),
    .Y(_03475_));
 AOI211x1_ASAP7_75t_R _10275_ (.A1(_03418_),
    .A2(_03467_),
    .B(_03475_),
    .C(_03384_),
    .Y(_03476_));
 OR3x4_ASAP7_75t_R _10276_ (.A(_03448_),
    .B(_03462_),
    .C(_03476_),
    .Y(_03477_));
 AND2x6_ASAP7_75t_R _10277_ (.A(_03441_),
    .B(_03477_),
    .Y(_03478_));
 CKINVDCx9p33_ASAP7_75t_R _10278_ (.A(_03478_),
    .Y(net99));
 INVx4_ASAP7_75t_R _10279_ (.A(_01116_),
    .Y(net73));
 INVx4_ASAP7_75t_R _10280_ (.A(_01113_),
    .Y(net72));
 INVx3_ASAP7_75t_R _10281_ (.A(_01122_),
    .Y(net75));
 INVx4_ASAP7_75t_R _10282_ (.A(_01119_),
    .Y(net74));
 INVx4_ASAP7_75t_R _10283_ (.A(_01128_),
    .Y(net78));
 INVx4_ASAP7_75t_R _10284_ (.A(_01125_),
    .Y(net77));
 INVx4_ASAP7_75t_R _10285_ (.A(_01134_),
    .Y(net80));
 INVx3_ASAP7_75t_R _10286_ (.A(_01131_),
    .Y(net79));
 INVx4_ASAP7_75t_R _10287_ (.A(_01140_),
    .Y(net82));
 INVx4_ASAP7_75t_R _10288_ (.A(_01137_),
    .Y(net81));
 INVx3_ASAP7_75t_R _10289_ (.A(_01146_),
    .Y(net84));
 INVx4_ASAP7_75t_R _10290_ (.A(_01143_),
    .Y(net83));
 INVx4_ASAP7_75t_R _10291_ (.A(_01152_),
    .Y(net86));
 INVx4_ASAP7_75t_R _10292_ (.A(_01149_),
    .Y(net85));
 INVx4_ASAP7_75t_R _10293_ (.A(_01155_),
    .Y(net88));
 INVx3_ASAP7_75t_R _10294_ (.A(_01092_),
    .Y(net96));
 CKINVDCx5p33_ASAP7_75t_R _10295_ (.A(_01089_),
    .Y(net95));
 INVx5_ASAP7_75t_R _10296_ (.A(_01098_),
    .Y(net67));
 INVx5_ASAP7_75t_R _10297_ (.A(_01095_),
    .Y(net66));
 INVx3_ASAP7_75t_R _10298_ (.A(_01104_),
    .Y(net69));
 INVx4_ASAP7_75t_R _10299_ (.A(_01101_),
    .Y(net68));
 INVx4_ASAP7_75t_R _10300_ (.A(_01110_),
    .Y(net71));
 INVx4_ASAP7_75t_R _10301_ (.A(_01107_),
    .Y(net70));
 INVx4_ASAP7_75t_R _10302_ (.A(_01080_),
    .Y(net92));
 INVx3_ASAP7_75t_R _10303_ (.A(_01077_),
    .Y(net91));
 INVx4_ASAP7_75t_R _10304_ (.A(_01086_),
    .Y(net94));
 BUFx6f_ASAP7_75t_R _10305_ (.A(_01083_),
    .Y(_03479_));
 INVx3_ASAP7_75t_R _10306_ (.A(_03479_),
    .Y(net93));
 INVx4_ASAP7_75t_R _10307_ (.A(_01070_),
    .Y(net76));
 INVx4_ASAP7_75t_R _10308_ (.A(_01068_),
    .Y(net65));
 BUFx12f_ASAP7_75t_R _10309_ (.A(_03415_),
    .Y(_03480_));
 BUFx12f_ASAP7_75t_R _10310_ (.A(_03480_),
    .Y(_03481_));
 BUFx12f_ASAP7_75t_R _10311_ (.A(_03481_),
    .Y(_03482_));
 BUFx4f_ASAP7_75t_R _10312_ (.A(net6),
    .Y(_03483_));
 AND4x2_ASAP7_75t_R _10313_ (.A(_01134_),
    .B(_01137_),
    .C(_01140_),
    .D(_01155_),
    .Y(_03484_));
 AND4x2_ASAP7_75t_R _10314_ (.A(_01143_),
    .B(_01146_),
    .C(_01149_),
    .D(_01152_),
    .Y(_03485_));
 AND2x6_ASAP7_75t_R _10315_ (.A(_03484_),
    .B(_03485_),
    .Y(_03486_));
 AND4x2_ASAP7_75t_R _10316_ (.A(_01159_),
    .B(_01113_),
    .C(_01116_),
    .D(_01131_),
    .Y(_03487_));
 AND4x2_ASAP7_75t_R _10317_ (.A(_01119_),
    .B(_01122_),
    .C(_01125_),
    .D(_01128_),
    .Y(_03488_));
 AND2x6_ASAP7_75t_R _10318_ (.A(_03487_),
    .B(_03488_),
    .Y(_03489_));
 INVx5_ASAP7_75t_R _10319_ (.A(_00033_),
    .Y(_03490_));
 AND4x2_ASAP7_75t_R _10320_ (.A(_01086_),
    .B(_01092_),
    .C(_01095_),
    .D(_01110_),
    .Y(_03491_));
 AND4x2_ASAP7_75t_R _10321_ (.A(_01098_),
    .B(_01101_),
    .C(_01104_),
    .D(_01107_),
    .Y(_03492_));
 AND4x2_ASAP7_75t_R _10322_ (.A(_01070_),
    .B(_01077_),
    .C(_01080_),
    .D(_03479_),
    .Y(_03493_));
 AND2x4_ASAP7_75t_R _10323_ (.A(_01068_),
    .B(_01089_),
    .Y(_03494_));
 AND5x2_ASAP7_75t_R _10324_ (.A(_03490_),
    .B(_03491_),
    .C(_03492_),
    .D(_03493_),
    .E(_03494_),
    .Y(_03495_));
 AO32x1_ASAP7_75t_R _10325_ (.A1(_03486_),
    .A2(_03489_),
    .A3(_03495_),
    .B1(net27),
    .B2(_03393_),
    .Y(_03496_));
 BUFx3_ASAP7_75t_R _10326_ (.A(_03496_),
    .Y(_03497_));
 AND2x2_ASAP7_75t_R _10327_ (.A(net11),
    .B(net26),
    .Y(_03498_));
 NOR2x1_ASAP7_75t_R _10328_ (.A(net21),
    .B(net24),
    .Y(_03499_));
 AND4x1_ASAP7_75t_R _10329_ (.A(net1),
    .B(_03372_),
    .C(_03498_),
    .D(_03499_),
    .Y(_03500_));
 BUFx4f_ASAP7_75t_R _10330_ (.A(_03500_),
    .Y(_03501_));
 NAND2x2_ASAP7_75t_R _10331_ (.A(_03393_),
    .B(net25),
    .Y(_03502_));
 AND2x4_ASAP7_75t_R _10332_ (.A(_03501_),
    .B(_03502_),
    .Y(_03503_));
 NAND2x2_ASAP7_75t_R _10333_ (.A(_03497_),
    .B(_03503_),
    .Y(_03504_));
 INVx1_ASAP7_75t_R _10334_ (.A(net24),
    .Y(_03505_));
 AND4x2_ASAP7_75t_R _10335_ (.A(net1),
    .B(_03372_),
    .C(net11),
    .D(_03505_),
    .Y(_03506_));
 INVx1_ASAP7_75t_R _10336_ (.A(net27),
    .Y(_03507_));
 AND4x2_ASAP7_75t_R _10337_ (.A(_03372_),
    .B(net21),
    .C(_03507_),
    .D(net25),
    .Y(_03508_));
 NAND2x2_ASAP7_75t_R _10338_ (.A(_03506_),
    .B(_03508_),
    .Y(_03509_));
 BUFx6f_ASAP7_75t_R _10339_ (.A(_00032_),
    .Y(_03510_));
 NAND2x2_ASAP7_75t_R _10340_ (.A(_03484_),
    .B(_03485_),
    .Y(_03511_));
 NAND2x2_ASAP7_75t_R _10341_ (.A(_03487_),
    .B(_03488_),
    .Y(_03512_));
 NAND2x2_ASAP7_75t_R _10342_ (.A(_03491_),
    .B(_03492_),
    .Y(_03513_));
 NAND2x2_ASAP7_75t_R _10343_ (.A(_03493_),
    .B(_03494_),
    .Y(_03514_));
 OR5x1_ASAP7_75t_R _10344_ (.A(_03510_),
    .B(_03511_),
    .C(_03512_),
    .D(_03513_),
    .E(_03514_),
    .Y(_03515_));
 BUFx6f_ASAP7_75t_R _10345_ (.A(_03515_),
    .Y(_03516_));
 AND2x2_ASAP7_75t_R _10346_ (.A(_03509_),
    .B(_03516_),
    .Y(_03517_));
 BUFx16f_ASAP7_75t_R _10347_ (.A(_03517_),
    .Y(_03518_));
 NAND2x2_ASAP7_75t_R _10348_ (.A(_03504_),
    .B(_03518_),
    .Y(_03519_));
 INVx1_ASAP7_75t_R _10349_ (.A(net1),
    .Y(_03520_));
 INVx1_ASAP7_75t_R _10350_ (.A(net11),
    .Y(_03521_));
 OR4x2_ASAP7_75t_R _10351_ (.A(_03520_),
    .B(_01159_),
    .C(_03521_),
    .D(net24),
    .Y(_03522_));
 BUFx6f_ASAP7_75t_R _10352_ (.A(_03522_),
    .Y(_03523_));
 BUFx12_ASAP7_75t_R _10353_ (.A(_03523_),
    .Y(_03524_));
 OR3x2_ASAP7_75t_R _10354_ (.A(net21),
    .B(net27),
    .C(net25),
    .Y(_03525_));
 NOR2x2_ASAP7_75t_R _10355_ (.A(_03524_),
    .B(_03525_),
    .Y(_03526_));
 OR4x2_ASAP7_75t_R _10356_ (.A(_03482_),
    .B(_03483_),
    .C(_03519_),
    .D(_03526_),
    .Y(_03527_));
 BUFx4f_ASAP7_75t_R _10357_ (.A(net5),
    .Y(_03528_));
 INVx1_ASAP7_75t_R _10358_ (.A(net25),
    .Y(_03529_));
 OR3x2_ASAP7_75t_R _10359_ (.A(_03414_),
    .B(net27),
    .C(_03529_),
    .Y(_03530_));
 NAND2x1_ASAP7_75t_R _10360_ (.A(net22),
    .B(_03501_),
    .Y(_03531_));
 AO21x2_ASAP7_75t_R _10361_ (.A1(_03530_),
    .A2(_03516_),
    .B(_03531_),
    .Y(_03532_));
 NAND2x1_ASAP7_75t_R _10362_ (.A(_03528_),
    .B(_03532_),
    .Y(_03533_));
 BUFx4f_ASAP7_75t_R _10363_ (.A(net4),
    .Y(_03534_));
 OR3x1_ASAP7_75t_R _10364_ (.A(_03528_),
    .B(_03534_),
    .C(_03532_),
    .Y(_03535_));
 AND2x2_ASAP7_75t_R _10365_ (.A(_03533_),
    .B(_03535_),
    .Y(_03536_));
 NOR2x2_ASAP7_75t_R _10366_ (.A(_03527_),
    .B(_03536_),
    .Y(_03537_));
 BUFx12f_ASAP7_75t_R _10367_ (.A(_03537_),
    .Y(_03538_));
 NAND2x2_ASAP7_75t_R _10368_ (.A(_03509_),
    .B(_03516_),
    .Y(_03539_));
 AND5x2_ASAP7_75t_R _10369_ (.A(net1),
    .B(_03393_),
    .C(net21),
    .D(net24),
    .E(_03498_),
    .Y(_03540_));
 OR2x2_ASAP7_75t_R _10370_ (.A(_03501_),
    .B(_03540_),
    .Y(_03541_));
 AND4x2_ASAP7_75t_R _10371_ (.A(_03497_),
    .B(_03502_),
    .C(_03516_),
    .D(_03541_),
    .Y(_03542_));
 NAND2x1_ASAP7_75t_R _10372_ (.A(net11),
    .B(net26),
    .Y(_03543_));
 OR2x2_ASAP7_75t_R _10373_ (.A(net21),
    .B(net24),
    .Y(_03544_));
 OR2x2_ASAP7_75t_R _10374_ (.A(net27),
    .B(net25),
    .Y(_03545_));
 OR5x1_ASAP7_75t_R _10375_ (.A(_03520_),
    .B(_01159_),
    .C(_03543_),
    .D(_03544_),
    .E(_03545_),
    .Y(_03546_));
 BUFx4f_ASAP7_75t_R _10376_ (.A(_03546_),
    .Y(_03547_));
 NAND2x2_ASAP7_75t_R _10377_ (.A(_03399_),
    .B(_03402_),
    .Y(_03548_));
 BUFx12f_ASAP7_75t_R _10378_ (.A(_03402_),
    .Y(_03549_));
 AOI21x1_ASAP7_75t_R _10379_ (.A1(_03549_),
    .A2(net28),
    .B(_03547_),
    .Y(_03550_));
 AO21x1_ASAP7_75t_R _10380_ (.A1(_03547_),
    .A2(_03548_),
    .B(_03550_),
    .Y(_03551_));
 OR3x4_ASAP7_75t_R _10381_ (.A(_03539_),
    .B(_03542_),
    .C(_03551_),
    .Y(_03552_));
 INVx4_ASAP7_75t_R _10382_ (.A(_03552_),
    .Y(_10106_));
 NAND2x2_ASAP7_75t_R _10383_ (.A(_03501_),
    .B(_03502_),
    .Y(_03553_));
 INVx4_ASAP7_75t_R _10384_ (.A(_03510_),
    .Y(_03554_));
 AND5x2_ASAP7_75t_R _10385_ (.A(_03554_),
    .B(_03491_),
    .C(_03492_),
    .D(_03493_),
    .E(_03494_),
    .Y(_03555_));
 NAND3x2_ASAP7_75t_R _10386_ (.B(_03489_),
    .C(_03555_),
    .Y(_03556_),
    .A(_03486_));
 BUFx6f_ASAP7_75t_R _10387_ (.A(_03556_),
    .Y(_03557_));
 OR5x1_ASAP7_75t_R _10388_ (.A(_03520_),
    .B(_01159_),
    .C(_03521_),
    .D(net24),
    .E(_03525_),
    .Y(_03558_));
 BUFx4f_ASAP7_75t_R _10389_ (.A(_03558_),
    .Y(_03559_));
 OR2x2_ASAP7_75t_R _10390_ (.A(_01159_),
    .B(net26),
    .Y(_03560_));
 OR2x2_ASAP7_75t_R _10391_ (.A(_03559_),
    .B(_03560_),
    .Y(_03561_));
 BUFx4f_ASAP7_75t_R _10392_ (.A(_03561_),
    .Y(_03562_));
 NAND2x1_ASAP7_75t_R _10393_ (.A(_03510_),
    .B(_00033_),
    .Y(_03563_));
 INVx1_ASAP7_75t_R _10394_ (.A(_03563_),
    .Y(_03564_));
 OR5x1_ASAP7_75t_R _10395_ (.A(_03511_),
    .B(_03512_),
    .C(_03513_),
    .D(_03514_),
    .E(_03564_),
    .Y(_03565_));
 BUFx4f_ASAP7_75t_R _10396_ (.A(_03565_),
    .Y(_03566_));
 INVx1_ASAP7_75t_R _10397_ (.A(net21),
    .Y(_03567_));
 AO21x1_ASAP7_75t_R _10398_ (.A1(_03567_),
    .A2(_03560_),
    .B(_03522_),
    .Y(_03568_));
 AO32x2_ASAP7_75t_R _10399_ (.A1(_03530_),
    .A2(_03557_),
    .A3(_03562_),
    .B1(_03566_),
    .B2(_03568_),
    .Y(_03569_));
 OR5x2_ASAP7_75t_R _10400_ (.A(_00033_),
    .B(_03511_),
    .C(_03512_),
    .D(_03513_),
    .E(_03514_),
    .Y(_03570_));
 OR5x2_ASAP7_75t_R _10401_ (.A(_03520_),
    .B(_03414_),
    .C(_03567_),
    .D(_03507_),
    .E(_03543_),
    .Y(_03571_));
 AND3x4_ASAP7_75t_R _10402_ (.A(_03486_),
    .B(_03489_),
    .C(_03555_),
    .Y(_03572_));
 AO221x1_ASAP7_75t_R _10403_ (.A1(_03394_),
    .A2(net25),
    .B1(_03570_),
    .B2(_03571_),
    .C(_03572_),
    .Y(_03573_));
 BUFx4f_ASAP7_75t_R _10404_ (.A(_03573_),
    .Y(_03574_));
 NAND3x2_ASAP7_75t_R _10405_ (.B(_03569_),
    .C(_03574_),
    .Y(_03575_),
    .A(_03553_));
 NAND2x2_ASAP7_75t_R _10406_ (.A(_10106_),
    .B(_03575_),
    .Y(_03576_));
 AO21x2_ASAP7_75t_R _10407_ (.A1(_03441_),
    .A2(_03477_),
    .B(_03575_),
    .Y(_03577_));
 AND2x2_ASAP7_75t_R _10408_ (.A(_03576_),
    .B(_03577_),
    .Y(_03578_));
 BUFx4f_ASAP7_75t_R _10409_ (.A(_03578_),
    .Y(_03579_));
 BUFx4f_ASAP7_75t_R _10410_ (.A(_03579_),
    .Y(_03580_));
 BUFx6f_ASAP7_75t_R _10411_ (.A(_03580_),
    .Y(_03581_));
 XNOR2x1_ASAP7_75t_R _10412_ (.B(_03581_),
    .Y(_09950_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _10413_ (.A(_09950_),
    .Y(_09948_));
 NAND2x2_ASAP7_75t_R _10414_ (.A(_03393_),
    .B(net7),
    .Y(_03582_));
 AO21x1_ASAP7_75t_R _10415_ (.A1(_03506_),
    .A2(_03508_),
    .B(_03582_),
    .Y(_03583_));
 BUFx6f_ASAP7_75t_R _10416_ (.A(_03583_),
    .Y(_03584_));
 BUFx12_ASAP7_75t_R _10417_ (.A(_03584_),
    .Y(_03585_));
 BUFx10_ASAP7_75t_R _10418_ (.A(_03585_),
    .Y(_03586_));
 BUFx12_ASAP7_75t_R _10419_ (.A(_03586_),
    .Y(_03587_));
 INVx1_ASAP7_75t_R _10420_ (.A(_03493_),
    .Y(_03588_));
 OR4x1_ASAP7_75t_R _10421_ (.A(_03554_),
    .B(_00033_),
    .C(net65),
    .D(net95),
    .Y(_03589_));
 OR5x2_ASAP7_75t_R _10422_ (.A(_03511_),
    .B(_03512_),
    .C(_03513_),
    .D(_03588_),
    .E(_03589_),
    .Y(_03590_));
 BUFx12f_ASAP7_75t_R _10423_ (.A(instr[16]),
    .Y(_03591_));
 NAND2x2_ASAP7_75t_R _10424_ (.A(_03393_),
    .B(_03591_),
    .Y(_03592_));
 BUFx10_ASAP7_75t_R _10425_ (.A(_03592_),
    .Y(_03593_));
 NAND2x2_ASAP7_75t_R _10426_ (.A(_03373_),
    .B(net10),
    .Y(_03594_));
 INVx3_ASAP7_75t_R _10427_ (.A(net8),
    .Y(_03595_));
 INVx1_ASAP7_75t_R _10428_ (.A(net9),
    .Y(_03596_));
 AO21x2_ASAP7_75t_R _10429_ (.A1(_03595_),
    .A2(_03596_),
    .B(_03414_),
    .Y(_03597_));
 AND3x1_ASAP7_75t_R _10430_ (.A(_03593_),
    .B(_03594_),
    .C(_03597_),
    .Y(_03598_));
 AND2x4_ASAP7_75t_R _10431_ (.A(_03506_),
    .B(_03508_),
    .Y(_03599_));
 BUFx6f_ASAP7_75t_R _10432_ (.A(_03599_),
    .Y(_03600_));
 AO211x2_ASAP7_75t_R _10433_ (.A1(_03590_),
    .A2(_03598_),
    .B(_03600_),
    .C(_03572_),
    .Y(_03601_));
 NAND2x2_ASAP7_75t_R _10434_ (.A(_03587_),
    .B(_03601_),
    .Y(_03602_));
 AND4x2_ASAP7_75t_R _10435_ (.A(_03491_),
    .B(_03492_),
    .C(_03493_),
    .D(_03494_),
    .Y(_03603_));
 AND5x2_ASAP7_75t_R _10436_ (.A(_03510_),
    .B(_03490_),
    .C(_03486_),
    .D(_03489_),
    .E(_03603_),
    .Y(_03604_));
 BUFx6f_ASAP7_75t_R _10437_ (.A(_03604_),
    .Y(_03605_));
 BUFx12_ASAP7_75t_R _10438_ (.A(_03605_),
    .Y(_03606_));
 BUFx10_ASAP7_75t_R _10439_ (.A(_03593_),
    .Y(_03607_));
 BUFx12f_ASAP7_75t_R _10440_ (.A(net8),
    .Y(_03608_));
 BUFx12f_ASAP7_75t_R _10441_ (.A(_03608_),
    .Y(_03609_));
 BUFx12_ASAP7_75t_R _10442_ (.A(_03609_),
    .Y(_03610_));
 OA21x2_ASAP7_75t_R _10443_ (.A1(_03610_),
    .A2(net9),
    .B(_03549_),
    .Y(_03611_));
 BUFx16f_ASAP7_75t_R _10444_ (.A(_03582_),
    .Y(_03612_));
 BUFx12f_ASAP7_75t_R _10445_ (.A(net7),
    .Y(_03613_));
 BUFx16f_ASAP7_75t_R _10446_ (.A(_03613_),
    .Y(_03614_));
 AND3x1_ASAP7_75t_R _10447_ (.A(_00003_),
    .B(_03374_),
    .C(_03614_),
    .Y(_03615_));
 AO21x1_ASAP7_75t_R _10448_ (.A1(_00002_),
    .A2(_03612_),
    .B(_03615_),
    .Y(_03616_));
 OR4x1_ASAP7_75t_R _10449_ (.A(_03606_),
    .B(_03607_),
    .C(_03611_),
    .D(_03616_),
    .Y(_03617_));
 CKINVDCx5p33_ASAP7_75t_R _10450_ (.A(net7),
    .Y(_03618_));
 BUFx12f_ASAP7_75t_R _10451_ (.A(_03591_),
    .Y(_03619_));
 OR3x4_ASAP7_75t_R _10452_ (.A(_03414_),
    .B(_03618_),
    .C(_03619_),
    .Y(_03620_));
 OR4x1_ASAP7_75t_R _10453_ (.A(_00001_),
    .B(_03606_),
    .C(_03611_),
    .D(_03620_),
    .Y(_03621_));
 NAND3x1_ASAP7_75t_R _10454_ (.A(_03594_),
    .B(_03617_),
    .C(_03621_),
    .Y(_03622_));
 BUFx10_ASAP7_75t_R _10455_ (.A(_03402_),
    .Y(_03623_));
 BUFx12f_ASAP7_75t_R _10456_ (.A(_03614_),
    .Y(_03624_));
 INVx1_ASAP7_75t_R _10457_ (.A(_00006_),
    .Y(_03625_));
 AO21x1_ASAP7_75t_R _10458_ (.A1(_03623_),
    .A2(_03624_),
    .B(_03625_),
    .Y(_03626_));
 INVx1_ASAP7_75t_R _10459_ (.A(_00007_),
    .Y(_03627_));
 BUFx6f_ASAP7_75t_R _10460_ (.A(_03414_),
    .Y(_03628_));
 BUFx10_ASAP7_75t_R _10461_ (.A(_03618_),
    .Y(_03629_));
 OR3x1_ASAP7_75t_R _10462_ (.A(_03627_),
    .B(_03628_),
    .C(_03629_),
    .Y(_03630_));
 INVx2_ASAP7_75t_R _10463_ (.A(_03591_),
    .Y(_03631_));
 BUFx12_ASAP7_75t_R _10464_ (.A(_03631_),
    .Y(_03632_));
 BUFx12f_ASAP7_75t_R _10465_ (.A(_03613_),
    .Y(_03633_));
 AND2x2_ASAP7_75t_R _10466_ (.A(_00007_),
    .B(_03633_),
    .Y(_03634_));
 AO21x1_ASAP7_75t_R _10467_ (.A1(_00006_),
    .A2(_03618_),
    .B(_03634_),
    .Y(_03635_));
 BUFx12f_ASAP7_75t_R _10468_ (.A(_03591_),
    .Y(_03636_));
 OR3x1_ASAP7_75t_R _10469_ (.A(_00005_),
    .B(_03618_),
    .C(_03636_),
    .Y(_03637_));
 OAI21x1_ASAP7_75t_R _10470_ (.A1(_03632_),
    .A2(_03635_),
    .B(_03637_),
    .Y(_03638_));
 BUFx12_ASAP7_75t_R _10471_ (.A(_03395_),
    .Y(_03639_));
 AO32x1_ASAP7_75t_R _10472_ (.A1(_03606_),
    .A2(_03626_),
    .A3(_03630_),
    .B1(_03638_),
    .B2(_03639_),
    .Y(_03640_));
 INVx1_ASAP7_75t_R _10473_ (.A(_00004_),
    .Y(_03641_));
 NAND2x2_ASAP7_75t_R _10474_ (.A(_03510_),
    .B(_03490_),
    .Y(_03642_));
 OR5x1_ASAP7_75t_R _10475_ (.A(_03511_),
    .B(_03512_),
    .C(_03513_),
    .D(_03514_),
    .E(_03642_),
    .Y(_03643_));
 BUFx4f_ASAP7_75t_R _10476_ (.A(_03643_),
    .Y(_03644_));
 BUFx12_ASAP7_75t_R _10477_ (.A(_03644_),
    .Y(_03645_));
 BUFx12_ASAP7_75t_R _10478_ (.A(_03645_),
    .Y(_03646_));
 AO21x2_ASAP7_75t_R _10479_ (.A1(_03618_),
    .A2(_03631_),
    .B(_03414_),
    .Y(_03647_));
 BUFx12_ASAP7_75t_R _10480_ (.A(_03647_),
    .Y(_03648_));
 AND3x1_ASAP7_75t_R _10481_ (.A(_03641_),
    .B(_03646_),
    .C(_03648_),
    .Y(_03649_));
 NAND2x2_ASAP7_75t_R _10482_ (.A(_03373_),
    .B(_03608_),
    .Y(_03650_));
 AND2x6_ASAP7_75t_R _10483_ (.A(_03373_),
    .B(net9),
    .Y(_03651_));
 AOI21x1_ASAP7_75t_R _10484_ (.A1(_03644_),
    .A2(_03650_),
    .B(_03651_),
    .Y(_03652_));
 BUFx10_ASAP7_75t_R _10485_ (.A(_03652_),
    .Y(_03653_));
 OA21x2_ASAP7_75t_R _10486_ (.A1(_03640_),
    .A2(_03649_),
    .B(_03653_),
    .Y(_03654_));
 BUFx10_ASAP7_75t_R _10487_ (.A(_03518_),
    .Y(_03655_));
 OA21x2_ASAP7_75t_R _10488_ (.A1(_03622_),
    .A2(_03654_),
    .B(_03655_),
    .Y(_03656_));
 AND3x4_ASAP7_75t_R _10489_ (.A(_03486_),
    .B(_03489_),
    .C(_03603_),
    .Y(_03657_));
 AO221x2_ASAP7_75t_R _10490_ (.A1(_03554_),
    .A2(_03657_),
    .B1(_03570_),
    .B2(_03593_),
    .C(_03599_),
    .Y(_03658_));
 BUFx10_ASAP7_75t_R _10491_ (.A(_03658_),
    .Y(_03659_));
 BUFx12f_ASAP7_75t_R _10492_ (.A(_03645_),
    .Y(_03660_));
 BUFx10_ASAP7_75t_R _10493_ (.A(_03650_),
    .Y(_03661_));
 AND2x6_ASAP7_75t_R _10494_ (.A(_03660_),
    .B(_03661_),
    .Y(_03662_));
 BUFx12f_ASAP7_75t_R _10495_ (.A(_03549_),
    .Y(_03663_));
 BUFx16f_ASAP7_75t_R _10496_ (.A(_03633_),
    .Y(_03664_));
 BUFx16f_ASAP7_75t_R _10497_ (.A(_03664_),
    .Y(_03665_));
 AO32x1_ASAP7_75t_R _10498_ (.A1(_00011_),
    .A2(_03663_),
    .A3(_03665_),
    .B1(_03585_),
    .B2(_00010_),
    .Y(_03666_));
 BUFx12f_ASAP7_75t_R _10499_ (.A(_03605_),
    .Y(_03667_));
 AND2x4_ASAP7_75t_R _10500_ (.A(_03393_),
    .B(_03608_),
    .Y(_03668_));
 BUFx6f_ASAP7_75t_R _10501_ (.A(_03668_),
    .Y(_03669_));
 BUFx16f_ASAP7_75t_R _10502_ (.A(_03669_),
    .Y(_03670_));
 BUFx16f_ASAP7_75t_R _10503_ (.A(_03582_),
    .Y(_03671_));
 BUFx16f_ASAP7_75t_R _10504_ (.A(_03613_),
    .Y(_03672_));
 AND3x1_ASAP7_75t_R _10505_ (.A(_00015_),
    .B(_03395_),
    .C(_03672_),
    .Y(_03673_));
 AO21x1_ASAP7_75t_R _10506_ (.A1(_00014_),
    .A2(_03671_),
    .B(_03673_),
    .Y(_03674_));
 OA21x2_ASAP7_75t_R _10507_ (.A1(_03667_),
    .A2(_03670_),
    .B(_03674_),
    .Y(_03675_));
 AOI21x1_ASAP7_75t_R _10508_ (.A1(_03662_),
    .A2(_03666_),
    .B(_03675_),
    .Y(_03676_));
 BUFx6f_ASAP7_75t_R _10509_ (.A(_03509_),
    .Y(_03677_));
 BUFx10_ASAP7_75t_R _10510_ (.A(_03516_),
    .Y(_03678_));
 BUFx12_ASAP7_75t_R _10511_ (.A(_03604_),
    .Y(_03679_));
 AND2x6_ASAP7_75t_R _10512_ (.A(_03373_),
    .B(_03591_),
    .Y(_03680_));
 BUFx12f_ASAP7_75t_R _10513_ (.A(_03680_),
    .Y(_03681_));
 INVx1_ASAP7_75t_R _10514_ (.A(_00009_),
    .Y(_03682_));
 BUFx12f_ASAP7_75t_R _10515_ (.A(_03595_),
    .Y(_03683_));
 AND3x1_ASAP7_75t_R _10516_ (.A(_03682_),
    .B(_03633_),
    .C(_03683_),
    .Y(_03684_));
 BUFx12_ASAP7_75t_R _10517_ (.A(_03608_),
    .Y(_03685_));
 NAND2x1_ASAP7_75t_R _10518_ (.A(_00013_),
    .B(_03613_),
    .Y(_03686_));
 OA211x2_ASAP7_75t_R _10519_ (.A1(_03433_),
    .A2(_03633_),
    .B(_03685_),
    .C(_03686_),
    .Y(_03687_));
 OA21x2_ASAP7_75t_R _10520_ (.A1(_03684_),
    .A2(_03687_),
    .B(_03443_),
    .Y(_03688_));
 OR3x1_ASAP7_75t_R _10521_ (.A(_03679_),
    .B(_03681_),
    .C(_03688_),
    .Y(_03689_));
 OR2x6_ASAP7_75t_R _10522_ (.A(net7),
    .B(net8),
    .Y(_03690_));
 NAND2x2_ASAP7_75t_R _10523_ (.A(_03394_),
    .B(_03690_),
    .Y(_03691_));
 AO211x2_ASAP7_75t_R _10524_ (.A1(_03590_),
    .A2(_03691_),
    .B(_03599_),
    .C(_03572_),
    .Y(_03692_));
 INVx1_ASAP7_75t_R _10525_ (.A(_00008_),
    .Y(_03693_));
 AO32x1_ASAP7_75t_R _10526_ (.A1(_03677_),
    .A2(_03678_),
    .A3(_03689_),
    .B1(_03692_),
    .B2(_03693_),
    .Y(_03694_));
 OR4x2_ASAP7_75t_R _10527_ (.A(_01159_),
    .B(_03567_),
    .C(net27),
    .D(_03529_),
    .Y(_03695_));
 BUFx6f_ASAP7_75t_R _10528_ (.A(_03695_),
    .Y(_03696_));
 OA21x2_ASAP7_75t_R _10529_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03651_),
    .Y(_03697_));
 BUFx12f_ASAP7_75t_R _10530_ (.A(_03697_),
    .Y(_03698_));
 OA211x2_ASAP7_75t_R _10531_ (.A1(_03659_),
    .A2(_03676_),
    .B(_03694_),
    .C(_03698_),
    .Y(_03699_));
 INVx2_ASAP7_75t_R _10532_ (.A(_00000_),
    .Y(_01222_));
 AO221x2_ASAP7_75t_R _10533_ (.A1(_03554_),
    .A2(_03657_),
    .B1(_03590_),
    .B2(_03597_),
    .C(_03599_),
    .Y(_03700_));
 BUFx10_ASAP7_75t_R _10534_ (.A(_03700_),
    .Y(_03701_));
 AO221x2_ASAP7_75t_R _10535_ (.A1(_03554_),
    .A2(_03657_),
    .B1(_03590_),
    .B2(_03647_),
    .C(_03599_),
    .Y(_03702_));
 BUFx6f_ASAP7_75t_R _10536_ (.A(_03702_),
    .Y(_03703_));
 AND3x1_ASAP7_75t_R _10537_ (.A(_01222_),
    .B(_03701_),
    .C(_03703_),
    .Y(_03704_));
 BUFx10_ASAP7_75t_R _10538_ (.A(_03646_),
    .Y(_03705_));
 OR3x1_ASAP7_75t_R _10539_ (.A(_03414_),
    .B(_03631_),
    .C(_03683_),
    .Y(_03706_));
 BUFx10_ASAP7_75t_R _10540_ (.A(_03706_),
    .Y(_03707_));
 NAND2x1_ASAP7_75t_R _10541_ (.A(_03705_),
    .B(_03707_),
    .Y(_03708_));
 BUFx12_ASAP7_75t_R _10542_ (.A(_03582_),
    .Y(_03709_));
 BUFx12_ASAP7_75t_R _10543_ (.A(_03709_),
    .Y(_03710_));
 BUFx12_ASAP7_75t_R _10544_ (.A(_03710_),
    .Y(_03711_));
 AND3x1_ASAP7_75t_R _10545_ (.A(_00023_),
    .B(_03663_),
    .C(_03665_),
    .Y(_03712_));
 AOI211x1_ASAP7_75t_R _10546_ (.A1(_00022_),
    .A2(_03711_),
    .B(_03651_),
    .C(_03712_),
    .Y(_03713_));
 BUFx12f_ASAP7_75t_R _10547_ (.A(_03710_),
    .Y(_03714_));
 BUFx12_ASAP7_75t_R _10548_ (.A(_03443_),
    .Y(_03715_));
 BUFx12f_ASAP7_75t_R _10549_ (.A(_03633_),
    .Y(_03716_));
 BUFx16f_ASAP7_75t_R _10550_ (.A(_03716_),
    .Y(_03717_));
 AND3x1_ASAP7_75t_R _10551_ (.A(_03471_),
    .B(_03715_),
    .C(_03717_),
    .Y(_03718_));
 AO21x1_ASAP7_75t_R _10552_ (.A1(_03468_),
    .A2(_03714_),
    .B(_03718_),
    .Y(_03719_));
 AND3x1_ASAP7_75t_R _10553_ (.A(_03596_),
    .B(_03592_),
    .C(_03668_),
    .Y(_03720_));
 AND2x6_ASAP7_75t_R _10554_ (.A(_03509_),
    .B(_03720_),
    .Y(_03721_));
 AO21x2_ASAP7_75t_R _10555_ (.A1(_03506_),
    .A2(_03508_),
    .B(_03594_),
    .Y(_03722_));
 BUFx10_ASAP7_75t_R _10556_ (.A(_03722_),
    .Y(_03723_));
 AO221x1_ASAP7_75t_R _10557_ (.A1(_03708_),
    .A2(_03713_),
    .B1(_03719_),
    .B2(_03721_),
    .C(_03723_),
    .Y(_03724_));
 NAND2x1_ASAP7_75t_R _10558_ (.A(_00026_),
    .B(_03585_),
    .Y(_03725_));
 AND2x2_ASAP7_75t_R _10559_ (.A(_03393_),
    .B(net7),
    .Y(_03726_));
 BUFx12_ASAP7_75t_R _10560_ (.A(_03726_),
    .Y(_03727_));
 BUFx12f_ASAP7_75t_R _10561_ (.A(_03727_),
    .Y(_03728_));
 NAND2x1_ASAP7_75t_R _10562_ (.A(_00027_),
    .B(_03728_),
    .Y(_03729_));
 AND4x1_ASAP7_75t_R _10563_ (.A(_03662_),
    .B(_03697_),
    .C(_03725_),
    .D(_03729_),
    .Y(_03730_));
 AO32x2_ASAP7_75t_R _10564_ (.A1(_03486_),
    .A2(_03489_),
    .A3(_03495_),
    .B1(_03591_),
    .B2(_03373_),
    .Y(_03731_));
 AND3x1_ASAP7_75t_R _10565_ (.A(_03509_),
    .B(_03557_),
    .C(_03731_),
    .Y(_03732_));
 BUFx12_ASAP7_75t_R _10566_ (.A(_03732_),
    .Y(_03733_));
 BUFx10_ASAP7_75t_R _10567_ (.A(_03650_),
    .Y(_03734_));
 BUFx12f_ASAP7_75t_R _10568_ (.A(_03734_),
    .Y(_03735_));
 BUFx6f_ASAP7_75t_R _10569_ (.A(_03644_),
    .Y(_03736_));
 BUFx12f_ASAP7_75t_R _10570_ (.A(_03736_),
    .Y(_03737_));
 AND2x2_ASAP7_75t_R _10571_ (.A(_00030_),
    .B(_03671_),
    .Y(_03738_));
 AO221x1_ASAP7_75t_R _10572_ (.A1(_00031_),
    .A2(_03728_),
    .B1(_03735_),
    .B2(_03737_),
    .C(_03738_),
    .Y(_03739_));
 NAND2x2_ASAP7_75t_R _10573_ (.A(_03509_),
    .B(_03651_),
    .Y(_03740_));
 AOI21x1_ASAP7_75t_R _10574_ (.A1(_03733_),
    .A2(_03739_),
    .B(_03740_),
    .Y(_03741_));
 BUFx10_ASAP7_75t_R _10575_ (.A(_03677_),
    .Y(_03742_));
 INVx1_ASAP7_75t_R _10576_ (.A(_00025_),
    .Y(_03743_));
 BUFx16f_ASAP7_75t_R _10577_ (.A(_03595_),
    .Y(_03744_));
 AND3x1_ASAP7_75t_R _10578_ (.A(_03743_),
    .B(_03614_),
    .C(_03744_),
    .Y(_03745_));
 NAND2x1_ASAP7_75t_R _10579_ (.A(_00029_),
    .B(_03613_),
    .Y(_03746_));
 OA211x2_ASAP7_75t_R _10580_ (.A1(_03436_),
    .A2(_03633_),
    .B(_03609_),
    .C(_03746_),
    .Y(_03747_));
 OA21x2_ASAP7_75t_R _10581_ (.A1(_03745_),
    .A2(_03747_),
    .B(_03623_),
    .Y(_03748_));
 OR3x1_ASAP7_75t_R _10582_ (.A(_03606_),
    .B(_03681_),
    .C(_03748_),
    .Y(_03749_));
 BUFx12_ASAP7_75t_R _10583_ (.A(_03692_),
    .Y(_03750_));
 INVx1_ASAP7_75t_R _10584_ (.A(_00024_),
    .Y(_03751_));
 AO32x1_ASAP7_75t_R _10585_ (.A1(_03742_),
    .A2(_03678_),
    .A3(_03749_),
    .B1(_03750_),
    .B2(_03751_),
    .Y(_03752_));
 OA21x2_ASAP7_75t_R _10586_ (.A1(_03730_),
    .A2(_03741_),
    .B(_03752_),
    .Y(_03753_));
 AND2x2_ASAP7_75t_R _10587_ (.A(_03491_),
    .B(_03492_),
    .Y(_03754_));
 AND4x1_ASAP7_75t_R _10588_ (.A(_03510_),
    .B(_03490_),
    .C(_03493_),
    .D(_03494_),
    .Y(_03755_));
 AND4x2_ASAP7_75t_R _10589_ (.A(_03486_),
    .B(_03489_),
    .C(_03754_),
    .D(_03755_),
    .Y(_03756_));
 NAND2x2_ASAP7_75t_R _10590_ (.A(_03582_),
    .B(_03592_),
    .Y(_03757_));
 OA211x2_ASAP7_75t_R _10591_ (.A1(_03756_),
    .A2(_03757_),
    .B(_03509_),
    .C(_03557_),
    .Y(_03758_));
 BUFx12f_ASAP7_75t_R _10592_ (.A(_03758_),
    .Y(_03759_));
 NOR2x1_ASAP7_75t_R _10593_ (.A(_00016_),
    .B(_03759_),
    .Y(_03760_));
 BUFx12_ASAP7_75t_R _10594_ (.A(_03671_),
    .Y(_03761_));
 BUFx16f_ASAP7_75t_R _10595_ (.A(_03672_),
    .Y(_03762_));
 AND3x1_ASAP7_75t_R _10596_ (.A(_00019_),
    .B(_03639_),
    .C(_03762_),
    .Y(_03763_));
 AO21x1_ASAP7_75t_R _10597_ (.A1(_00018_),
    .A2(_03761_),
    .B(_03763_),
    .Y(_03764_));
 BUFx10_ASAP7_75t_R _10598_ (.A(_03680_),
    .Y(_03765_));
 OR4x1_ASAP7_75t_R _10599_ (.A(_00017_),
    .B(_03606_),
    .C(_03585_),
    .D(_03765_),
    .Y(_03766_));
 OAI21x1_ASAP7_75t_R _10600_ (.A1(_03659_),
    .A2(_03764_),
    .B(_03766_),
    .Y(_03767_));
 OA21x2_ASAP7_75t_R _10601_ (.A1(_03760_),
    .A2(_03767_),
    .B(_03701_),
    .Y(_03768_));
 OA33x2_ASAP7_75t_R _10602_ (.A1(_03656_),
    .A2(_03699_),
    .A3(_03704_),
    .B1(_03724_),
    .B2(_03753_),
    .B3(_03768_),
    .Y(_03769_));
 BUFx6f_ASAP7_75t_R _10603_ (.A(_03769_),
    .Y(_03770_));
 AND2x4_ASAP7_75t_R _10604_ (.A(_03602_),
    .B(_03770_),
    .Y(_09949_));
 BUFx10_ASAP7_75t_R _10605_ (.A(_03597_),
    .Y(_03771_));
 AND2x6_ASAP7_75t_R _10606_ (.A(_03645_),
    .B(_03771_),
    .Y(_03772_));
 BUFx12f_ASAP7_75t_R _10607_ (.A(_03772_),
    .Y(_03773_));
 BUFx6f_ASAP7_75t_R _10608_ (.A(_03728_),
    .Y(_03774_));
 BUFx12f_ASAP7_75t_R _10609_ (.A(_03593_),
    .Y(_03775_));
 BUFx12f_ASAP7_75t_R _10610_ (.A(_03775_),
    .Y(_03776_));
 BUFx12_ASAP7_75t_R _10611_ (.A(_03737_),
    .Y(_03777_));
 AND2x2_ASAP7_75t_R _10612_ (.A(_00053_),
    .B(_03761_),
    .Y(_03778_));
 AO221x1_ASAP7_75t_R _10613_ (.A1(_00054_),
    .A2(_03774_),
    .B1(_03776_),
    .B2(_03777_),
    .C(_03778_),
    .Y(_03779_));
 BUFx12_ASAP7_75t_R _10614_ (.A(_03679_),
    .Y(_03780_));
 BUFx16f_ASAP7_75t_R _10615_ (.A(_03612_),
    .Y(_03781_));
 BUFx12_ASAP7_75t_R _10616_ (.A(_03781_),
    .Y(_03782_));
 BUFx10_ASAP7_75t_R _10617_ (.A(_03681_),
    .Y(_03783_));
 OR4x1_ASAP7_75t_R _10618_ (.A(_00052_),
    .B(_03780_),
    .C(_03782_),
    .D(_03783_),
    .Y(_03784_));
 BUFx16f_ASAP7_75t_R _10619_ (.A(_03539_),
    .Y(_03785_));
 BUFx12f_ASAP7_75t_R _10620_ (.A(_03785_),
    .Y(_03786_));
 AO31x2_ASAP7_75t_R _10621_ (.A1(_03773_),
    .A2(_03779_),
    .A3(_03784_),
    .B(_03786_),
    .Y(_03787_));
 INVx2_ASAP7_75t_R _10622_ (.A(_00051_),
    .Y(_03788_));
 NAND2x1_ASAP7_75t_R _10623_ (.A(_03788_),
    .B(_03703_),
    .Y(_03789_));
 AND2x2_ASAP7_75t_R _10624_ (.A(_03517_),
    .B(_03652_),
    .Y(_03790_));
 BUFx12f_ASAP7_75t_R _10625_ (.A(_03790_),
    .Y(_03791_));
 BUFx12f_ASAP7_75t_R _10626_ (.A(_03791_),
    .Y(_03792_));
 NAND2x1_ASAP7_75t_R _10627_ (.A(_03644_),
    .B(_03592_),
    .Y(_03793_));
 BUFx10_ASAP7_75t_R _10628_ (.A(_03793_),
    .Y(_03794_));
 BUFx10_ASAP7_75t_R _10629_ (.A(_03794_),
    .Y(_03795_));
 BUFx12_ASAP7_75t_R _10630_ (.A(_03714_),
    .Y(_03796_));
 BUFx10_ASAP7_75t_R _10631_ (.A(_03715_),
    .Y(_03797_));
 BUFx12f_ASAP7_75t_R _10632_ (.A(_03717_),
    .Y(_03798_));
 AND3x1_ASAP7_75t_R _10633_ (.A(_03797_),
    .B(_03798_),
    .C(_00056_),
    .Y(_03799_));
 AO21x1_ASAP7_75t_R _10634_ (.A1(_00055_),
    .A2(_03796_),
    .B(_03799_),
    .Y(_03800_));
 BUFx10_ASAP7_75t_R _10635_ (.A(_03593_),
    .Y(_03801_));
 BUFx12f_ASAP7_75t_R _10636_ (.A(_03801_),
    .Y(_03802_));
 BUFx10_ASAP7_75t_R _10637_ (.A(_03802_),
    .Y(_03803_));
 BUFx10_ASAP7_75t_R _10638_ (.A(_03737_),
    .Y(_03804_));
 BUFx6f_ASAP7_75t_R _10639_ (.A(_03710_),
    .Y(_03805_));
 AND2x2_ASAP7_75t_R _10640_ (.A(_00057_),
    .B(_03805_),
    .Y(_03806_));
 AO221x1_ASAP7_75t_R _10641_ (.A1(_00058_),
    .A2(_03774_),
    .B1(_03803_),
    .B2(_03804_),
    .C(_03806_),
    .Y(_03807_));
 OA21x2_ASAP7_75t_R _10642_ (.A1(_03795_),
    .A2(_03800_),
    .B(_03807_),
    .Y(_03808_));
 BUFx6f_ASAP7_75t_R _10643_ (.A(_03723_),
    .Y(_03809_));
 AO221x1_ASAP7_75t_R _10644_ (.A1(_03787_),
    .A2(_03789_),
    .B1(_03792_),
    .B2(_03808_),
    .C(_03809_),
    .Y(_03810_));
 BUFx12_ASAP7_75t_R _10645_ (.A(_03750_),
    .Y(_03811_));
 AND2x2_ASAP7_75t_R _10646_ (.A(_00059_),
    .B(_03811_),
    .Y(_03812_));
 OA21x2_ASAP7_75t_R _10647_ (.A1(_03522_),
    .A2(_03696_),
    .B(_03727_),
    .Y(_03813_));
 BUFx12_ASAP7_75t_R _10648_ (.A(_03813_),
    .Y(_03814_));
 BUFx12f_ASAP7_75t_R _10649_ (.A(_03663_),
    .Y(_03815_));
 BUFx6f_ASAP7_75t_R _10650_ (.A(_03636_),
    .Y(_03816_));
 BUFx6f_ASAP7_75t_R _10651_ (.A(_03670_),
    .Y(_03817_));
 AND3x1_ASAP7_75t_R _10652_ (.A(_03639_),
    .B(_03762_),
    .C(_00064_),
    .Y(_03818_));
 AO21x1_ASAP7_75t_R _10653_ (.A1(_00063_),
    .A2(_03805_),
    .B(_03818_),
    .Y(_03819_));
 BUFx12_ASAP7_75t_R _10654_ (.A(_03667_),
    .Y(_03820_));
 AO221x1_ASAP7_75t_R _10655_ (.A1(_03815_),
    .A2(_03816_),
    .B1(_03817_),
    .B2(_03819_),
    .C(_03820_),
    .Y(_03821_));
 BUFx12f_ASAP7_75t_R _10656_ (.A(_03518_),
    .Y(_03822_));
 AO32x1_ASAP7_75t_R _10657_ (.A1(_00060_),
    .A2(_03814_),
    .A3(_03662_),
    .B1(_03821_),
    .B2(_03822_),
    .Y(_03823_));
 AND2x6_ASAP7_75t_R _10658_ (.A(_03644_),
    .B(_03592_),
    .Y(_03824_));
 BUFx12f_ASAP7_75t_R _10659_ (.A(_03824_),
    .Y(_03825_));
 BUFx10_ASAP7_75t_R _10660_ (.A(_03825_),
    .Y(_03826_));
 BUFx12_ASAP7_75t_R _10661_ (.A(_03644_),
    .Y(_03827_));
 BUFx12f_ASAP7_75t_R _10662_ (.A(_03827_),
    .Y(_03828_));
 BUFx10_ASAP7_75t_R _10663_ (.A(_03828_),
    .Y(_03829_));
 BUFx12f_ASAP7_75t_R _10664_ (.A(_03691_),
    .Y(_03830_));
 BUFx6f_ASAP7_75t_R _10665_ (.A(_03830_),
    .Y(_03831_));
 AND3x1_ASAP7_75t_R _10666_ (.A(_00061_),
    .B(_03829_),
    .C(_03831_),
    .Y(_03832_));
 AND3x4_ASAP7_75t_R _10667_ (.A(_03395_),
    .B(_03672_),
    .C(_03744_),
    .Y(_03833_));
 BUFx10_ASAP7_75t_R _10668_ (.A(_03833_),
    .Y(_03834_));
 AND2x2_ASAP7_75t_R _10669_ (.A(_00062_),
    .B(_03834_),
    .Y(_03835_));
 BUFx12f_ASAP7_75t_R _10670_ (.A(_03660_),
    .Y(_03836_));
 BUFx10_ASAP7_75t_R _10671_ (.A(_03836_),
    .Y(_03837_));
 BUFx12f_ASAP7_75t_R _10672_ (.A(_03735_),
    .Y(_03838_));
 BUFx12_ASAP7_75t_R _10673_ (.A(_03419_),
    .Y(_03839_));
 BUFx10_ASAP7_75t_R _10674_ (.A(_03629_),
    .Y(_03840_));
 INVx1_ASAP7_75t_R _10675_ (.A(_00066_),
    .Y(_03841_));
 OR3x1_ASAP7_75t_R _10676_ (.A(_03839_),
    .B(_03840_),
    .C(_03841_),
    .Y(_03842_));
 BUFx16f_ASAP7_75t_R _10677_ (.A(_03374_),
    .Y(_03843_));
 BUFx10_ASAP7_75t_R _10678_ (.A(_03843_),
    .Y(_03844_));
 BUFx12_ASAP7_75t_R _10679_ (.A(_03762_),
    .Y(_03845_));
 INVx1_ASAP7_75t_R _10680_ (.A(_00065_),
    .Y(_03846_));
 AO21x1_ASAP7_75t_R _10681_ (.A1(_03844_),
    .A2(_03845_),
    .B(_03846_),
    .Y(_03847_));
 AOI22x1_ASAP7_75t_R _10682_ (.A1(_03837_),
    .A2(_03838_),
    .B1(_03842_),
    .B2(_03847_),
    .Y(_03848_));
 OR4x1_ASAP7_75t_R _10683_ (.A(_03826_),
    .B(_03832_),
    .C(_03835_),
    .D(_03848_),
    .Y(_03849_));
 BUFx6f_ASAP7_75t_R _10684_ (.A(_03698_),
    .Y(_03850_));
 OA211x2_ASAP7_75t_R _10685_ (.A1(_03812_),
    .A2(_03823_),
    .B(_03849_),
    .C(_03850_),
    .Y(_03851_));
 BUFx12f_ASAP7_75t_R _10686_ (.A(_03794_),
    .Y(_03852_));
 BUFx10_ASAP7_75t_R _10687_ (.A(_03664_),
    .Y(_03853_));
 AND3x1_ASAP7_75t_R _10688_ (.A(_03663_),
    .B(_03853_),
    .C(_00048_),
    .Y(_03854_));
 AO21x1_ASAP7_75t_R _10689_ (.A1(_00047_),
    .A2(_03711_),
    .B(_03854_),
    .Y(_03855_));
 AND2x2_ASAP7_75t_R _10690_ (.A(_03817_),
    .B(_03855_),
    .Y(_03856_));
 OA21x2_ASAP7_75t_R _10691_ (.A1(_03852_),
    .A2(_03856_),
    .B(_03822_),
    .Y(_03857_));
 AO32x1_ASAP7_75t_R _10692_ (.A1(_00044_),
    .A2(_03814_),
    .A3(_03662_),
    .B1(_03811_),
    .B2(_00043_),
    .Y(_03858_));
 OR3x1_ASAP7_75t_R _10693_ (.A(_00045_),
    .B(_03820_),
    .C(_03817_),
    .Y(_03859_));
 BUFx6f_ASAP7_75t_R _10694_ (.A(_03645_),
    .Y(_03860_));
 BUFx12f_ASAP7_75t_R _10695_ (.A(_03860_),
    .Y(_03861_));
 BUFx12f_ASAP7_75t_R _10696_ (.A(_03861_),
    .Y(_03862_));
 AO21x1_ASAP7_75t_R _10697_ (.A1(_03862_),
    .A2(_03838_),
    .B(_00049_),
    .Y(_03863_));
 AO21x2_ASAP7_75t_R _10698_ (.A1(_03590_),
    .A2(_03592_),
    .B(_03726_),
    .Y(_03864_));
 BUFx10_ASAP7_75t_R _10699_ (.A(_03864_),
    .Y(_03865_));
 BUFx16f_ASAP7_75t_R _10700_ (.A(_03865_),
    .Y(_03866_));
 AO21x1_ASAP7_75t_R _10701_ (.A1(_03859_),
    .A2(_03863_),
    .B(_03866_),
    .Y(_03867_));
 BUFx12_ASAP7_75t_R _10702_ (.A(_03697_),
    .Y(_03868_));
 OR3x4_ASAP7_75t_R _10703_ (.A(_03415_),
    .B(_03629_),
    .C(_03632_),
    .Y(_03869_));
 AND3x1_ASAP7_75t_R _10704_ (.A(_00050_),
    .B(_03742_),
    .C(_03651_),
    .Y(_03870_));
 NAND2x2_ASAP7_75t_R _10705_ (.A(_03645_),
    .B(_03650_),
    .Y(_03871_));
 BUFx16f_ASAP7_75t_R _10706_ (.A(_03871_),
    .Y(_03872_));
 BUFx6f_ASAP7_75t_R _10707_ (.A(_03646_),
    .Y(_03873_));
 BUFx10_ASAP7_75t_R _10708_ (.A(_03661_),
    .Y(_03874_));
 AND5x1_ASAP7_75t_R _10709_ (.A(_00046_),
    .B(_03742_),
    .C(_03873_),
    .D(_03651_),
    .E(_03874_),
    .Y(_03875_));
 AO221x1_ASAP7_75t_R _10710_ (.A1(_03868_),
    .A2(_03869_),
    .B1(_03870_),
    .B2(_03872_),
    .C(_03875_),
    .Y(_03876_));
 OA211x2_ASAP7_75t_R _10711_ (.A1(_03857_),
    .A2(_03858_),
    .B(_03867_),
    .C(_03876_),
    .Y(_03877_));
 BUFx12f_ASAP7_75t_R _10712_ (.A(_03584_),
    .Y(_03878_));
 BUFx12f_ASAP7_75t_R _10713_ (.A(_03878_),
    .Y(_03879_));
 BUFx10_ASAP7_75t_R _10714_ (.A(_03696_),
    .Y(_03880_));
 BUFx16f_ASAP7_75t_R _10715_ (.A(_03727_),
    .Y(_03881_));
 BUFx12_ASAP7_75t_R _10716_ (.A(_03881_),
    .Y(_03882_));
 OA211x2_ASAP7_75t_R _10717_ (.A1(_03524_),
    .A2(_03880_),
    .B(_03882_),
    .C(_00040_),
    .Y(_03883_));
 AO21x1_ASAP7_75t_R _10718_ (.A1(_00039_),
    .A2(_03879_),
    .B(_03883_),
    .Y(_03884_));
 BUFx12_ASAP7_75t_R _10719_ (.A(_03726_),
    .Y(_03885_));
 BUFx12f_ASAP7_75t_R _10720_ (.A(_03885_),
    .Y(_03886_));
 BUFx12_ASAP7_75t_R _10721_ (.A(_03886_),
    .Y(_03887_));
 BUFx12f_ASAP7_75t_R _10722_ (.A(_03801_),
    .Y(_03888_));
 BUFx12f_ASAP7_75t_R _10723_ (.A(_03888_),
    .Y(_03889_));
 BUFx12f_ASAP7_75t_R _10724_ (.A(_03612_),
    .Y(_03890_));
 BUFx12f_ASAP7_75t_R _10725_ (.A(_03890_),
    .Y(_03891_));
 AND2x2_ASAP7_75t_R _10726_ (.A(_00041_),
    .B(_03891_),
    .Y(_03892_));
 AO221x1_ASAP7_75t_R _10727_ (.A1(_00042_),
    .A2(_03887_),
    .B1(_03889_),
    .B2(_03862_),
    .C(_03892_),
    .Y(_03893_));
 OA21x2_ASAP7_75t_R _10728_ (.A1(_03852_),
    .A2(_03884_),
    .B(_03893_),
    .Y(_03894_));
 INVx1_ASAP7_75t_R _10729_ (.A(_00038_),
    .Y(_03895_));
 NAND2x1_ASAP7_75t_R _10730_ (.A(_03895_),
    .B(_03814_),
    .Y(_03896_));
 BUFx12f_ASAP7_75t_R _10731_ (.A(_03619_),
    .Y(_03897_));
 INVx1_ASAP7_75t_R _10732_ (.A(net10),
    .Y(_03898_));
 AND3x1_ASAP7_75t_R _10733_ (.A(_03395_),
    .B(_03897_),
    .C(_03898_),
    .Y(_03899_));
 OA211x2_ASAP7_75t_R _10734_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03771_),
    .C(_03899_),
    .Y(_03900_));
 BUFx6f_ASAP7_75t_R _10735_ (.A(_03900_),
    .Y(_03901_));
 OA21x2_ASAP7_75t_R _10736_ (.A1(_00037_),
    .A2(_03887_),
    .B(_03901_),
    .Y(_03902_));
 INVx2_ASAP7_75t_R _10737_ (.A(_00036_),
    .Y(_03903_));
 NAND2x1_ASAP7_75t_R _10738_ (.A(_03903_),
    .B(_03814_),
    .Y(_03904_));
 AND2x4_ASAP7_75t_R _10739_ (.A(_03393_),
    .B(net10),
    .Y(_03905_));
 OA21x2_ASAP7_75t_R _10740_ (.A1(_03522_),
    .A2(_03695_),
    .B(_03905_),
    .Y(_03906_));
 BUFx6f_ASAP7_75t_R _10741_ (.A(_03906_),
    .Y(_03907_));
 AO221x1_ASAP7_75t_R _10742_ (.A1(_03896_),
    .A2(_03902_),
    .B1(_03904_),
    .B2(_03601_),
    .C(_03907_),
    .Y(_03908_));
 AO21x1_ASAP7_75t_R _10743_ (.A1(_03792_),
    .A2(_03894_),
    .B(_03908_),
    .Y(_03909_));
 OA22x2_ASAP7_75t_R _10744_ (.A1(_03810_),
    .A2(_03851_),
    .B1(_03877_),
    .B2(_03909_),
    .Y(_03910_));
 INVx3_ASAP7_75t_R _10745_ (.A(_03910_),
    .Y(_03911_));
 BUFx4f_ASAP7_75t_R _10746_ (.A(_03911_),
    .Y(_09953_));
 OR2x2_ASAP7_75t_R _10747_ (.A(_03527_),
    .B(_03536_),
    .Y(_03912_));
 BUFx12_ASAP7_75t_R _10748_ (.A(_03912_),
    .Y(_03913_));
 BUFx12_ASAP7_75t_R _10749_ (.A(_03913_),
    .Y(_03914_));
 BUFx6f_ASAP7_75t_R _10750_ (.A(_03575_),
    .Y(_03915_));
 BUFx10_ASAP7_75t_R _10751_ (.A(_03384_),
    .Y(_03916_));
 BUFx10_ASAP7_75t_R _10752_ (.A(_03916_),
    .Y(_03917_));
 AND2x2_ASAP7_75t_R _10753_ (.A(_03442_),
    .B(_03375_),
    .Y(_03918_));
 BUFx10_ASAP7_75t_R _10754_ (.A(_03918_),
    .Y(_03919_));
 BUFx10_ASAP7_75t_R _10755_ (.A(_03919_),
    .Y(_03920_));
 BUFx10_ASAP7_75t_R _10756_ (.A(_03920_),
    .Y(_03921_));
 BUFx6f_ASAP7_75t_R _10757_ (.A(_03392_),
    .Y(_03922_));
 BUFx6f_ASAP7_75t_R _10758_ (.A(_03922_),
    .Y(_03923_));
 BUFx6f_ASAP7_75t_R _10759_ (.A(_03923_),
    .Y(_03924_));
 BUFx12_ASAP7_75t_R _10760_ (.A(_03924_),
    .Y(_03925_));
 BUFx12f_ASAP7_75t_R _10761_ (.A(_03925_),
    .Y(_03926_));
 BUFx10_ASAP7_75t_R _10762_ (.A(_03926_),
    .Y(_03927_));
 BUFx12_ASAP7_75t_R _10763_ (.A(_03423_),
    .Y(_03928_));
 BUFx10_ASAP7_75t_R _10764_ (.A(_03928_),
    .Y(_03929_));
 BUFx12f_ASAP7_75t_R _10765_ (.A(_03929_),
    .Y(_03930_));
 BUFx6f_ASAP7_75t_R _10766_ (.A(_03400_),
    .Y(_03931_));
 BUFx6f_ASAP7_75t_R _10767_ (.A(_03931_),
    .Y(_03932_));
 BUFx6f_ASAP7_75t_R _10768_ (.A(_03932_),
    .Y(_03933_));
 AND2x2_ASAP7_75t_R _10769_ (.A(_03933_),
    .B(_00050_),
    .Y(_03934_));
 AO21x1_ASAP7_75t_R _10770_ (.A1(_03930_),
    .A2(_00049_),
    .B(_03934_),
    .Y(_03935_));
 NAND2x2_ASAP7_75t_R _10771_ (.A(_03922_),
    .B(_03715_),
    .Y(_03936_));
 BUFx10_ASAP7_75t_R _10772_ (.A(_03936_),
    .Y(_03937_));
 BUFx6f_ASAP7_75t_R _10773_ (.A(_03937_),
    .Y(_03938_));
 BUFx6f_ASAP7_75t_R _10774_ (.A(_03548_),
    .Y(_03939_));
 BUFx6f_ASAP7_75t_R _10775_ (.A(_03931_),
    .Y(_03940_));
 BUFx12_ASAP7_75t_R _10776_ (.A(_03940_),
    .Y(_03941_));
 BUFx10_ASAP7_75t_R _10777_ (.A(_03941_),
    .Y(_03942_));
 BUFx10_ASAP7_75t_R _10778_ (.A(_03378_),
    .Y(_03943_));
 AND3x1_ASAP7_75t_R _10779_ (.A(_03942_),
    .B(_03943_),
    .C(_00048_),
    .Y(_03944_));
 AO21x1_ASAP7_75t_R _10780_ (.A1(_00047_),
    .A2(_03939_),
    .B(_03944_),
    .Y(_03945_));
 BUFx6f_ASAP7_75t_R _10781_ (.A(_03449_),
    .Y(_03946_));
 BUFx6f_ASAP7_75t_R _10782_ (.A(_03946_),
    .Y(_03947_));
 AO221x2_ASAP7_75t_R _10783_ (.A1(_03927_),
    .A2(_03935_),
    .B1(_03938_),
    .B2(_03945_),
    .C(_03947_),
    .Y(_03948_));
 BUFx10_ASAP7_75t_R _10784_ (.A(_03928_),
    .Y(_03949_));
 BUFx6f_ASAP7_75t_R _10785_ (.A(_03949_),
    .Y(_03950_));
 BUFx12_ASAP7_75t_R _10786_ (.A(_03950_),
    .Y(_03951_));
 BUFx6f_ASAP7_75t_R _10787_ (.A(_03424_),
    .Y(_03952_));
 BUFx10_ASAP7_75t_R _10788_ (.A(_03952_),
    .Y(_03953_));
 BUFx6f_ASAP7_75t_R _10789_ (.A(_03953_),
    .Y(_03954_));
 BUFx12_ASAP7_75t_R _10790_ (.A(_03954_),
    .Y(_03955_));
 BUFx6f_ASAP7_75t_R _10791_ (.A(_03923_),
    .Y(_03956_));
 BUFx10_ASAP7_75t_R _10792_ (.A(_03956_),
    .Y(_03957_));
 AND2x2_ASAP7_75t_R _10793_ (.A(_03957_),
    .B(_00045_),
    .Y(_03958_));
 AO21x1_ASAP7_75t_R _10794_ (.A1(_03955_),
    .A2(_00043_),
    .B(_03958_),
    .Y(_03959_));
 AND2x6_ASAP7_75t_R _10795_ (.A(_03399_),
    .B(_03391_),
    .Y(_03960_));
 BUFx6f_ASAP7_75t_R _10796_ (.A(_03960_),
    .Y(_03961_));
 BUFx10_ASAP7_75t_R _10797_ (.A(_03961_),
    .Y(_03962_));
 AND3x4_ASAP7_75t_R _10798_ (.A(_03399_),
    .B(_03385_),
    .C(_03373_),
    .Y(_03963_));
 BUFx12f_ASAP7_75t_R _10799_ (.A(_03963_),
    .Y(_03964_));
 BUFx6f_ASAP7_75t_R _10800_ (.A(_03412_),
    .Y(_03965_));
 BUFx10_ASAP7_75t_R _10801_ (.A(_03965_),
    .Y(_03966_));
 AO21x1_ASAP7_75t_R _10802_ (.A1(_00044_),
    .A2(_03964_),
    .B(_03966_),
    .Y(_03967_));
 AO221x1_ASAP7_75t_R _10803_ (.A1(_03951_),
    .A2(_03959_),
    .B1(_03962_),
    .B2(_00046_),
    .C(_03967_),
    .Y(_03968_));
 BUFx10_ASAP7_75t_R _10804_ (.A(_03844_),
    .Y(_03969_));
 BUFx10_ASAP7_75t_R _10805_ (.A(_03969_),
    .Y(_03970_));
 BUFx10_ASAP7_75t_R _10806_ (.A(_03970_),
    .Y(_03971_));
 BUFx12f_ASAP7_75t_R _10807_ (.A(_03971_),
    .Y(_03972_));
 BUFx10_ASAP7_75t_R _10808_ (.A(_03923_),
    .Y(_03973_));
 BUFx12f_ASAP7_75t_R _10809_ (.A(_03973_),
    .Y(_03974_));
 BUFx10_ASAP7_75t_R _10810_ (.A(_03974_),
    .Y(_03975_));
 BUFx10_ASAP7_75t_R _10811_ (.A(_03949_),
    .Y(_03976_));
 BUFx10_ASAP7_75t_R _10812_ (.A(_03931_),
    .Y(_03977_));
 BUFx10_ASAP7_75t_R _10813_ (.A(_03977_),
    .Y(_03978_));
 AND2x2_ASAP7_75t_R _10814_ (.A(_03978_),
    .B(_00038_),
    .Y(_03979_));
 AO21x1_ASAP7_75t_R _10815_ (.A1(_03976_),
    .A2(_00037_),
    .B(_03979_),
    .Y(_03980_));
 BUFx10_ASAP7_75t_R _10816_ (.A(_03965_),
    .Y(_03981_));
 AO21x1_ASAP7_75t_R _10817_ (.A1(_03975_),
    .A2(_03980_),
    .B(_03981_),
    .Y(_03982_));
 BUFx12f_ASAP7_75t_R _10818_ (.A(_03482_),
    .Y(_03983_));
 BUFx6f_ASAP7_75t_R _10819_ (.A(_03983_),
    .Y(_03984_));
 BUFx10_ASAP7_75t_R _10820_ (.A(_03928_),
    .Y(_03985_));
 BUFx6f_ASAP7_75t_R _10821_ (.A(_03985_),
    .Y(_03986_));
 AND2x2_ASAP7_75t_R _10822_ (.A(_03399_),
    .B(_03373_),
    .Y(_03987_));
 BUFx12_ASAP7_75t_R _10823_ (.A(_03987_),
    .Y(_03988_));
 BUFx6f_ASAP7_75t_R _10824_ (.A(_03988_),
    .Y(_03989_));
 AO22x1_ASAP7_75t_R _10825_ (.A1(_03986_),
    .A2(_00035_),
    .B1(_00036_),
    .B2(_03989_),
    .Y(_03990_));
 BUFx12f_ASAP7_75t_R _10826_ (.A(_03953_),
    .Y(_03991_));
 BUFx10_ASAP7_75t_R _10827_ (.A(_03991_),
    .Y(_03992_));
 AO22x1_ASAP7_75t_R _10828_ (.A1(_03984_),
    .A2(_00035_),
    .B1(_03990_),
    .B2(_03992_),
    .Y(_03993_));
 AO21x1_ASAP7_75t_R _10829_ (.A1(_03972_),
    .A2(_03982_),
    .B(_03993_),
    .Y(_03994_));
 BUFx6f_ASAP7_75t_R _10830_ (.A(_03444_),
    .Y(_03995_));
 BUFx10_ASAP7_75t_R _10831_ (.A(_03995_),
    .Y(_03996_));
 BUFx10_ASAP7_75t_R _10832_ (.A(_03996_),
    .Y(_03997_));
 BUFx12_ASAP7_75t_R _10833_ (.A(_03928_),
    .Y(_03998_));
 AND2x2_ASAP7_75t_R _10834_ (.A(_03941_),
    .B(_00042_),
    .Y(_03999_));
 AO21x1_ASAP7_75t_R _10835_ (.A1(_03998_),
    .A2(_00041_),
    .B(_03999_),
    .Y(_04000_));
 BUFx10_ASAP7_75t_R _10836_ (.A(_03548_),
    .Y(_04001_));
 AND3x1_ASAP7_75t_R _10837_ (.A(_03941_),
    .B(_03378_),
    .C(_00040_),
    .Y(_04002_));
 AO21x1_ASAP7_75t_R _10838_ (.A1(_00039_),
    .A2(_04001_),
    .B(_04002_),
    .Y(_04003_));
 BUFx10_ASAP7_75t_R _10839_ (.A(_03936_),
    .Y(_04004_));
 AO221x1_ASAP7_75t_R _10840_ (.A1(_03926_),
    .A2(_04000_),
    .B1(_04003_),
    .B2(_04004_),
    .C(_03946_),
    .Y(_04005_));
 AND2x2_ASAP7_75t_R _10841_ (.A(_03997_),
    .B(_04005_),
    .Y(_04006_));
 AO32x1_ASAP7_75t_R _10842_ (.A1(_03921_),
    .A2(_03948_),
    .A3(_03968_),
    .B1(_03994_),
    .B2(_04006_),
    .Y(_04007_));
 BUFx10_ASAP7_75t_R _10843_ (.A(_03947_),
    .Y(_04008_));
 BUFx10_ASAP7_75t_R _10844_ (.A(_03413_),
    .Y(_04009_));
 AND2x2_ASAP7_75t_R _10845_ (.A(_03978_),
    .B(_00066_),
    .Y(_04010_));
 AO21x1_ASAP7_75t_R _10846_ (.A1(_03976_),
    .A2(_00065_),
    .B(_04010_),
    .Y(_04011_));
 AO221x1_ASAP7_75t_R _10847_ (.A1(_03998_),
    .A2(_00063_),
    .B1(_00064_),
    .B2(_03989_),
    .C(_03974_),
    .Y(_04012_));
 OA21x2_ASAP7_75t_R _10848_ (.A1(_03992_),
    .A2(_04011_),
    .B(_04012_),
    .Y(_04013_));
 BUFx6f_ASAP7_75t_R _10849_ (.A(_03940_),
    .Y(_04014_));
 BUFx10_ASAP7_75t_R _10850_ (.A(_04014_),
    .Y(_04015_));
 BUFx6f_ASAP7_75t_R _10851_ (.A(_04015_),
    .Y(_04016_));
 BUFx10_ASAP7_75t_R _10852_ (.A(_03924_),
    .Y(_04017_));
 BUFx10_ASAP7_75t_R _10853_ (.A(_04017_),
    .Y(_04018_));
 NOR2x2_ASAP7_75t_R _10854_ (.A(net13),
    .B(_03414_),
    .Y(_04019_));
 BUFx6f_ASAP7_75t_R _10855_ (.A(_04019_),
    .Y(_04020_));
 BUFx6f_ASAP7_75t_R _10856_ (.A(_04020_),
    .Y(_04021_));
 AO22x1_ASAP7_75t_R _10857_ (.A1(_04018_),
    .A2(_00058_),
    .B1(_04021_),
    .B2(_00056_),
    .Y(_04022_));
 BUFx10_ASAP7_75t_R _10858_ (.A(_03482_),
    .Y(_04023_));
 BUFx10_ASAP7_75t_R _10859_ (.A(_03953_),
    .Y(_04024_));
 BUFx6f_ASAP7_75t_R _10860_ (.A(_03923_),
    .Y(_04025_));
 AND2x2_ASAP7_75t_R _10861_ (.A(_04025_),
    .B(_00057_),
    .Y(_04026_));
 AO21x1_ASAP7_75t_R _10862_ (.A1(_04024_),
    .A2(_00055_),
    .B(_04026_),
    .Y(_04027_));
 BUFx10_ASAP7_75t_R _10863_ (.A(_03985_),
    .Y(_04028_));
 AO221x1_ASAP7_75t_R _10864_ (.A1(_04023_),
    .A2(_00055_),
    .B1(_04027_),
    .B2(_04028_),
    .C(_03919_),
    .Y(_04029_));
 AO21x1_ASAP7_75t_R _10865_ (.A1(_04016_),
    .A2(_04022_),
    .B(_04029_),
    .Y(_04030_));
 OA21x2_ASAP7_75t_R _10866_ (.A1(_04009_),
    .A2(_04013_),
    .B(_04030_),
    .Y(_04031_));
 BUFx10_ASAP7_75t_R _10867_ (.A(_03966_),
    .Y(_04032_));
 BUFx10_ASAP7_75t_R _10868_ (.A(_03977_),
    .Y(_04033_));
 BUFx10_ASAP7_75t_R _10869_ (.A(_04033_),
    .Y(_04034_));
 AND2x2_ASAP7_75t_R _10870_ (.A(_03973_),
    .B(_00053_),
    .Y(_04035_));
 AO21x1_ASAP7_75t_R _10871_ (.A1(_03991_),
    .A2(_00051_),
    .B(_04035_),
    .Y(_04036_));
 BUFx12_ASAP7_75t_R _10872_ (.A(_03928_),
    .Y(_04037_));
 AO221x1_ASAP7_75t_R _10873_ (.A1(_04017_),
    .A2(_00054_),
    .B1(_04021_),
    .B2(_00052_),
    .C(_04037_),
    .Y(_04038_));
 OA211x2_ASAP7_75t_R _10874_ (.A1(_04034_),
    .A2(_04036_),
    .B(_04038_),
    .C(_03996_),
    .Y(_04039_));
 BUFx6f_ASAP7_75t_R _10875_ (.A(_03953_),
    .Y(_04040_));
 AND2x2_ASAP7_75t_R _10876_ (.A(_03973_),
    .B(_00061_),
    .Y(_04041_));
 AO21x1_ASAP7_75t_R _10877_ (.A1(_04040_),
    .A2(_00059_),
    .B(_04041_),
    .Y(_04042_));
 BUFx12_ASAP7_75t_R _10878_ (.A(_03924_),
    .Y(_04043_));
 INVx1_ASAP7_75t_R _10879_ (.A(_00060_),
    .Y(_04044_));
 NAND2x1_ASAP7_75t_R _10880_ (.A(_04025_),
    .B(_00062_),
    .Y(_04045_));
 OA211x2_ASAP7_75t_R _10881_ (.A1(_04043_),
    .A2(_04044_),
    .B(_04045_),
    .C(_04014_),
    .Y(_04046_));
 INVx1_ASAP7_75t_R _10882_ (.A(_04046_),
    .Y(_04047_));
 OA211x2_ASAP7_75t_R _10883_ (.A1(_04034_),
    .A2(_04042_),
    .B(_04047_),
    .C(_03919_),
    .Y(_04048_));
 OR3x1_ASAP7_75t_R _10884_ (.A(_04032_),
    .B(_04039_),
    .C(_04048_),
    .Y(_04049_));
 AND2x6_ASAP7_75t_R _10885_ (.A(_03396_),
    .B(_03375_),
    .Y(_04050_));
 BUFx10_ASAP7_75t_R _10886_ (.A(_04050_),
    .Y(_04051_));
 OA211x2_ASAP7_75t_R _10887_ (.A1(_04008_),
    .A2(_04031_),
    .B(_04049_),
    .C(_04051_),
    .Y(_04052_));
 BUFx12f_ASAP7_75t_R _10888_ (.A(_03376_),
    .Y(_04053_));
 NAND2x2_ASAP7_75t_R _10889_ (.A(_04053_),
    .B(_03445_),
    .Y(_04054_));
 BUFx10_ASAP7_75t_R _10890_ (.A(_04054_),
    .Y(_04055_));
 AOI211x1_ASAP7_75t_R _10891_ (.A1(_03917_),
    .A2(_04007_),
    .B(_04052_),
    .C(_04055_),
    .Y(_04056_));
 AND3x1_ASAP7_75t_R _10892_ (.A(_03553_),
    .B(_03569_),
    .C(_03574_),
    .Y(_04057_));
 BUFx6f_ASAP7_75t_R _10893_ (.A(_04057_),
    .Y(_04058_));
 BUFx4f_ASAP7_75t_R _10894_ (.A(_04058_),
    .Y(_04059_));
 BUFx12_ASAP7_75t_R _10895_ (.A(_03972_),
    .Y(_04060_));
 AND4x2_ASAP7_75t_R _10896_ (.A(_03554_),
    .B(_03486_),
    .C(_03489_),
    .D(_03603_),
    .Y(_04061_));
 AO21x2_ASAP7_75t_R _10897_ (.A1(_04060_),
    .A2(net23),
    .B(_04061_),
    .Y(_04062_));
 OR2x2_ASAP7_75t_R _10898_ (.A(_04059_),
    .B(_04062_),
    .Y(_04063_));
 OA21x2_ASAP7_75t_R _10899_ (.A1(_03915_),
    .A2(_04056_),
    .B(_04063_),
    .Y(_04064_));
 XNOR2x2_ASAP7_75t_R _10900_ (.A(_03914_),
    .B(_04064_),
    .Y(_09952_));
 INVx1_ASAP7_75t_R _10901_ (.A(_09952_),
    .Y(_09954_));
 BUFx6f_ASAP7_75t_R _10902_ (.A(_04059_),
    .Y(_04065_));
 BUFx6f_ASAP7_75t_R _10903_ (.A(_04016_),
    .Y(_04066_));
 BUFx4f_ASAP7_75t_R _10904_ (.A(_03927_),
    .Y(_04067_));
 BUFx6f_ASAP7_75t_R _10905_ (.A(_04021_),
    .Y(_04068_));
 BUFx6f_ASAP7_75t_R _10906_ (.A(_04068_),
    .Y(_04069_));
 AO22x1_ASAP7_75t_R _10907_ (.A1(_04067_),
    .A2(_00090_),
    .B1(_04069_),
    .B2(_00088_),
    .Y(_04070_));
 BUFx6f_ASAP7_75t_R _10908_ (.A(_03983_),
    .Y(_04071_));
 BUFx10_ASAP7_75t_R _10909_ (.A(_04071_),
    .Y(_04072_));
 BUFx10_ASAP7_75t_R _10910_ (.A(_04024_),
    .Y(_04073_));
 BUFx10_ASAP7_75t_R _10911_ (.A(_04073_),
    .Y(_04074_));
 BUFx6f_ASAP7_75t_R _10912_ (.A(_04025_),
    .Y(_04075_));
 BUFx10_ASAP7_75t_R _10913_ (.A(_04075_),
    .Y(_04076_));
 AND2x2_ASAP7_75t_R _10914_ (.A(_04076_),
    .B(_00089_),
    .Y(_04077_));
 AO21x1_ASAP7_75t_R _10915_ (.A1(_04074_),
    .A2(_00087_),
    .B(_04077_),
    .Y(_04078_));
 BUFx6f_ASAP7_75t_R _10916_ (.A(_04028_),
    .Y(_04079_));
 BUFx6f_ASAP7_75t_R _10917_ (.A(_04079_),
    .Y(_04080_));
 AO221x1_ASAP7_75t_R _10918_ (.A1(_04072_),
    .A2(_00087_),
    .B1(_04078_),
    .B2(_04080_),
    .C(_03921_),
    .Y(_04081_));
 AO21x1_ASAP7_75t_R _10919_ (.A1(_04066_),
    .A2(_04070_),
    .B(_04081_),
    .Y(_04082_));
 BUFx6f_ASAP7_75t_R _10920_ (.A(_03964_),
    .Y(_04083_));
 BUFx10_ASAP7_75t_R _10921_ (.A(_03991_),
    .Y(_04084_));
 BUFx4f_ASAP7_75t_R _10922_ (.A(_04084_),
    .Y(_04085_));
 AND2x2_ASAP7_75t_R _10923_ (.A(_03927_),
    .B(_00097_),
    .Y(_04086_));
 AO21x1_ASAP7_75t_R _10924_ (.A1(_04085_),
    .A2(_00095_),
    .B(_04086_),
    .Y(_04087_));
 BUFx10_ASAP7_75t_R _10925_ (.A(_03976_),
    .Y(_04088_));
 BUFx12_ASAP7_75t_R _10926_ (.A(_04088_),
    .Y(_04089_));
 BUFx12_ASAP7_75t_R _10927_ (.A(_03960_),
    .Y(_04090_));
 BUFx6f_ASAP7_75t_R _10928_ (.A(_04090_),
    .Y(_04091_));
 AO21x1_ASAP7_75t_R _10929_ (.A1(_00098_),
    .A2(_04091_),
    .B(_04009_),
    .Y(_04092_));
 AO221x1_ASAP7_75t_R _10930_ (.A1(_00096_),
    .A2(_04083_),
    .B1(_04087_),
    .B2(_04089_),
    .C(_04092_),
    .Y(_04093_));
 BUFx12_ASAP7_75t_R _10931_ (.A(_03946_),
    .Y(_04094_));
 BUFx6f_ASAP7_75t_R _10932_ (.A(_04094_),
    .Y(_04095_));
 AO21x1_ASAP7_75t_R _10933_ (.A1(_04082_),
    .A2(_04093_),
    .B(_04095_),
    .Y(_04096_));
 BUFx6f_ASAP7_75t_R _10934_ (.A(_03996_),
    .Y(_04097_));
 BUFx6f_ASAP7_75t_R _10935_ (.A(_04097_),
    .Y(_04098_));
 BUFx10_ASAP7_75t_R _10936_ (.A(_04098_),
    .Y(_04099_));
 AND3x1_ASAP7_75t_R _10937_ (.A(_04066_),
    .B(_04067_),
    .C(_00094_),
    .Y(_04100_));
 BUFx6f_ASAP7_75t_R _10938_ (.A(_03988_),
    .Y(_04101_));
 BUFx12_ASAP7_75t_R _10939_ (.A(_04101_),
    .Y(_04102_));
 BUFx10_ASAP7_75t_R _10940_ (.A(_04024_),
    .Y(_04103_));
 BUFx6f_ASAP7_75t_R _10941_ (.A(_04103_),
    .Y(_04104_));
 BUFx10_ASAP7_75t_R _10942_ (.A(_04025_),
    .Y(_04105_));
 BUFx12f_ASAP7_75t_R _10943_ (.A(_04105_),
    .Y(_04106_));
 AND2x2_ASAP7_75t_R _10944_ (.A(_04106_),
    .B(_00093_),
    .Y(_04107_));
 AO21x1_ASAP7_75t_R _10945_ (.A1(_04104_),
    .A2(_00091_),
    .B(_04107_),
    .Y(_04108_));
 AO32x1_ASAP7_75t_R _10946_ (.A1(_04085_),
    .A2(_00092_),
    .A3(_04102_),
    .B1(_04108_),
    .B2(_04080_),
    .Y(_04109_));
 OR3x1_ASAP7_75t_R _10947_ (.A(_04099_),
    .B(_04100_),
    .C(_04109_),
    .Y(_04110_));
 BUFx6f_ASAP7_75t_R _10948_ (.A(_03442_),
    .Y(_04111_));
 BUFx6f_ASAP7_75t_R _10949_ (.A(_04111_),
    .Y(_04112_));
 BUFx12_ASAP7_75t_R _10950_ (.A(_04024_),
    .Y(_04113_));
 BUFx10_ASAP7_75t_R _10951_ (.A(_04113_),
    .Y(_04114_));
 AND2x2_ASAP7_75t_R _10952_ (.A(_03926_),
    .B(_00085_),
    .Y(_04115_));
 AO21x1_ASAP7_75t_R _10953_ (.A1(_04114_),
    .A2(_00083_),
    .B(_04115_),
    .Y(_04116_));
 AO32x1_ASAP7_75t_R _10954_ (.A1(_04085_),
    .A2(_00084_),
    .A3(_04102_),
    .B1(_04116_),
    .B2(_04080_),
    .Y(_04117_));
 AO221x1_ASAP7_75t_R _10955_ (.A1(_04112_),
    .A2(_03382_),
    .B1(_00086_),
    .B2(_04091_),
    .C(_04117_),
    .Y(_04118_));
 BUFx10_ASAP7_75t_R _10956_ (.A(_03981_),
    .Y(_04119_));
 BUFx6f_ASAP7_75t_R _10957_ (.A(_04119_),
    .Y(_04120_));
 AO21x1_ASAP7_75t_R _10958_ (.A1(_04110_),
    .A2(_04118_),
    .B(_04120_),
    .Y(_04121_));
 BUFx12_ASAP7_75t_R _10959_ (.A(_03916_),
    .Y(_04122_));
 AOI21x1_ASAP7_75t_R _10960_ (.A1(_04096_),
    .A2(_04121_),
    .B(_04122_),
    .Y(_04123_));
 BUFx12_ASAP7_75t_R _10961_ (.A(_04051_),
    .Y(_04124_));
 BUFx10_ASAP7_75t_R _10962_ (.A(_04037_),
    .Y(_04125_));
 BUFx6f_ASAP7_75t_R _10963_ (.A(_04125_),
    .Y(_04126_));
 BUFx6f_ASAP7_75t_R _10964_ (.A(_03933_),
    .Y(_04127_));
 AND2x2_ASAP7_75t_R _10965_ (.A(_04127_),
    .B(_00070_),
    .Y(_04128_));
 AO21x1_ASAP7_75t_R _10966_ (.A1(_04126_),
    .A2(_00069_),
    .B(_04128_),
    .Y(_04129_));
 BUFx10_ASAP7_75t_R _10967_ (.A(_03965_),
    .Y(_04130_));
 BUFx10_ASAP7_75t_R _10968_ (.A(_04130_),
    .Y(_04131_));
 AO21x1_ASAP7_75t_R _10969_ (.A1(_04067_),
    .A2(_04129_),
    .B(_04131_),
    .Y(_04132_));
 AO22x1_ASAP7_75t_R _10970_ (.A1(_03951_),
    .A2(_00067_),
    .B1(_00068_),
    .B2(_04102_),
    .Y(_04133_));
 AO22x1_ASAP7_75t_R _10971_ (.A1(_04072_),
    .A2(_00067_),
    .B1(_04133_),
    .B2(_04085_),
    .Y(_04134_));
 AO21x1_ASAP7_75t_R _10972_ (.A1(_03382_),
    .A2(_04132_),
    .B(_04134_),
    .Y(_04135_));
 BUFx6f_ASAP7_75t_R _10973_ (.A(_03930_),
    .Y(_04136_));
 BUFx10_ASAP7_75t_R _10974_ (.A(_03941_),
    .Y(_04137_));
 BUFx6f_ASAP7_75t_R _10975_ (.A(_04137_),
    .Y(_04138_));
 AND2x2_ASAP7_75t_R _10976_ (.A(_04138_),
    .B(_00074_),
    .Y(_04139_));
 AO21x1_ASAP7_75t_R _10977_ (.A1(_04136_),
    .A2(_00073_),
    .B(_04139_),
    .Y(_04140_));
 BUFx6f_ASAP7_75t_R _10978_ (.A(_03939_),
    .Y(_04141_));
 BUFx12_ASAP7_75t_R _10979_ (.A(_03943_),
    .Y(_04142_));
 AND3x1_ASAP7_75t_R _10980_ (.A(_04016_),
    .B(_04142_),
    .C(_00072_),
    .Y(_04143_));
 AO21x1_ASAP7_75t_R _10981_ (.A1(_00071_),
    .A2(_04141_),
    .B(_04143_),
    .Y(_04144_));
 BUFx4f_ASAP7_75t_R _10982_ (.A(_03938_),
    .Y(_04145_));
 AO221x1_ASAP7_75t_R _10983_ (.A1(_04067_),
    .A2(_04140_),
    .B1(_04144_),
    .B2(_04145_),
    .C(_04095_),
    .Y(_04146_));
 AND2x2_ASAP7_75t_R _10984_ (.A(_04138_),
    .B(_00082_),
    .Y(_04147_));
 AO21x1_ASAP7_75t_R _10985_ (.A1(_04136_),
    .A2(_00081_),
    .B(_04147_),
    .Y(_04148_));
 AND3x1_ASAP7_75t_R _10986_ (.A(_04016_),
    .B(_04142_),
    .C(_00080_),
    .Y(_04149_));
 AO21x1_ASAP7_75t_R _10987_ (.A1(_00079_),
    .A2(_04141_),
    .B(_04149_),
    .Y(_04150_));
 AO221x1_ASAP7_75t_R _10988_ (.A1(_04067_),
    .A2(_04148_),
    .B1(_04150_),
    .B2(_04145_),
    .C(_04095_),
    .Y(_04151_));
 AND2x2_ASAP7_75t_R _10989_ (.A(_03926_),
    .B(_00077_),
    .Y(_04152_));
 AO21x1_ASAP7_75t_R _10990_ (.A1(_04114_),
    .A2(_00075_),
    .B(_04152_),
    .Y(_04153_));
 AO22x1_ASAP7_75t_R _10991_ (.A1(_00078_),
    .A2(_04091_),
    .B1(_04153_),
    .B2(_04136_),
    .Y(_04154_));
 AO21x1_ASAP7_75t_R _10992_ (.A1(_00076_),
    .A2(_04083_),
    .B(_04119_),
    .Y(_04155_));
 BUFx10_ASAP7_75t_R _10993_ (.A(_03919_),
    .Y(_04156_));
 BUFx10_ASAP7_75t_R _10994_ (.A(_04156_),
    .Y(_04157_));
 OA21x2_ASAP7_75t_R _10995_ (.A1(_04154_),
    .A2(_04155_),
    .B(_04157_),
    .Y(_04158_));
 AO32x1_ASAP7_75t_R _10996_ (.A1(_04099_),
    .A2(_04135_),
    .A3(_04146_),
    .B1(_04151_),
    .B2(_04158_),
    .Y(_04159_));
 NOR2x1_ASAP7_75t_R _10997_ (.A(_04124_),
    .B(_04159_),
    .Y(_04160_));
 OA21x2_ASAP7_75t_R _10998_ (.A1(_04123_),
    .A2(_04160_),
    .B(_03447_),
    .Y(_04161_));
 BUFx4f_ASAP7_75t_R _10999_ (.A(_03915_),
    .Y(_04162_));
 BUFx12f_ASAP7_75t_R _11000_ (.A(_03539_),
    .Y(_04163_));
 BUFx12f_ASAP7_75t_R _11001_ (.A(_04163_),
    .Y(_04164_));
 BUFx12f_ASAP7_75t_R _11002_ (.A(_04164_),
    .Y(_04165_));
 INVx1_ASAP7_75t_R _11003_ (.A(_03547_),
    .Y(_04166_));
 BUFx12_ASAP7_75t_R _11004_ (.A(_04166_),
    .Y(net64));
 OR4x2_ASAP7_75t_R _11005_ (.A(_04165_),
    .B(_03542_),
    .C(net64),
    .D(_04062_),
    .Y(_04167_));
 BUFx4f_ASAP7_75t_R _11006_ (.A(_04167_),
    .Y(_04168_));
 AND2x6_ASAP7_75t_R _11007_ (.A(_04142_),
    .B(net22),
    .Y(_04169_));
 AND3x1_ASAP7_75t_R _11008_ (.A(_03497_),
    .B(_03502_),
    .C(_03557_),
    .Y(_04170_));
 BUFx4f_ASAP7_75t_R _11009_ (.A(_04170_),
    .Y(_04171_));
 BUFx3_ASAP7_75t_R _11010_ (.A(_03540_),
    .Y(_04172_));
 AND2x2_ASAP7_75t_R _11011_ (.A(_04171_),
    .B(_04172_),
    .Y(_04173_));
 NAND2x2_ASAP7_75t_R _11012_ (.A(_04171_),
    .B(_03541_),
    .Y(_04174_));
 AO32x1_ASAP7_75t_R _11013_ (.A1(_03822_),
    .A2(_04174_),
    .A3(_03547_),
    .B1(_04062_),
    .B2(_03503_),
    .Y(_04175_));
 AO21x1_ASAP7_75t_R _11014_ (.A1(_04062_),
    .A2(_04173_),
    .B(_04175_),
    .Y(_04176_));
 AO21x1_ASAP7_75t_R _11015_ (.A1(_03600_),
    .A2(_04169_),
    .B(_04176_),
    .Y(_04177_));
 AND2x2_ASAP7_75t_R _11016_ (.A(_04168_),
    .B(_04177_),
    .Y(_10168_));
 AND2x2_ASAP7_75t_R _11017_ (.A(_04162_),
    .B(_10168_),
    .Y(_04178_));
 AO21x1_ASAP7_75t_R _11018_ (.A1(_04065_),
    .A2(_04161_),
    .B(_04178_),
    .Y(_04179_));
 XNOR2x2_ASAP7_75t_R _11019_ (.A(_03914_),
    .B(_04179_),
    .Y(_09960_));
 INVx1_ASAP7_75t_R _11020_ (.A(_09960_),
    .Y(_09958_));
 OA211x2_ASAP7_75t_R _11021_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03727_),
    .C(_00072_),
    .Y(_04180_));
 AO21x1_ASAP7_75t_R _11022_ (.A1(_00071_),
    .A2(_03584_),
    .B(_04180_),
    .Y(_04181_));
 OA222x2_ASAP7_75t_R _11023_ (.A1(_00073_),
    .A2(_03885_),
    .B1(_03584_),
    .B2(_00074_),
    .C1(_03680_),
    .C2(_03605_),
    .Y(_04182_));
 AO21x1_ASAP7_75t_R _11024_ (.A1(_03824_),
    .A2(_04181_),
    .B(_04182_),
    .Y(_04183_));
 INVx1_ASAP7_75t_R _11025_ (.A(_00069_),
    .Y(_04184_));
 AND2x6_ASAP7_75t_R _11026_ (.A(_03618_),
    .B(_03591_),
    .Y(_04185_));
 INVx1_ASAP7_75t_R _11027_ (.A(_00068_),
    .Y(_04186_));
 NAND2x1_ASAP7_75t_R _11028_ (.A(_03591_),
    .B(_00070_),
    .Y(_04187_));
 OA211x2_ASAP7_75t_R _11029_ (.A1(_03619_),
    .A2(_04186_),
    .B(_04187_),
    .C(_03613_),
    .Y(_04188_));
 AOI21x1_ASAP7_75t_R _11030_ (.A1(_04184_),
    .A2(_04185_),
    .B(_04188_),
    .Y(_04189_));
 OA211x2_ASAP7_75t_R _11031_ (.A1(_03628_),
    .A2(_04189_),
    .B(_03771_),
    .C(_03827_),
    .Y(_04190_));
 OA22x2_ASAP7_75t_R _11032_ (.A1(_00067_),
    .A2(_03758_),
    .B1(_04190_),
    .B2(_03539_),
    .Y(_04191_));
 AND2x2_ASAP7_75t_R _11033_ (.A(_03594_),
    .B(_03597_),
    .Y(_04192_));
 AND2x2_ASAP7_75t_R _11034_ (.A(_03590_),
    .B(_04192_),
    .Y(_04193_));
 OR3x4_ASAP7_75t_R _11035_ (.A(_03599_),
    .B(_04061_),
    .C(_03906_),
    .Y(_04194_));
 AO21x2_ASAP7_75t_R _11036_ (.A1(_03648_),
    .A2(_04193_),
    .B(_04194_),
    .Y(_04195_));
 AO211x2_ASAP7_75t_R _11037_ (.A1(_03790_),
    .A2(_04183_),
    .B(_04191_),
    .C(_04195_),
    .Y(_04196_));
 OA21x2_ASAP7_75t_R _11038_ (.A1(_03756_),
    .A2(_03668_),
    .B(_03726_),
    .Y(_04197_));
 BUFx12f_ASAP7_75t_R _11039_ (.A(_04197_),
    .Y(_04198_));
 OA21x2_ASAP7_75t_R _11040_ (.A1(_03756_),
    .A2(_03668_),
    .B(_03709_),
    .Y(_04199_));
 AND3x1_ASAP7_75t_R _11041_ (.A(_00077_),
    .B(_03827_),
    .C(_03691_),
    .Y(_04200_));
 AO221x1_ASAP7_75t_R _11042_ (.A1(_00082_),
    .A2(_04198_),
    .B1(_04199_),
    .B2(_00081_),
    .C(_04200_),
    .Y(_04201_));
 AO21x1_ASAP7_75t_R _11043_ (.A1(_00078_),
    .A2(_03833_),
    .B(_03824_),
    .Y(_04202_));
 INVx1_ASAP7_75t_R _11044_ (.A(_00075_),
    .Y(_04203_));
 AND2x4_ASAP7_75t_R _11045_ (.A(_03393_),
    .B(_03690_),
    .Y(_04204_));
 OA211x2_ASAP7_75t_R _11046_ (.A1(_03756_),
    .A2(_04204_),
    .B(_03509_),
    .C(_03556_),
    .Y(_04205_));
 BUFx4f_ASAP7_75t_R _11047_ (.A(_04205_),
    .Y(_04206_));
 AND2x2_ASAP7_75t_R _11048_ (.A(_03608_),
    .B(_00080_),
    .Y(_04207_));
 AO21x1_ASAP7_75t_R _11049_ (.A1(_03683_),
    .A2(_00076_),
    .B(_04207_),
    .Y(_04208_));
 AND2x2_ASAP7_75t_R _11050_ (.A(_03618_),
    .B(net8),
    .Y(_04209_));
 BUFx12f_ASAP7_75t_R _11051_ (.A(_04209_),
    .Y(_04210_));
 AOI22x1_ASAP7_75t_R _11052_ (.A1(_03716_),
    .A2(_04208_),
    .B1(_04210_),
    .B2(_00079_),
    .Y(_04211_));
 BUFx6f_ASAP7_75t_R _11053_ (.A(_03592_),
    .Y(_04212_));
 OA211x2_ASAP7_75t_R _11054_ (.A1(_03628_),
    .A2(_04211_),
    .B(_04212_),
    .C(_03827_),
    .Y(_04213_));
 BUFx12f_ASAP7_75t_R _11055_ (.A(_03539_),
    .Y(_04214_));
 OAI22x1_ASAP7_75t_R _11056_ (.A1(_04203_),
    .A2(_04206_),
    .B1(_04213_),
    .B2(_04214_),
    .Y(_04215_));
 OA211x2_ASAP7_75t_R _11057_ (.A1(_04201_),
    .A2(_04202_),
    .B(_03697_),
    .C(_04215_),
    .Y(_04216_));
 INVx1_ASAP7_75t_R _11058_ (.A(_00091_),
    .Y(_04217_));
 BUFx12_ASAP7_75t_R _11059_ (.A(_04206_),
    .Y(_04218_));
 AND2x2_ASAP7_75t_R _11060_ (.A(_03608_),
    .B(_00096_),
    .Y(_04219_));
 AO21x1_ASAP7_75t_R _11061_ (.A1(_03683_),
    .A2(_00092_),
    .B(_04219_),
    .Y(_04220_));
 AOI22x1_ASAP7_75t_R _11062_ (.A1(_00095_),
    .A2(_04210_),
    .B1(_04220_),
    .B2(_03664_),
    .Y(_04221_));
 OA211x2_ASAP7_75t_R _11063_ (.A1(_03419_),
    .A2(_04221_),
    .B(_04212_),
    .C(_03736_),
    .Y(_04222_));
 OAI22x1_ASAP7_75t_R _11064_ (.A1(_04217_),
    .A2(_04218_),
    .B1(_04222_),
    .B2(_04214_),
    .Y(_04223_));
 AND3x1_ASAP7_75t_R _11065_ (.A(_03394_),
    .B(_03613_),
    .C(_00094_),
    .Y(_04224_));
 AO21x1_ASAP7_75t_R _11066_ (.A1(_00093_),
    .A2(_03709_),
    .B(_04224_),
    .Y(_04225_));
 OR3x1_ASAP7_75t_R _11067_ (.A(_03605_),
    .B(_03669_),
    .C(_04225_),
    .Y(_04226_));
 AND2x2_ASAP7_75t_R _11068_ (.A(_00097_),
    .B(_03582_),
    .Y(_04227_));
 AO221x1_ASAP7_75t_R _11069_ (.A1(_00098_),
    .A2(_03727_),
    .B1(_03734_),
    .B2(_03827_),
    .C(_04227_),
    .Y(_04228_));
 AO21x1_ASAP7_75t_R _11070_ (.A1(_03736_),
    .A2(_04212_),
    .B(_03722_),
    .Y(_04229_));
 AO21x1_ASAP7_75t_R _11071_ (.A1(_04226_),
    .A2(_04228_),
    .B(_04229_),
    .Y(_04230_));
 OR2x2_ASAP7_75t_R _11072_ (.A(_03697_),
    .B(_03722_),
    .Y(_04231_));
 OA211x2_ASAP7_75t_R _11073_ (.A1(_03722_),
    .A2(_04223_),
    .B(_04230_),
    .C(_04231_),
    .Y(_04232_));
 BUFx6f_ASAP7_75t_R _11074_ (.A(_03604_),
    .Y(_04233_));
 OR3x1_ASAP7_75t_R _11075_ (.A(_00084_),
    .B(_04233_),
    .C(_03680_),
    .Y(_04234_));
 AO21x1_ASAP7_75t_R _11076_ (.A1(_03660_),
    .A2(_03801_),
    .B(_00086_),
    .Y(_04235_));
 BUFx12_ASAP7_75t_R _11077_ (.A(_03671_),
    .Y(_04236_));
 AO21x1_ASAP7_75t_R _11078_ (.A1(_04234_),
    .A2(_04235_),
    .B(_04236_),
    .Y(_04237_));
 OR2x2_ASAP7_75t_R _11079_ (.A(_00085_),
    .B(_03864_),
    .Y(_04238_));
 OA21x2_ASAP7_75t_R _11080_ (.A1(_00083_),
    .A2(_03758_),
    .B(_03700_),
    .Y(_04239_));
 OR3x1_ASAP7_75t_R _11081_ (.A(_00088_),
    .B(_04233_),
    .C(_03680_),
    .Y(_04240_));
 AO21x1_ASAP7_75t_R _11082_ (.A1(_03660_),
    .A2(_03801_),
    .B(_00090_),
    .Y(_04241_));
 BUFx16f_ASAP7_75t_R _11083_ (.A(_03671_),
    .Y(_04242_));
 AO21x1_ASAP7_75t_R _11084_ (.A1(_04240_),
    .A2(_04241_),
    .B(_04242_),
    .Y(_04243_));
 BUFx6f_ASAP7_75t_R _11085_ (.A(_03517_),
    .Y(_04244_));
 OR3x1_ASAP7_75t_R _11086_ (.A(_00087_),
    .B(_03605_),
    .C(_03757_),
    .Y(_04245_));
 AO221x1_ASAP7_75t_R _11087_ (.A1(_03395_),
    .A2(_03716_),
    .B1(_03645_),
    .B2(_03593_),
    .C(_00089_),
    .Y(_04246_));
 AND4x1_ASAP7_75t_R _11088_ (.A(_04244_),
    .B(_03652_),
    .C(_04245_),
    .D(_04246_),
    .Y(_04247_));
 AO32x1_ASAP7_75t_R _11089_ (.A1(_04237_),
    .A2(_04238_),
    .A3(_04239_),
    .B1(_04243_),
    .B2(_04247_),
    .Y(_04248_));
 OA22x2_ASAP7_75t_R _11090_ (.A1(_04196_),
    .A2(_04216_),
    .B1(_04232_),
    .B2(_04248_),
    .Y(_04249_));
 BUFx6f_ASAP7_75t_R _11091_ (.A(_04249_),
    .Y(_09957_));
 INVx5_ASAP7_75t_R _11092_ (.A(_09957_),
    .Y(_09959_));
 BUFx6f_ASAP7_75t_R _11093_ (.A(_04162_),
    .Y(_04250_));
 BUFx3_ASAP7_75t_R _11094_ (.A(_04176_),
    .Y(_04251_));
 AND3x1_ASAP7_75t_R _11095_ (.A(net89),
    .B(net20),
    .C(_03600_),
    .Y(_04252_));
 BUFx3_ASAP7_75t_R _11096_ (.A(_04168_),
    .Y(_04253_));
 OA21x2_ASAP7_75t_R _11097_ (.A1(_04251_),
    .A2(_04252_),
    .B(_04253_),
    .Y(_10166_));
 BUFx6f_ASAP7_75t_R _11098_ (.A(_03915_),
    .Y(_04254_));
 BUFx10_ASAP7_75t_R _11099_ (.A(_04018_),
    .Y(_04255_));
 BUFx6f_ASAP7_75t_R _11100_ (.A(_03932_),
    .Y(_04256_));
 AND2x2_ASAP7_75t_R _11101_ (.A(_04256_),
    .B(_00116_),
    .Y(_04257_));
 AO21x1_ASAP7_75t_R _11102_ (.A1(_04125_),
    .A2(_00115_),
    .B(_04257_),
    .Y(_04258_));
 AND3x1_ASAP7_75t_R _11103_ (.A(_03933_),
    .B(_03379_),
    .C(_00114_),
    .Y(_04259_));
 AO21x1_ASAP7_75t_R _11104_ (.A1(_00113_),
    .A2(_03939_),
    .B(_04259_),
    .Y(_04260_));
 AO221x1_ASAP7_75t_R _11105_ (.A1(_04255_),
    .A2(_04258_),
    .B1(_04260_),
    .B2(_03938_),
    .C(_03947_),
    .Y(_04261_));
 BUFx10_ASAP7_75t_R _11106_ (.A(_03960_),
    .Y(_04262_));
 AND2x2_ASAP7_75t_R _11107_ (.A(_03957_),
    .B(_00111_),
    .Y(_04263_));
 AO21x1_ASAP7_75t_R _11108_ (.A1(_03955_),
    .A2(_00109_),
    .B(_04263_),
    .Y(_04264_));
 BUFx6f_ASAP7_75t_R _11109_ (.A(_03976_),
    .Y(_04265_));
 BUFx12_ASAP7_75t_R _11110_ (.A(_03963_),
    .Y(_04266_));
 AO21x1_ASAP7_75t_R _11111_ (.A1(_00110_),
    .A2(_04266_),
    .B(_03966_),
    .Y(_04267_));
 AO221x1_ASAP7_75t_R _11112_ (.A1(_00112_),
    .A2(_04262_),
    .B1(_04264_),
    .B2(_04265_),
    .C(_04267_),
    .Y(_04268_));
 BUFx6f_ASAP7_75t_R _11113_ (.A(_03956_),
    .Y(_04269_));
 BUFx6f_ASAP7_75t_R _11114_ (.A(_04269_),
    .Y(_04270_));
 AND2x2_ASAP7_75t_R _11115_ (.A(_03978_),
    .B(_00104_),
    .Y(_04271_));
 AO21x1_ASAP7_75t_R _11116_ (.A1(_03976_),
    .A2(_00103_),
    .B(_04271_),
    .Y(_04272_));
 AO21x1_ASAP7_75t_R _11117_ (.A1(_04270_),
    .A2(_04272_),
    .B(_03981_),
    .Y(_04273_));
 BUFx10_ASAP7_75t_R _11118_ (.A(_03985_),
    .Y(_04274_));
 AO22x1_ASAP7_75t_R _11119_ (.A1(_04274_),
    .A2(_00101_),
    .B1(_00102_),
    .B2(_03989_),
    .Y(_04275_));
 BUFx10_ASAP7_75t_R _11120_ (.A(_03954_),
    .Y(_04276_));
 AO22x1_ASAP7_75t_R _11121_ (.A1(_03984_),
    .A2(_00101_),
    .B1(_04275_),
    .B2(_04276_),
    .Y(_04277_));
 AO21x1_ASAP7_75t_R _11122_ (.A1(_03972_),
    .A2(_04273_),
    .B(_04277_),
    .Y(_04278_));
 BUFx10_ASAP7_75t_R _11123_ (.A(_03919_),
    .Y(_04279_));
 BUFx12_ASAP7_75t_R _11124_ (.A(_04279_),
    .Y(_04280_));
 BUFx10_ASAP7_75t_R _11125_ (.A(_03949_),
    .Y(_04281_));
 AND2x2_ASAP7_75t_R _11126_ (.A(_04256_),
    .B(_00108_),
    .Y(_04282_));
 AO21x1_ASAP7_75t_R _11127_ (.A1(_04281_),
    .A2(_00107_),
    .B(_04282_),
    .Y(_04283_));
 AND3x1_ASAP7_75t_R _11128_ (.A(_04256_),
    .B(_03379_),
    .C(_00106_),
    .Y(_04284_));
 AO21x1_ASAP7_75t_R _11129_ (.A1(_00105_),
    .A2(_03939_),
    .B(_04284_),
    .Y(_04285_));
 AOI221x1_ASAP7_75t_R _11130_ (.A1(_04255_),
    .A2(_04283_),
    .B1(_04285_),
    .B2(_03938_),
    .C(_03947_),
    .Y(_04286_));
 NOR2x1_ASAP7_75t_R _11131_ (.A(_04280_),
    .B(_04286_),
    .Y(_04287_));
 AO32x1_ASAP7_75t_R _11132_ (.A1(_03921_),
    .A2(_04261_),
    .A3(_04268_),
    .B1(_04278_),
    .B2(_04287_),
    .Y(_04288_));
 BUFx6f_ASAP7_75t_R _11133_ (.A(_04106_),
    .Y(_04289_));
 AND2x2_ASAP7_75t_R _11134_ (.A(_04137_),
    .B(_00124_),
    .Y(_04290_));
 AO21x1_ASAP7_75t_R _11135_ (.A1(_03930_),
    .A2(_00123_),
    .B(_04290_),
    .Y(_04291_));
 BUFx10_ASAP7_75t_R _11136_ (.A(_04001_),
    .Y(_04292_));
 AND3x1_ASAP7_75t_R _11137_ (.A(_03942_),
    .B(_03943_),
    .C(_00122_),
    .Y(_04293_));
 AO21x1_ASAP7_75t_R _11138_ (.A1(_00121_),
    .A2(_04292_),
    .B(_04293_),
    .Y(_04294_));
 BUFx6f_ASAP7_75t_R _11139_ (.A(_04004_),
    .Y(_04295_));
 BUFx10_ASAP7_75t_R _11140_ (.A(_03418_),
    .Y(_04296_));
 OR3x2_ASAP7_75t_R _11141_ (.A(_04296_),
    .B(_04111_),
    .C(_03482_),
    .Y(_04297_));
 BUFx6f_ASAP7_75t_R _11142_ (.A(_04297_),
    .Y(_04298_));
 AO221x1_ASAP7_75t_R _11143_ (.A1(_04289_),
    .A2(_04291_),
    .B1(_04294_),
    .B2(_04295_),
    .C(_04298_),
    .Y(_04299_));
 AND2x2_ASAP7_75t_R _11144_ (.A(_04137_),
    .B(_00132_),
    .Y(_04300_));
 AO21x1_ASAP7_75t_R _11145_ (.A1(_03930_),
    .A2(_00131_),
    .B(_04300_),
    .Y(_04301_));
 AND3x1_ASAP7_75t_R _11146_ (.A(_03942_),
    .B(_03943_),
    .C(_00130_),
    .Y(_04302_));
 AO21x1_ASAP7_75t_R _11147_ (.A1(_00129_),
    .A2(_04292_),
    .B(_04302_),
    .Y(_04303_));
 BUFx6f_ASAP7_75t_R _11148_ (.A(_03420_),
    .Y(_04304_));
 AO221x1_ASAP7_75t_R _11149_ (.A1(_03927_),
    .A2(_04301_),
    .B1(_04303_),
    .B2(_03938_),
    .C(_04304_),
    .Y(_04305_));
 AND3x1_ASAP7_75t_R _11150_ (.A(_04051_),
    .B(_04299_),
    .C(_04305_),
    .Y(_04306_));
 BUFx12f_ASAP7_75t_R _11151_ (.A(_03978_),
    .Y(_04307_));
 BUFx10_ASAP7_75t_R _11152_ (.A(_04307_),
    .Y(_04308_));
 AO221x1_ASAP7_75t_R _11153_ (.A1(_04106_),
    .A2(_00128_),
    .B1(_04068_),
    .B2(_00126_),
    .C(_04097_),
    .Y(_04309_));
 AO221x1_ASAP7_75t_R _11154_ (.A1(_04106_),
    .A2(_00120_),
    .B1(_04068_),
    .B2(_00118_),
    .C(_04279_),
    .Y(_04310_));
 AND3x1_ASAP7_75t_R _11155_ (.A(_04308_),
    .B(_04309_),
    .C(_04310_),
    .Y(_04311_));
 AND2x2_ASAP7_75t_R _11156_ (.A(_04269_),
    .B(_00127_),
    .Y(_04312_));
 AO21x1_ASAP7_75t_R _11157_ (.A1(_04276_),
    .A2(_00125_),
    .B(_04312_),
    .Y(_04313_));
 BUFx6f_ASAP7_75t_R _11158_ (.A(_03969_),
    .Y(_04314_));
 BUFx12f_ASAP7_75t_R _11159_ (.A(_04314_),
    .Y(_04315_));
 AND2x2_ASAP7_75t_R _11160_ (.A(_04105_),
    .B(_00119_),
    .Y(_04316_));
 AO221x1_ASAP7_75t_R _11161_ (.A1(_04111_),
    .A2(_04315_),
    .B1(_00117_),
    .B2(_04103_),
    .C(_04316_),
    .Y(_04317_));
 OA211x2_ASAP7_75t_R _11162_ (.A1(_03997_),
    .A2(_04313_),
    .B(_04317_),
    .C(_04265_),
    .Y(_04318_));
 OR3x1_ASAP7_75t_R _11163_ (.A(_04131_),
    .B(_04311_),
    .C(_04318_),
    .Y(_04319_));
 AO221x2_ASAP7_75t_R _11164_ (.A1(_03917_),
    .A2(_04288_),
    .B1(_04306_),
    .B2(_04319_),
    .C(_04055_),
    .Y(_04320_));
 NOR2x1_ASAP7_75t_R _11165_ (.A(_04254_),
    .B(_04320_),
    .Y(_04321_));
 AOI21x1_ASAP7_75t_R _11166_ (.A1(_04250_),
    .A2(_10166_),
    .B(_04321_),
    .Y(_04322_));
 XNOR2x1_ASAP7_75t_R _11167_ (.B(_04322_),
    .Y(_09965_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _11168_ (.A(_09965_),
    .Y(_09963_));
 INVx1_ASAP7_75t_R _11169_ (.A(_00125_),
    .Y(_04323_));
 AND2x2_ASAP7_75t_R _11170_ (.A(_03685_),
    .B(_00130_),
    .Y(_04324_));
 AO21x1_ASAP7_75t_R _11171_ (.A1(_03683_),
    .A2(_00126_),
    .B(_04324_),
    .Y(_04325_));
 AOI22x1_ASAP7_75t_R _11172_ (.A1(_00129_),
    .A2(_04210_),
    .B1(_04325_),
    .B2(_03664_),
    .Y(_04326_));
 OA211x2_ASAP7_75t_R _11173_ (.A1(_03419_),
    .A2(_04326_),
    .B(_04212_),
    .C(_03736_),
    .Y(_04327_));
 OAI22x1_ASAP7_75t_R _11174_ (.A1(_04323_),
    .A2(_04218_),
    .B1(_04327_),
    .B2(_04214_),
    .Y(_04328_));
 AND3x1_ASAP7_75t_R _11175_ (.A(_03374_),
    .B(_03614_),
    .C(_00128_),
    .Y(_04329_));
 AND2x2_ASAP7_75t_R _11176_ (.A(_00127_),
    .B(_03582_),
    .Y(_04330_));
 OR4x1_ASAP7_75t_R _11177_ (.A(_03605_),
    .B(_03669_),
    .C(_04329_),
    .D(_04330_),
    .Y(_04331_));
 AND2x2_ASAP7_75t_R _11178_ (.A(_00131_),
    .B(_03582_),
    .Y(_04332_));
 AO221x1_ASAP7_75t_R _11179_ (.A1(_00132_),
    .A2(_03727_),
    .B1(_03734_),
    .B2(_03827_),
    .C(_04332_),
    .Y(_04333_));
 AO21x1_ASAP7_75t_R _11180_ (.A1(_04331_),
    .A2(_04333_),
    .B(_04229_),
    .Y(_04334_));
 OA211x2_ASAP7_75t_R _11181_ (.A1(_03723_),
    .A2(_04328_),
    .B(_04334_),
    .C(_04231_),
    .Y(_04335_));
 OR3x1_ASAP7_75t_R _11182_ (.A(_00118_),
    .B(_04233_),
    .C(_03680_),
    .Y(_04336_));
 AO21x1_ASAP7_75t_R _11183_ (.A1(_03660_),
    .A2(_03801_),
    .B(_00120_),
    .Y(_04337_));
 AO21x1_ASAP7_75t_R _11184_ (.A1(_04336_),
    .A2(_04337_),
    .B(_04236_),
    .Y(_04338_));
 OR2x2_ASAP7_75t_R _11185_ (.A(_00119_),
    .B(_03865_),
    .Y(_04339_));
 OA21x2_ASAP7_75t_R _11186_ (.A1(_00117_),
    .A2(_03758_),
    .B(_03700_),
    .Y(_04340_));
 OR3x1_ASAP7_75t_R _11187_ (.A(_00122_),
    .B(_04233_),
    .C(_03680_),
    .Y(_04341_));
 AO21x1_ASAP7_75t_R _11188_ (.A1(_03660_),
    .A2(_03801_),
    .B(_00124_),
    .Y(_04342_));
 AO21x1_ASAP7_75t_R _11189_ (.A1(_04341_),
    .A2(_04342_),
    .B(_04236_),
    .Y(_04343_));
 BUFx12_ASAP7_75t_R _11190_ (.A(_03757_),
    .Y(_04344_));
 OR3x1_ASAP7_75t_R _11191_ (.A(_00121_),
    .B(_03605_),
    .C(_04344_),
    .Y(_04345_));
 AO221x1_ASAP7_75t_R _11192_ (.A1(_03443_),
    .A2(_03716_),
    .B1(_03645_),
    .B2(_03593_),
    .C(_00123_),
    .Y(_04346_));
 AND4x1_ASAP7_75t_R _11193_ (.A(_04244_),
    .B(_03652_),
    .C(_04345_),
    .D(_04346_),
    .Y(_04347_));
 AO32x1_ASAP7_75t_R _11194_ (.A1(_04338_),
    .A2(_04339_),
    .A3(_04340_),
    .B1(_04343_),
    .B2(_04347_),
    .Y(_04348_));
 OR3x1_ASAP7_75t_R _11195_ (.A(_00112_),
    .B(_04233_),
    .C(_03669_),
    .Y(_04349_));
 BUFx10_ASAP7_75t_R _11196_ (.A(_03645_),
    .Y(_04350_));
 AO21x1_ASAP7_75t_R _11197_ (.A1(_04350_),
    .A2(_03734_),
    .B(_00116_),
    .Y(_04351_));
 AO21x1_ASAP7_75t_R _11198_ (.A1(_04349_),
    .A2(_04351_),
    .B(_03869_),
    .Y(_04352_));
 INVx1_ASAP7_75t_R _11199_ (.A(_00109_),
    .Y(_04353_));
 AND2x2_ASAP7_75t_R _11200_ (.A(_03608_),
    .B(_00114_),
    .Y(_04354_));
 AO21x1_ASAP7_75t_R _11201_ (.A1(_03683_),
    .A2(_00110_),
    .B(_04354_),
    .Y(_04355_));
 AOI22x1_ASAP7_75t_R _11202_ (.A1(_00113_),
    .A2(_04210_),
    .B1(_04355_),
    .B2(_03716_),
    .Y(_04356_));
 OA211x2_ASAP7_75t_R _11203_ (.A1(_03419_),
    .A2(_04356_),
    .B(_04212_),
    .C(_03736_),
    .Y(_04357_));
 OAI22x1_ASAP7_75t_R _11204_ (.A1(_04353_),
    .A2(_04218_),
    .B1(_04357_),
    .B2(_04214_),
    .Y(_04358_));
 OR3x1_ASAP7_75t_R _11205_ (.A(_00111_),
    .B(_03605_),
    .C(_03669_),
    .Y(_04359_));
 AO21x1_ASAP7_75t_R _11206_ (.A1(_04350_),
    .A2(_03734_),
    .B(_00115_),
    .Y(_04360_));
 AO21x1_ASAP7_75t_R _11207_ (.A1(_04359_),
    .A2(_04360_),
    .B(_03865_),
    .Y(_04361_));
 AND4x1_ASAP7_75t_R _11208_ (.A(_03697_),
    .B(_04352_),
    .C(_04358_),
    .D(_04361_),
    .Y(_04362_));
 OA211x2_ASAP7_75t_R _11209_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03727_),
    .C(_00106_),
    .Y(_04363_));
 AO21x1_ASAP7_75t_R _11210_ (.A1(_00105_),
    .A2(_03584_),
    .B(_04363_),
    .Y(_04364_));
 OA222x2_ASAP7_75t_R _11211_ (.A1(_00107_),
    .A2(_03885_),
    .B1(_03584_),
    .B2(_00108_),
    .C1(_03680_),
    .C2(_03605_),
    .Y(_04365_));
 AO21x1_ASAP7_75t_R _11212_ (.A1(_03824_),
    .A2(_04364_),
    .B(_04365_),
    .Y(_04366_));
 INVx1_ASAP7_75t_R _11213_ (.A(_00103_),
    .Y(_04367_));
 INVx2_ASAP7_75t_R _11214_ (.A(_00102_),
    .Y(_04368_));
 NAND2x1_ASAP7_75t_R _11215_ (.A(_03591_),
    .B(_00104_),
    .Y(_04369_));
 OA211x2_ASAP7_75t_R _11216_ (.A1(_03619_),
    .A2(_04368_),
    .B(_04369_),
    .C(_03613_),
    .Y(_04370_));
 AOI21x1_ASAP7_75t_R _11217_ (.A1(_04367_),
    .A2(_04185_),
    .B(_04370_),
    .Y(_04371_));
 OA211x2_ASAP7_75t_R _11218_ (.A1(_03628_),
    .A2(_04371_),
    .B(_03771_),
    .C(_03827_),
    .Y(_04372_));
 OA22x2_ASAP7_75t_R _11219_ (.A1(_00101_),
    .A2(_03759_),
    .B1(_04372_),
    .B2(_04214_),
    .Y(_04373_));
 AO211x2_ASAP7_75t_R _11220_ (.A1(_03791_),
    .A2(_04366_),
    .B(_04373_),
    .C(_04195_),
    .Y(_04374_));
 OA22x2_ASAP7_75t_R _11221_ (.A1(_04335_),
    .A2(_04348_),
    .B1(_04362_),
    .B2(_04374_),
    .Y(_04375_));
 BUFx6f_ASAP7_75t_R _11222_ (.A(_04375_),
    .Y(_09962_));
 INVx4_ASAP7_75t_R _11223_ (.A(_09962_),
    .Y(_09964_));
 AND3x1_ASAP7_75t_R _11224_ (.A(net89),
    .B(net19),
    .C(_03600_),
    .Y(_04376_));
 OA21x2_ASAP7_75t_R _11225_ (.A1(_04251_),
    .A2(_04376_),
    .B(_04253_),
    .Y(_10164_));
 AND2x2_ASAP7_75t_R _11226_ (.A(_04014_),
    .B(_00166_),
    .Y(_04377_));
 AO21x1_ASAP7_75t_R _11227_ (.A1(_04274_),
    .A2(_00165_),
    .B(_04377_),
    .Y(_04378_));
 AND3x1_ASAP7_75t_R _11228_ (.A(_04014_),
    .B(_03970_),
    .C(_00164_),
    .Y(_04379_));
 AO21x1_ASAP7_75t_R _11229_ (.A1(_00163_),
    .A2(_04001_),
    .B(_04379_),
    .Y(_04380_));
 AO221x1_ASAP7_75t_R _11230_ (.A1(_04076_),
    .A2(_04378_),
    .B1(_04380_),
    .B2(_04004_),
    .C(_03420_),
    .Y(_04381_));
 AND2x2_ASAP7_75t_R _11231_ (.A(_04014_),
    .B(_00158_),
    .Y(_04382_));
 AO21x1_ASAP7_75t_R _11232_ (.A1(_04274_),
    .A2(_00157_),
    .B(_04382_),
    .Y(_04383_));
 AND3x1_ASAP7_75t_R _11233_ (.A(_04014_),
    .B(_03970_),
    .C(_00156_),
    .Y(_04384_));
 AO21x1_ASAP7_75t_R _11234_ (.A1(_00155_),
    .A2(_04001_),
    .B(_04384_),
    .Y(_04385_));
 AO221x1_ASAP7_75t_R _11235_ (.A1(_04076_),
    .A2(_04383_),
    .B1(_04385_),
    .B2(_04004_),
    .C(_04297_),
    .Y(_04386_));
 AO22x1_ASAP7_75t_R _11236_ (.A1(_03956_),
    .A2(_00162_),
    .B1(_04020_),
    .B2(_00160_),
    .Y(_04387_));
 AND2x2_ASAP7_75t_R _11237_ (.A(_03923_),
    .B(_00154_),
    .Y(_04388_));
 AO221x1_ASAP7_75t_R _11238_ (.A1(_04111_),
    .A2(_03378_),
    .B1(_00152_),
    .B2(_04020_),
    .C(_04388_),
    .Y(_04389_));
 OA211x2_ASAP7_75t_R _11239_ (.A1(_03996_),
    .A2(_04387_),
    .B(_04389_),
    .C(_04256_),
    .Y(_04390_));
 AND2x2_ASAP7_75t_R _11240_ (.A(_03924_),
    .B(_00161_),
    .Y(_04391_));
 AO21x1_ASAP7_75t_R _11241_ (.A1(_04024_),
    .A2(_00159_),
    .B(_04391_),
    .Y(_04392_));
 AND2x2_ASAP7_75t_R _11242_ (.A(_03923_),
    .B(_00153_),
    .Y(_04393_));
 AO221x1_ASAP7_75t_R _11243_ (.A1(_03442_),
    .A2(_03378_),
    .B1(_00151_),
    .B2(_03953_),
    .C(_04393_),
    .Y(_04394_));
 OA211x2_ASAP7_75t_R _11244_ (.A1(_03996_),
    .A2(_04392_),
    .B(_04394_),
    .C(_03929_),
    .Y(_04395_));
 OR3x1_ASAP7_75t_R _11245_ (.A(_03981_),
    .B(_04390_),
    .C(_04395_),
    .Y(_04396_));
 AND3x1_ASAP7_75t_R _11246_ (.A(_04381_),
    .B(_04386_),
    .C(_04396_),
    .Y(_04397_));
 AND2x2_ASAP7_75t_R _11247_ (.A(_03973_),
    .B(_00145_),
    .Y(_04398_));
 AO21x1_ASAP7_75t_R _11248_ (.A1(_03991_),
    .A2(_00143_),
    .B(_04398_),
    .Y(_04399_));
 AO221x1_ASAP7_75t_R _11249_ (.A1(_04105_),
    .A2(_00146_),
    .B1(_04021_),
    .B2(_00144_),
    .C(_03929_),
    .Y(_04400_));
 OAI21x1_ASAP7_75t_R _11250_ (.A1(_04127_),
    .A2(_04399_),
    .B(_04400_),
    .Y(_04401_));
 INVx2_ASAP7_75t_R _11251_ (.A(_00149_),
    .Y(_04402_));
 BUFx10_ASAP7_75t_R _11252_ (.A(_03940_),
    .Y(_04403_));
 NAND2x1_ASAP7_75t_R _11253_ (.A(_04403_),
    .B(_00150_),
    .Y(_04404_));
 OA21x2_ASAP7_75t_R _11254_ (.A1(_04033_),
    .A2(_04402_),
    .B(_04404_),
    .Y(_04405_));
 BUFx12_ASAP7_75t_R _11255_ (.A(_03474_),
    .Y(_04406_));
 OA21x2_ASAP7_75t_R _11256_ (.A1(_04103_),
    .A2(_04405_),
    .B(_04406_),
    .Y(_04407_));
 INVx2_ASAP7_75t_R _11257_ (.A(_00148_),
    .Y(_04408_));
 OR3x1_ASAP7_75t_R _11258_ (.A(_04037_),
    .B(_03983_),
    .C(_04408_),
    .Y(_04409_));
 INVx1_ASAP7_75t_R _11259_ (.A(_00147_),
    .Y(_04410_));
 AO21x1_ASAP7_75t_R _11260_ (.A1(_03933_),
    .A2(_03379_),
    .B(_04410_),
    .Y(_04411_));
 AND2x6_ASAP7_75t_R _11261_ (.A(_03388_),
    .B(_03402_),
    .Y(_04412_));
 AO21x1_ASAP7_75t_R _11262_ (.A1(_04409_),
    .A2(_04411_),
    .B(_04412_),
    .Y(_04413_));
 BUFx12f_ASAP7_75t_R _11263_ (.A(_03996_),
    .Y(_04414_));
 AOI221x1_ASAP7_75t_R _11264_ (.A1(_04296_),
    .A2(_04401_),
    .B1(_04407_),
    .B2(_04413_),
    .C(_04414_),
    .Y(_04415_));
 AND2x2_ASAP7_75t_R _11265_ (.A(_03977_),
    .B(_00142_),
    .Y(_04416_));
 AO21x1_ASAP7_75t_R _11266_ (.A1(_03949_),
    .A2(_00141_),
    .B(_04416_),
    .Y(_04417_));
 AO21x1_ASAP7_75t_R _11267_ (.A1(_03974_),
    .A2(_04417_),
    .B(_03946_),
    .Y(_04418_));
 AND3x1_ASAP7_75t_R _11268_ (.A(_03941_),
    .B(_03970_),
    .C(_00140_),
    .Y(_04419_));
 OA21x2_ASAP7_75t_R _11269_ (.A1(_03985_),
    .A2(_03983_),
    .B(_00139_),
    .Y(_04420_));
 OA21x2_ASAP7_75t_R _11270_ (.A1(_04419_),
    .A2(_04420_),
    .B(_03937_),
    .Y(_04421_));
 AND2x2_ASAP7_75t_R _11271_ (.A(_03985_),
    .B(_00135_),
    .Y(_04422_));
 AND3x1_ASAP7_75t_R _11272_ (.A(_03941_),
    .B(_03378_),
    .C(_00136_),
    .Y(_04423_));
 OA21x2_ASAP7_75t_R _11273_ (.A1(_04422_),
    .A2(_04423_),
    .B(_03991_),
    .Y(_04424_));
 AND2x2_ASAP7_75t_R _11274_ (.A(_03940_),
    .B(_00138_),
    .Y(_04425_));
 AO21x1_ASAP7_75t_R _11275_ (.A1(_03928_),
    .A2(_00137_),
    .B(_04425_),
    .Y(_04426_));
 AO221x1_ASAP7_75t_R _11276_ (.A1(_03983_),
    .A2(_00135_),
    .B1(_04412_),
    .B2(_04426_),
    .C(_04406_),
    .Y(_04427_));
 OA222x2_ASAP7_75t_R _11277_ (.A1(_03413_),
    .A2(_03984_),
    .B1(_04418_),
    .B2(_04421_),
    .C1(_04424_),
    .C2(_04427_),
    .Y(_04428_));
 NAND2x2_ASAP7_75t_R _11278_ (.A(_03916_),
    .B(_03447_),
    .Y(_04429_));
 OR3x1_ASAP7_75t_R _11279_ (.A(_04415_),
    .B(_04428_),
    .C(_04429_),
    .Y(_04430_));
 OA21x2_ASAP7_75t_R _11280_ (.A1(_03916_),
    .A2(_04397_),
    .B(_04430_),
    .Y(_04431_));
 NOR2x1_ASAP7_75t_R _11281_ (.A(_04254_),
    .B(_04431_),
    .Y(_04432_));
 AOI21x1_ASAP7_75t_R _11282_ (.A1(_04250_),
    .A2(_10164_),
    .B(_04432_),
    .Y(_04433_));
 XNOR2x2_ASAP7_75t_R _11283_ (.A(_03538_),
    .B(_04433_),
    .Y(_09970_));
 INVx1_ASAP7_75t_R _11284_ (.A(_09970_),
    .Y(_09968_));
 BUFx12f_ASAP7_75t_R _11285_ (.A(_04236_),
    .Y(_04434_));
 BUFx12f_ASAP7_75t_R _11286_ (.A(_03614_),
    .Y(_04435_));
 BUFx10_ASAP7_75t_R _11287_ (.A(_04435_),
    .Y(_04436_));
 AND3x1_ASAP7_75t_R _11288_ (.A(_03376_),
    .B(_04436_),
    .C(_00142_),
    .Y(_04437_));
 AO21x1_ASAP7_75t_R _11289_ (.A1(_00141_),
    .A2(_04434_),
    .B(_04437_),
    .Y(_04438_));
 AND3x1_ASAP7_75t_R _11290_ (.A(_04244_),
    .B(_03793_),
    .C(_03652_),
    .Y(_04439_));
 BUFx10_ASAP7_75t_R _11291_ (.A(_04439_),
    .Y(_04440_));
 INVx1_ASAP7_75t_R _11292_ (.A(_00137_),
    .Y(_04441_));
 BUFx12f_ASAP7_75t_R _11293_ (.A(_04185_),
    .Y(_04442_));
 INVx3_ASAP7_75t_R _11294_ (.A(_00136_),
    .Y(_04443_));
 NAND2x1_ASAP7_75t_R _11295_ (.A(_03636_),
    .B(_00138_),
    .Y(_04444_));
 OA211x2_ASAP7_75t_R _11296_ (.A1(_03897_),
    .A2(_04443_),
    .B(_04444_),
    .C(_03664_),
    .Y(_04445_));
 AO21x1_ASAP7_75t_R _11297_ (.A1(_04441_),
    .A2(_04442_),
    .B(_04445_),
    .Y(_04446_));
 NAND2x1_ASAP7_75t_R _11298_ (.A(_03844_),
    .B(_04446_),
    .Y(_04447_));
 AO21x1_ASAP7_75t_R _11299_ (.A1(_03677_),
    .A2(_04344_),
    .B(_00135_),
    .Y(_04448_));
 OA211x2_ASAP7_75t_R _11300_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03885_),
    .C(_00140_),
    .Y(_04449_));
 AO21x1_ASAP7_75t_R _11301_ (.A1(_00139_),
    .A2(_03878_),
    .B(_04449_),
    .Y(_04450_));
 AO32x1_ASAP7_75t_R _11302_ (.A1(_03773_),
    .A2(_04447_),
    .A3(_04448_),
    .B1(_04450_),
    .B2(_03721_),
    .Y(_04451_));
 BUFx10_ASAP7_75t_R _11303_ (.A(_04195_),
    .Y(_04452_));
 AOI211x1_ASAP7_75t_R _11304_ (.A1(_04438_),
    .A2(_04440_),
    .B(_04451_),
    .C(_04452_),
    .Y(_04453_));
 BUFx10_ASAP7_75t_R _11305_ (.A(_03824_),
    .Y(_04454_));
 BUFx12f_ASAP7_75t_R _11306_ (.A(_03623_),
    .Y(_04455_));
 BUFx12_ASAP7_75t_R _11307_ (.A(_04210_),
    .Y(_04456_));
 BUFx12f_ASAP7_75t_R _11308_ (.A(_03683_),
    .Y(_04457_));
 AND2x2_ASAP7_75t_R _11309_ (.A(_03609_),
    .B(_00148_),
    .Y(_04458_));
 AO21x1_ASAP7_75t_R _11310_ (.A1(_04457_),
    .A2(_00144_),
    .B(_04458_),
    .Y(_04459_));
 BUFx16f_ASAP7_75t_R _11311_ (.A(_03672_),
    .Y(_04460_));
 AO22x1_ASAP7_75t_R _11312_ (.A1(_00147_),
    .A2(_04456_),
    .B1(_04459_),
    .B2(_04460_),
    .Y(_04461_));
 NAND2x1_ASAP7_75t_R _11313_ (.A(_04455_),
    .B(_04461_),
    .Y(_04462_));
 AO21x1_ASAP7_75t_R _11314_ (.A1(_04454_),
    .A2(_04462_),
    .B(_04163_),
    .Y(_04463_));
 NAND2x1_ASAP7_75t_R _11315_ (.A(_00143_),
    .B(_03750_),
    .Y(_04464_));
 AND3x1_ASAP7_75t_R _11316_ (.A(_00145_),
    .B(_03828_),
    .C(_03830_),
    .Y(_04465_));
 AOI221x1_ASAP7_75t_R _11317_ (.A1(_00150_),
    .A2(_04198_),
    .B1(_04199_),
    .B2(_00149_),
    .C(_04465_),
    .Y(_04466_));
 AOI21x1_ASAP7_75t_R _11318_ (.A1(_00146_),
    .A2(_03834_),
    .B(_03825_),
    .Y(_04467_));
 BUFx12f_ASAP7_75t_R _11319_ (.A(_03740_),
    .Y(_04468_));
 AO221x2_ASAP7_75t_R _11320_ (.A1(_04463_),
    .A2(_04464_),
    .B1(_04466_),
    .B2(_04467_),
    .C(_04468_),
    .Y(_04469_));
 AND2x2_ASAP7_75t_R _11321_ (.A(_03609_),
    .B(_00164_),
    .Y(_04470_));
 AO21x1_ASAP7_75t_R _11322_ (.A1(_04457_),
    .A2(_00160_),
    .B(_04470_),
    .Y(_04471_));
 AO22x1_ASAP7_75t_R _11323_ (.A1(_00163_),
    .A2(_04456_),
    .B1(_04471_),
    .B2(_03762_),
    .Y(_04472_));
 AND2x2_ASAP7_75t_R _11324_ (.A(_03376_),
    .B(_04472_),
    .Y(_04473_));
 OA21x2_ASAP7_75t_R _11325_ (.A1(_03794_),
    .A2(_04473_),
    .B(_03698_),
    .Y(_04474_));
 AND3x1_ASAP7_75t_R _11326_ (.A(_00159_),
    .B(_03750_),
    .C(_03698_),
    .Y(_04475_));
 BUFx10_ASAP7_75t_R _11327_ (.A(_04199_),
    .Y(_04476_));
 AND2x2_ASAP7_75t_R _11328_ (.A(_00161_),
    .B(_03830_),
    .Y(_04477_));
 BUFx10_ASAP7_75t_R _11329_ (.A(_03660_),
    .Y(_04478_));
 OA21x2_ASAP7_75t_R _11330_ (.A1(_03802_),
    .A2(_04477_),
    .B(_04478_),
    .Y(_04479_));
 AO21x1_ASAP7_75t_R _11331_ (.A1(_00165_),
    .A2(_04476_),
    .B(_04479_),
    .Y(_04480_));
 AND3x1_ASAP7_75t_R _11332_ (.A(_00162_),
    .B(_03836_),
    .C(_03735_),
    .Y(_04481_));
 OA21x2_ASAP7_75t_R _11333_ (.A1(_03667_),
    .A2(_03670_),
    .B(_00166_),
    .Y(_04482_));
 OA21x2_ASAP7_75t_R _11334_ (.A1(_04481_),
    .A2(_04482_),
    .B(_03774_),
    .Y(_04483_));
 OAI22x1_ASAP7_75t_R _11335_ (.A1(_04474_),
    .A2(_04475_),
    .B1(_04480_),
    .B2(_04483_),
    .Y(_04484_));
 INVx1_ASAP7_75t_R _11336_ (.A(_00157_),
    .Y(_04485_));
 AND2x2_ASAP7_75t_R _11337_ (.A(_04485_),
    .B(_03805_),
    .Y(_04486_));
 INVx1_ASAP7_75t_R _11338_ (.A(_00158_),
    .Y(_04487_));
 NAND2x1_ASAP7_75t_R _11339_ (.A(_03632_),
    .B(_00156_),
    .Y(_04488_));
 OA211x2_ASAP7_75t_R _11340_ (.A1(_03632_),
    .A2(_04487_),
    .B(_03886_),
    .C(_04488_),
    .Y(_04489_));
 AOI21x1_ASAP7_75t_R _11341_ (.A1(_03794_),
    .A2(_04486_),
    .B(_04489_),
    .Y(_04490_));
 NAND2x2_ASAP7_75t_R _11342_ (.A(_03827_),
    .B(_03647_),
    .Y(_04491_));
 BUFx10_ASAP7_75t_R _11343_ (.A(_04491_),
    .Y(_04492_));
 OA211x2_ASAP7_75t_R _11344_ (.A1(_00155_),
    .A2(_04492_),
    .B(_03653_),
    .C(_03518_),
    .Y(_04493_));
 AND2x2_ASAP7_75t_R _11345_ (.A(_03897_),
    .B(_00154_),
    .Y(_04494_));
 AO21x1_ASAP7_75t_R _11346_ (.A1(_03632_),
    .A2(_00152_),
    .B(_04494_),
    .Y(_04495_));
 OA222x2_ASAP7_75t_R _11347_ (.A1(_04163_),
    .A2(_03773_),
    .B1(_04495_),
    .B2(_03711_),
    .C1(_03865_),
    .C2(_00153_),
    .Y(_04496_));
 INVx2_ASAP7_75t_R _11348_ (.A(_00151_),
    .Y(_04497_));
 NAND2x1_ASAP7_75t_R _11349_ (.A(_04497_),
    .B(_03702_),
    .Y(_04498_));
 BUFx6f_ASAP7_75t_R _11350_ (.A(_03723_),
    .Y(_04499_));
 AOI221x1_ASAP7_75t_R _11351_ (.A1(_04490_),
    .A2(_04493_),
    .B1(_04496_),
    .B2(_04498_),
    .C(_04499_),
    .Y(_04500_));
 AO22x1_ASAP7_75t_R _11352_ (.A1(_04453_),
    .A2(_04469_),
    .B1(_04484_),
    .B2(_04500_),
    .Y(_04501_));
 BUFx4f_ASAP7_75t_R _11353_ (.A(_04501_),
    .Y(_09969_));
 BUFx12_ASAP7_75t_R _11354_ (.A(_04106_),
    .Y(_04502_));
 AO22x1_ASAP7_75t_R _11355_ (.A1(_04502_),
    .A2(_00191_),
    .B1(_04069_),
    .B2(_00189_),
    .Y(_04503_));
 BUFx6f_ASAP7_75t_R _11356_ (.A(_04023_),
    .Y(_04504_));
 AND2x2_ASAP7_75t_R _11357_ (.A(_03957_),
    .B(_00190_),
    .Y(_04505_));
 AO21x1_ASAP7_75t_R _11358_ (.A1(_03955_),
    .A2(_00188_),
    .B(_04505_),
    .Y(_04506_));
 AO221x1_ASAP7_75t_R _11359_ (.A1(_04504_),
    .A2(_00188_),
    .B1(_04506_),
    .B2(_04265_),
    .C(_04156_),
    .Y(_04507_));
 AO21x1_ASAP7_75t_R _11360_ (.A1(_04066_),
    .A2(_04503_),
    .B(_04507_),
    .Y(_04508_));
 AND2x2_ASAP7_75t_R _11361_ (.A(_04106_),
    .B(_00198_),
    .Y(_04509_));
 AO21x1_ASAP7_75t_R _11362_ (.A1(_04104_),
    .A2(_00196_),
    .B(_04509_),
    .Y(_04510_));
 AO21x1_ASAP7_75t_R _11363_ (.A1(_00199_),
    .A2(_03962_),
    .B(_04009_),
    .Y(_04511_));
 AO221x1_ASAP7_75t_R _11364_ (.A1(_00197_),
    .A2(_04083_),
    .B1(_04510_),
    .B2(_04080_),
    .C(_04511_),
    .Y(_04512_));
 AO21x1_ASAP7_75t_R _11365_ (.A1(_04508_),
    .A2(_04512_),
    .B(_04095_),
    .Y(_04513_));
 BUFx6f_ASAP7_75t_R _11366_ (.A(_04414_),
    .Y(_04514_));
 AND3x1_ASAP7_75t_R _11367_ (.A(_04016_),
    .B(_03927_),
    .C(_00195_),
    .Y(_04515_));
 AND2x2_ASAP7_75t_R _11368_ (.A(_04075_),
    .B(_00194_),
    .Y(_04516_));
 AO21x1_ASAP7_75t_R _11369_ (.A1(_03955_),
    .A2(_00192_),
    .B(_04516_),
    .Y(_04517_));
 AO32x1_ASAP7_75t_R _11370_ (.A1(_04114_),
    .A2(_00193_),
    .A3(_04102_),
    .B1(_04517_),
    .B2(_03951_),
    .Y(_04518_));
 OR3x1_ASAP7_75t_R _11371_ (.A(_04514_),
    .B(_04515_),
    .C(_04518_),
    .Y(_04519_));
 BUFx12_ASAP7_75t_R _11372_ (.A(_04024_),
    .Y(_04520_));
 BUFx6f_ASAP7_75t_R _11373_ (.A(_04520_),
    .Y(_04521_));
 BUFx6f_ASAP7_75t_R _11374_ (.A(_03989_),
    .Y(_04522_));
 AND2x2_ASAP7_75t_R _11375_ (.A(_04105_),
    .B(_00186_),
    .Y(_04523_));
 AO21x1_ASAP7_75t_R _11376_ (.A1(_04073_),
    .A2(_00184_),
    .B(_04523_),
    .Y(_04524_));
 AO32x1_ASAP7_75t_R _11377_ (.A1(_04521_),
    .A2(_00185_),
    .A3(_04522_),
    .B1(_04524_),
    .B2(_04088_),
    .Y(_04525_));
 AO221x1_ASAP7_75t_R _11378_ (.A1(_04112_),
    .A2(_03381_),
    .B1(_00187_),
    .B2(_04091_),
    .C(_04525_),
    .Y(_04526_));
 AO21x1_ASAP7_75t_R _11379_ (.A1(_04519_),
    .A2(_04526_),
    .B(_04120_),
    .Y(_04527_));
 AO21x1_ASAP7_75t_R _11380_ (.A1(_04513_),
    .A2(_04527_),
    .B(_04122_),
    .Y(_04528_));
 BUFx10_ASAP7_75t_R _11381_ (.A(_03957_),
    .Y(_04529_));
 BUFx10_ASAP7_75t_R _11382_ (.A(_04529_),
    .Y(_04530_));
 BUFx12_ASAP7_75t_R _11383_ (.A(_03986_),
    .Y(_04531_));
 BUFx10_ASAP7_75t_R _11384_ (.A(_04403_),
    .Y(_04532_));
 AND2x2_ASAP7_75t_R _11385_ (.A(_04532_),
    .B(_00183_),
    .Y(_04533_));
 AO21x1_ASAP7_75t_R _11386_ (.A1(_04531_),
    .A2(_00182_),
    .B(_04533_),
    .Y(_04534_));
 BUFx12_ASAP7_75t_R _11387_ (.A(_04001_),
    .Y(_04535_));
 BUFx6f_ASAP7_75t_R _11388_ (.A(_03977_),
    .Y(_04536_));
 BUFx10_ASAP7_75t_R _11389_ (.A(_04536_),
    .Y(_04537_));
 AND3x1_ASAP7_75t_R _11390_ (.A(_04537_),
    .B(_03971_),
    .C(_00181_),
    .Y(_04538_));
 AO21x1_ASAP7_75t_R _11391_ (.A1(_00180_),
    .A2(_04535_),
    .B(_04538_),
    .Y(_04539_));
 BUFx10_ASAP7_75t_R _11392_ (.A(_04004_),
    .Y(_04540_));
 BUFx4f_ASAP7_75t_R _11393_ (.A(_03449_),
    .Y(_04541_));
 BUFx6f_ASAP7_75t_R _11394_ (.A(_04541_),
    .Y(_04542_));
 AO221x2_ASAP7_75t_R _11395_ (.A1(_04530_),
    .A2(_04534_),
    .B1(_04539_),
    .B2(_04540_),
    .C(_04542_),
    .Y(_04543_));
 BUFx10_ASAP7_75t_R _11396_ (.A(_04043_),
    .Y(_04544_));
 AND2x2_ASAP7_75t_R _11397_ (.A(_04544_),
    .B(_00178_),
    .Y(_04545_));
 AO21x1_ASAP7_75t_R _11398_ (.A1(_04084_),
    .A2(_00176_),
    .B(_04545_),
    .Y(_04546_));
 AO21x1_ASAP7_75t_R _11399_ (.A1(_00177_),
    .A2(_03964_),
    .B(_04130_),
    .Y(_04547_));
 AO221x1_ASAP7_75t_R _11400_ (.A1(_00179_),
    .A2(_03962_),
    .B1(_04546_),
    .B2(_04136_),
    .C(_04547_),
    .Y(_04548_));
 AND3x1_ASAP7_75t_R _11401_ (.A(_04157_),
    .B(_04543_),
    .C(_04548_),
    .Y(_04549_));
 AND2x2_ASAP7_75t_R _11402_ (.A(_03933_),
    .B(_00171_),
    .Y(_04550_));
 AO21x1_ASAP7_75t_R _11403_ (.A1(_04125_),
    .A2(_00170_),
    .B(_04550_),
    .Y(_04551_));
 AO21x1_ASAP7_75t_R _11404_ (.A1(_03927_),
    .A2(_04551_),
    .B(_04032_),
    .Y(_04552_));
 AO22x1_ASAP7_75t_R _11405_ (.A1(_03950_),
    .A2(_00168_),
    .B1(_00169_),
    .B2(_04101_),
    .Y(_04553_));
 AO22x1_ASAP7_75t_R _11406_ (.A1(_04071_),
    .A2(_00168_),
    .B1(_04553_),
    .B2(_04521_),
    .Y(_04554_));
 AO21x1_ASAP7_75t_R _11407_ (.A1(_03381_),
    .A2(_04552_),
    .B(_04554_),
    .Y(_04555_));
 BUFx10_ASAP7_75t_R _11408_ (.A(_04274_),
    .Y(_04556_));
 AND2x2_ASAP7_75t_R _11409_ (.A(_04015_),
    .B(_00175_),
    .Y(_04557_));
 AO21x1_ASAP7_75t_R _11410_ (.A1(_04556_),
    .A2(_00174_),
    .B(_04557_),
    .Y(_04558_));
 BUFx12_ASAP7_75t_R _11411_ (.A(_03970_),
    .Y(_04559_));
 AND3x1_ASAP7_75t_R _11412_ (.A(_04532_),
    .B(_04559_),
    .C(_00173_),
    .Y(_04560_));
 AO21x1_ASAP7_75t_R _11413_ (.A1(_00172_),
    .A2(_04535_),
    .B(_04560_),
    .Y(_04561_));
 AO221x1_ASAP7_75t_R _11414_ (.A1(_04530_),
    .A2(_04558_),
    .B1(_04561_),
    .B2(_04540_),
    .C(_04542_),
    .Y(_04562_));
 AND3x2_ASAP7_75t_R _11415_ (.A(_04099_),
    .B(_04555_),
    .C(_04562_),
    .Y(_04563_));
 OR3x1_ASAP7_75t_R _11416_ (.A(_04124_),
    .B(_04549_),
    .C(_04563_),
    .Y(_04564_));
 BUFx12_ASAP7_75t_R _11417_ (.A(_04055_),
    .Y(_04565_));
 AO21x2_ASAP7_75t_R _11418_ (.A1(_04528_),
    .A2(_04564_),
    .B(_04565_),
    .Y(_04566_));
 AND3x1_ASAP7_75t_R _11419_ (.A(_03382_),
    .B(net18),
    .C(_03600_),
    .Y(_04567_));
 OA21x2_ASAP7_75t_R _11420_ (.A1(_04251_),
    .A2(_04567_),
    .B(_04168_),
    .Y(_10162_));
 NAND2x1_ASAP7_75t_R _11421_ (.A(_04254_),
    .B(_10162_),
    .Y(_04568_));
 OAI21x1_ASAP7_75t_R _11422_ (.A1(_04250_),
    .A2(_04566_),
    .B(_04568_),
    .Y(_04569_));
 XNOR2x1_ASAP7_75t_R _11423_ (.B(_04569_),
    .Y(_09975_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _11424_ (.A(_09975_),
    .Y(_09973_));
 AO221x1_ASAP7_75t_R _11425_ (.A1(_00199_),
    .A2(_04198_),
    .B1(_03833_),
    .B2(_00195_),
    .C(_04454_),
    .Y(_04570_));
 AND3x1_ASAP7_75t_R _11426_ (.A(_00194_),
    .B(_03737_),
    .C(_03735_),
    .Y(_04571_));
 OA21x2_ASAP7_75t_R _11427_ (.A1(_03667_),
    .A2(_03670_),
    .B(_00198_),
    .Y(_04572_));
 OA21x2_ASAP7_75t_R _11428_ (.A1(_04571_),
    .A2(_04572_),
    .B(_03782_),
    .Y(_04573_));
 INVx1_ASAP7_75t_R _11429_ (.A(_00192_),
    .Y(_04574_));
 BUFx16f_ASAP7_75t_R _11430_ (.A(_04206_),
    .Y(_04575_));
 BUFx16f_ASAP7_75t_R _11431_ (.A(_04210_),
    .Y(_04576_));
 AND2x2_ASAP7_75t_R _11432_ (.A(_03609_),
    .B(_00197_),
    .Y(_04577_));
 AO21x1_ASAP7_75t_R _11433_ (.A1(_04457_),
    .A2(_00193_),
    .B(_04577_),
    .Y(_04578_));
 AOI22x1_ASAP7_75t_R _11434_ (.A1(_00196_),
    .A2(_04576_),
    .B1(_04578_),
    .B2(_03762_),
    .Y(_04579_));
 OA211x2_ASAP7_75t_R _11435_ (.A1(_03839_),
    .A2(_04579_),
    .B(_03775_),
    .C(_03828_),
    .Y(_04580_));
 OAI22x1_ASAP7_75t_R _11436_ (.A1(_04574_),
    .A2(_04575_),
    .B1(_04580_),
    .B2(_03785_),
    .Y(_04581_));
 OA211x2_ASAP7_75t_R _11437_ (.A1(_04570_),
    .A2(_04573_),
    .B(_03868_),
    .C(_04581_),
    .Y(_04582_));
 BUFx6f_ASAP7_75t_R _11438_ (.A(_03659_),
    .Y(_04583_));
 BUFx12f_ASAP7_75t_R _11439_ (.A(_03624_),
    .Y(_04584_));
 AND3x1_ASAP7_75t_R _11440_ (.A(_04455_),
    .B(_04584_),
    .C(_00191_),
    .Y(_04585_));
 AO21x1_ASAP7_75t_R _11441_ (.A1(_00190_),
    .A2(_03782_),
    .B(_04585_),
    .Y(_04586_));
 BUFx6f_ASAP7_75t_R _11442_ (.A(_03731_),
    .Y(_04587_));
 AND2x2_ASAP7_75t_R _11443_ (.A(_00188_),
    .B(_03585_),
    .Y(_04588_));
 AO221x1_ASAP7_75t_R _11444_ (.A1(_00189_),
    .A2(_03813_),
    .B1(_04587_),
    .B2(_03518_),
    .C(_04588_),
    .Y(_04589_));
 OA211x2_ASAP7_75t_R _11445_ (.A1(_04583_),
    .A2(_04586_),
    .B(_04589_),
    .C(_03791_),
    .Y(_04590_));
 BUFx10_ASAP7_75t_R _11446_ (.A(_03813_),
    .Y(_04591_));
 BUFx10_ASAP7_75t_R _11447_ (.A(_03775_),
    .Y(_04592_));
 AO32x1_ASAP7_75t_R _11448_ (.A1(_00185_),
    .A2(_04591_),
    .A3(_04592_),
    .B1(_03702_),
    .B2(_00184_),
    .Y(_04593_));
 AND2x2_ASAP7_75t_R _11449_ (.A(_03701_),
    .B(_04593_),
    .Y(_04594_));
 BUFx10_ASAP7_75t_R _11450_ (.A(_04242_),
    .Y(_04595_));
 BUFx12f_ASAP7_75t_R _11451_ (.A(_03375_),
    .Y(_04596_));
 BUFx12f_ASAP7_75t_R _11452_ (.A(_04435_),
    .Y(_04597_));
 AND3x1_ASAP7_75t_R _11453_ (.A(_04596_),
    .B(_04597_),
    .C(_00187_),
    .Y(_04598_));
 AO21x1_ASAP7_75t_R _11454_ (.A1(_00186_),
    .A2(_04595_),
    .B(_04598_),
    .Y(_04599_));
 AND3x1_ASAP7_75t_R _11455_ (.A(_03733_),
    .B(_03701_),
    .C(_04599_),
    .Y(_04600_));
 OR5x2_ASAP7_75t_R _11456_ (.A(_03809_),
    .B(_04582_),
    .C(_04590_),
    .D(_04594_),
    .E(_04600_),
    .Y(_04601_));
 BUFx6f_ASAP7_75t_R _11457_ (.A(_03871_),
    .Y(_04602_));
 AO21x1_ASAP7_75t_R _11458_ (.A1(_00178_),
    .A2(_03830_),
    .B(_03802_),
    .Y(_04603_));
 AO32x1_ASAP7_75t_R _11459_ (.A1(_00182_),
    .A2(_04595_),
    .A3(_04602_),
    .B1(_04603_),
    .B2(_03829_),
    .Y(_04604_));
 AND3x1_ASAP7_75t_R _11460_ (.A(_00179_),
    .B(_03836_),
    .C(_03735_),
    .Y(_04605_));
 OA21x2_ASAP7_75t_R _11461_ (.A1(_03667_),
    .A2(_03670_),
    .B(_00183_),
    .Y(_04606_));
 OA21x2_ASAP7_75t_R _11462_ (.A1(_04605_),
    .A2(_04606_),
    .B(_03774_),
    .Y(_04607_));
 INVx1_ASAP7_75t_R _11463_ (.A(_00176_),
    .Y(_04608_));
 BUFx16f_ASAP7_75t_R _11464_ (.A(_03744_),
    .Y(_04609_));
 BUFx12f_ASAP7_75t_R _11465_ (.A(_03685_),
    .Y(_04610_));
 AND2x2_ASAP7_75t_R _11466_ (.A(_04610_),
    .B(_00181_),
    .Y(_04611_));
 AO21x1_ASAP7_75t_R _11467_ (.A1(_04609_),
    .A2(_00177_),
    .B(_04611_),
    .Y(_04612_));
 AOI22x1_ASAP7_75t_R _11468_ (.A1(_00180_),
    .A2(_04576_),
    .B1(_04612_),
    .B2(_03665_),
    .Y(_04613_));
 OA211x2_ASAP7_75t_R _11469_ (.A1(_03481_),
    .A2(_04613_),
    .B(_03802_),
    .C(_03836_),
    .Y(_04614_));
 OAI22x1_ASAP7_75t_R _11470_ (.A1(_04608_),
    .A2(_04575_),
    .B1(_04614_),
    .B2(_04164_),
    .Y(_04615_));
 OA211x2_ASAP7_75t_R _11471_ (.A1(_04604_),
    .A2(_04607_),
    .B(_03868_),
    .C(_04615_),
    .Y(_04616_));
 AND4x1_ASAP7_75t_R _11472_ (.A(_00175_),
    .B(_03677_),
    .C(_03516_),
    .D(_03731_),
    .Y(_04617_));
 AO21x1_ASAP7_75t_R _11473_ (.A1(_00173_),
    .A2(_03659_),
    .B(_04617_),
    .Y(_04618_));
 OA211x2_ASAP7_75t_R _11474_ (.A1(_00172_),
    .A2(_04492_),
    .B(_03653_),
    .C(_03518_),
    .Y(_04619_));
 OA221x2_ASAP7_75t_R _11475_ (.A1(_00174_),
    .A2(_03866_),
    .B1(_04618_),
    .B2(_03879_),
    .C(_04619_),
    .Y(_04620_));
 OR3x4_ASAP7_75t_R _11476_ (.A(_04452_),
    .B(_04616_),
    .C(_04620_),
    .Y(_04621_));
 AND2x4_ASAP7_75t_R _11477_ (.A(_03878_),
    .B(_03601_),
    .Y(_04622_));
 BUFx12_ASAP7_75t_R _11478_ (.A(_04434_),
    .Y(_04623_));
 BUFx10_ASAP7_75t_R _11479_ (.A(_04597_),
    .Y(_04624_));
 AND3x1_ASAP7_75t_R _11480_ (.A(_04053_),
    .B(_04624_),
    .C(_00171_),
    .Y(_04625_));
 AO21x1_ASAP7_75t_R _11481_ (.A1(_00170_),
    .A2(_04623_),
    .B(_04625_),
    .Y(_04626_));
 BUFx6f_ASAP7_75t_R _11482_ (.A(_04193_),
    .Y(_04627_));
 AND2x6_ASAP7_75t_R _11483_ (.A(_03813_),
    .B(_03607_),
    .Y(_04628_));
 AND2x4_ASAP7_75t_R _11484_ (.A(_04627_),
    .B(_04628_),
    .Y(_04629_));
 AO222x2_ASAP7_75t_R _11485_ (.A1(_00168_),
    .A2(_04622_),
    .B1(_03901_),
    .B2(_04626_),
    .C1(_04629_),
    .C2(_00169_),
    .Y(_04630_));
 AO21x2_ASAP7_75t_R _11486_ (.A1(_04601_),
    .A2(_04621_),
    .B(_04630_),
    .Y(_09972_));
 INVx3_ASAP7_75t_R _11487_ (.A(_09972_),
    .Y(_09974_));
 AND3x1_ASAP7_75t_R _11488_ (.A(net89),
    .B(net17),
    .C(_03600_),
    .Y(_04631_));
 OA21x2_ASAP7_75t_R _11489_ (.A1(_04251_),
    .A2(_04631_),
    .B(_04253_),
    .Y(_10160_));
 BUFx6f_ASAP7_75t_R _11490_ (.A(_04021_),
    .Y(_04632_));
 AO22x1_ASAP7_75t_R _11491_ (.A1(_04255_),
    .A2(_00225_),
    .B1(_04632_),
    .B2(_00223_),
    .Y(_04633_));
 AND2x2_ASAP7_75t_R _11492_ (.A(_03925_),
    .B(_00224_),
    .Y(_04634_));
 AO21x1_ASAP7_75t_R _11493_ (.A1(_04103_),
    .A2(_00222_),
    .B(_04634_),
    .Y(_04635_));
 AO221x1_ASAP7_75t_R _11494_ (.A1(_04071_),
    .A2(_00222_),
    .B1(_04635_),
    .B2(_04079_),
    .C(_03920_),
    .Y(_04636_));
 AO21x1_ASAP7_75t_R _11495_ (.A1(_04066_),
    .A2(_04633_),
    .B(_04636_),
    .Y(_04637_));
 AND2x2_ASAP7_75t_R _11496_ (.A(_04018_),
    .B(_00232_),
    .Y(_04638_));
 AO21x1_ASAP7_75t_R _11497_ (.A1(_04521_),
    .A2(_00230_),
    .B(_04638_),
    .Y(_04639_));
 AO21x1_ASAP7_75t_R _11498_ (.A1(_00233_),
    .A2(_04262_),
    .B(_04009_),
    .Y(_04640_));
 AO221x1_ASAP7_75t_R _11499_ (.A1(_00231_),
    .A2(_04083_),
    .B1(_04639_),
    .B2(_04136_),
    .C(_04640_),
    .Y(_04641_));
 AO21x1_ASAP7_75t_R _11500_ (.A1(_04637_),
    .A2(_04641_),
    .B(_04095_),
    .Y(_04642_));
 BUFx6f_ASAP7_75t_R _11501_ (.A(_04544_),
    .Y(_04643_));
 AND3x1_ASAP7_75t_R _11502_ (.A(_04016_),
    .B(_04643_),
    .C(_00229_),
    .Y(_04644_));
 AND2x2_ASAP7_75t_R _11503_ (.A(_03925_),
    .B(_00228_),
    .Y(_04645_));
 AO21x1_ASAP7_75t_R _11504_ (.A1(_04113_),
    .A2(_00226_),
    .B(_04645_),
    .Y(_04646_));
 BUFx6f_ASAP7_75t_R _11505_ (.A(_04274_),
    .Y(_04647_));
 AO32x1_ASAP7_75t_R _11506_ (.A1(_04521_),
    .A2(_00227_),
    .A3(_04522_),
    .B1(_04646_),
    .B2(_04647_),
    .Y(_04648_));
 OR3x1_ASAP7_75t_R _11507_ (.A(_04098_),
    .B(_04644_),
    .C(_04648_),
    .Y(_04649_));
 AND2x2_ASAP7_75t_R _11508_ (.A(_04017_),
    .B(_00220_),
    .Y(_04650_));
 AO21x1_ASAP7_75t_R _11509_ (.A1(_04520_),
    .A2(_00218_),
    .B(_04650_),
    .Y(_04651_));
 AO32x1_ASAP7_75t_R _11510_ (.A1(_04084_),
    .A2(_00219_),
    .A3(_04522_),
    .B1(_04651_),
    .B2(_04556_),
    .Y(_04652_));
 AO221x1_ASAP7_75t_R _11511_ (.A1(_04112_),
    .A2(_03381_),
    .B1(_00221_),
    .B2(_04091_),
    .C(_04652_),
    .Y(_04653_));
 AO21x1_ASAP7_75t_R _11512_ (.A1(_04649_),
    .A2(_04653_),
    .B(_04120_),
    .Y(_04654_));
 AOI21x1_ASAP7_75t_R _11513_ (.A1(_04642_),
    .A2(_04654_),
    .B(_04122_),
    .Y(_04655_));
 BUFx10_ASAP7_75t_R _11514_ (.A(_04270_),
    .Y(_04656_));
 AND2x2_ASAP7_75t_R _11515_ (.A(_04307_),
    .B(_00205_),
    .Y(_04657_));
 AO21x1_ASAP7_75t_R _11516_ (.A1(_03951_),
    .A2(_00204_),
    .B(_04657_),
    .Y(_04658_));
 AO21x1_ASAP7_75t_R _11517_ (.A1(_04656_),
    .A2(_04658_),
    .B(_04119_),
    .Y(_04659_));
 AO22x1_ASAP7_75t_R _11518_ (.A1(_04647_),
    .A2(_00202_),
    .B1(_00203_),
    .B2(_04522_),
    .Y(_04660_));
 AO22x1_ASAP7_75t_R _11519_ (.A1(_04504_),
    .A2(_00202_),
    .B1(_04660_),
    .B2(_04085_),
    .Y(_04661_));
 AO21x1_ASAP7_75t_R _11520_ (.A1(_04060_),
    .A2(_04659_),
    .B(_04661_),
    .Y(_04662_));
 BUFx12_ASAP7_75t_R _11521_ (.A(_03998_),
    .Y(_04663_));
 AND2x2_ASAP7_75t_R _11522_ (.A(_04137_),
    .B(_00209_),
    .Y(_04664_));
 AO21x1_ASAP7_75t_R _11523_ (.A1(_04663_),
    .A2(_00208_),
    .B(_04664_),
    .Y(_04665_));
 BUFx10_ASAP7_75t_R _11524_ (.A(_03941_),
    .Y(_04666_));
 AND3x1_ASAP7_75t_R _11525_ (.A(_04666_),
    .B(_03943_),
    .C(_00207_),
    .Y(_04667_));
 AO21x1_ASAP7_75t_R _11526_ (.A1(_00206_),
    .A2(_04292_),
    .B(_04667_),
    .Y(_04668_));
 AO221x1_ASAP7_75t_R _11527_ (.A1(_04289_),
    .A2(_04665_),
    .B1(_04668_),
    .B2(_04295_),
    .C(_04094_),
    .Y(_04669_));
 AND2x2_ASAP7_75t_R _11528_ (.A(_04514_),
    .B(_04669_),
    .Y(_04670_));
 BUFx10_ASAP7_75t_R _11529_ (.A(_03998_),
    .Y(_04671_));
 AND2x2_ASAP7_75t_R _11530_ (.A(_04666_),
    .B(_00217_),
    .Y(_04672_));
 AO21x1_ASAP7_75t_R _11531_ (.A1(_04671_),
    .A2(_00216_),
    .B(_04672_),
    .Y(_04673_));
 AND3x1_ASAP7_75t_R _11532_ (.A(_04015_),
    .B(_04559_),
    .C(_00215_),
    .Y(_04674_));
 AO21x1_ASAP7_75t_R _11533_ (.A1(_00214_),
    .A2(_04292_),
    .B(_04674_),
    .Y(_04675_));
 AO221x1_ASAP7_75t_R _11534_ (.A1(_04502_),
    .A2(_04673_),
    .B1(_04675_),
    .B2(_04295_),
    .C(_04094_),
    .Y(_04676_));
 AND2x2_ASAP7_75t_R _11535_ (.A(_03974_),
    .B(_00212_),
    .Y(_04677_));
 AO21x1_ASAP7_75t_R _11536_ (.A1(_03992_),
    .A2(_00210_),
    .B(_04677_),
    .Y(_04678_));
 AO21x1_ASAP7_75t_R _11537_ (.A1(_00211_),
    .A2(_03964_),
    .B(_03981_),
    .Y(_04679_));
 AO221x1_ASAP7_75t_R _11538_ (.A1(_00213_),
    .A2(_03962_),
    .B1(_04678_),
    .B2(_04126_),
    .C(_04679_),
    .Y(_04680_));
 AND3x1_ASAP7_75t_R _11539_ (.A(_04157_),
    .B(_04676_),
    .C(_04680_),
    .Y(_04681_));
 AOI211x1_ASAP7_75t_R _11540_ (.A1(_04662_),
    .A2(_04670_),
    .B(_04124_),
    .C(_04681_),
    .Y(_04682_));
 OA21x2_ASAP7_75t_R _11541_ (.A1(_04655_),
    .A2(_04682_),
    .B(_03447_),
    .Y(_04683_));
 AND2x2_ASAP7_75t_R _11542_ (.A(_04059_),
    .B(_04683_),
    .Y(_04684_));
 AO21x1_ASAP7_75t_R _11543_ (.A1(_04250_),
    .A2(_10160_),
    .B(_04684_),
    .Y(_04685_));
 XNOR2x1_ASAP7_75t_R _11544_ (.B(_04685_),
    .Y(_09980_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _11545_ (.A(_09980_),
    .Y(_09978_));
 INVx1_ASAP7_75t_R _11546_ (.A(_00226_),
    .Y(_04686_));
 AND2x2_ASAP7_75t_R _11547_ (.A(_03685_),
    .B(_00231_),
    .Y(_04687_));
 AO21x1_ASAP7_75t_R _11548_ (.A1(_03744_),
    .A2(_00227_),
    .B(_04687_),
    .Y(_04688_));
 AOI22x1_ASAP7_75t_R _11549_ (.A1(_00230_),
    .A2(_04456_),
    .B1(_04688_),
    .B2(_03664_),
    .Y(_04689_));
 OA211x2_ASAP7_75t_R _11550_ (.A1(_03480_),
    .A2(_04689_),
    .B(_04212_),
    .C(_04350_),
    .Y(_04690_));
 OAI22x1_ASAP7_75t_R _11551_ (.A1(_04686_),
    .A2(_04218_),
    .B1(_04690_),
    .B2(_04163_),
    .Y(_04691_));
 AND3x1_ASAP7_75t_R _11552_ (.A(_03402_),
    .B(_03633_),
    .C(_00229_),
    .Y(_04692_));
 AO21x1_ASAP7_75t_R _11553_ (.A1(_00228_),
    .A2(_03709_),
    .B(_04692_),
    .Y(_04693_));
 OR3x1_ASAP7_75t_R _11554_ (.A(_04233_),
    .B(_03669_),
    .C(_04693_),
    .Y(_04694_));
 AND2x2_ASAP7_75t_R _11555_ (.A(_00232_),
    .B(_03709_),
    .Y(_04695_));
 AO221x1_ASAP7_75t_R _11556_ (.A1(_00233_),
    .A2(_03727_),
    .B1(_03734_),
    .B2(_03736_),
    .C(_04695_),
    .Y(_04696_));
 AO21x1_ASAP7_75t_R _11557_ (.A1(_04694_),
    .A2(_04696_),
    .B(_04229_),
    .Y(_04697_));
 OA211x2_ASAP7_75t_R _11558_ (.A1(_03723_),
    .A2(_04691_),
    .B(_04697_),
    .C(_04231_),
    .Y(_04698_));
 OR3x1_ASAP7_75t_R _11559_ (.A(_00219_),
    .B(_04233_),
    .C(_03681_),
    .Y(_04699_));
 AO21x1_ASAP7_75t_R _11560_ (.A1(_03860_),
    .A2(_03801_),
    .B(_00221_),
    .Y(_04700_));
 AO21x1_ASAP7_75t_R _11561_ (.A1(_04699_),
    .A2(_04700_),
    .B(_03761_),
    .Y(_04701_));
 OR2x2_ASAP7_75t_R _11562_ (.A(_00220_),
    .B(_03865_),
    .Y(_04702_));
 OA21x2_ASAP7_75t_R _11563_ (.A1(_00218_),
    .A2(_03759_),
    .B(_03700_),
    .Y(_04703_));
 OR3x1_ASAP7_75t_R _11564_ (.A(_00223_),
    .B(_04233_),
    .C(_03680_),
    .Y(_04704_));
 AO21x1_ASAP7_75t_R _11565_ (.A1(_03860_),
    .A2(_03801_),
    .B(_00225_),
    .Y(_04705_));
 AO21x1_ASAP7_75t_R _11566_ (.A1(_04704_),
    .A2(_04705_),
    .B(_04236_),
    .Y(_04706_));
 OR3x1_ASAP7_75t_R _11567_ (.A(_00222_),
    .B(_03605_),
    .C(_04344_),
    .Y(_04707_));
 AO221x1_ASAP7_75t_R _11568_ (.A1(_03443_),
    .A2(_03716_),
    .B1(_03645_),
    .B2(_03593_),
    .C(_00224_),
    .Y(_04708_));
 AND4x1_ASAP7_75t_R _11569_ (.A(_04244_),
    .B(_03652_),
    .C(_04707_),
    .D(_04708_),
    .Y(_04709_));
 AO32x2_ASAP7_75t_R _11570_ (.A1(_04701_),
    .A2(_04702_),
    .A3(_04703_),
    .B1(_04706_),
    .B2(_04709_),
    .Y(_04710_));
 AO21x1_ASAP7_75t_R _11571_ (.A1(_00212_),
    .A2(_03830_),
    .B(_04212_),
    .Y(_04711_));
 AO32x1_ASAP7_75t_R _11572_ (.A1(_00216_),
    .A2(_03781_),
    .A3(_03871_),
    .B1(_04711_),
    .B2(_03828_),
    .Y(_04712_));
 AND3x1_ASAP7_75t_R _11573_ (.A(_00213_),
    .B(_03736_),
    .C(_03734_),
    .Y(_04713_));
 OA21x2_ASAP7_75t_R _11574_ (.A1(_04233_),
    .A2(_03669_),
    .B(_00217_),
    .Y(_04714_));
 OA21x2_ASAP7_75t_R _11575_ (.A1(_04713_),
    .A2(_04714_),
    .B(_03728_),
    .Y(_04715_));
 INVx1_ASAP7_75t_R _11576_ (.A(_00210_),
    .Y(_04716_));
 AND2x2_ASAP7_75t_R _11577_ (.A(_03608_),
    .B(_00215_),
    .Y(_04717_));
 AO21x1_ASAP7_75t_R _11578_ (.A1(_03683_),
    .A2(_00211_),
    .B(_04717_),
    .Y(_04718_));
 AOI22x1_ASAP7_75t_R _11579_ (.A1(_00214_),
    .A2(_04210_),
    .B1(_04718_),
    .B2(_03664_),
    .Y(_04719_));
 OA211x2_ASAP7_75t_R _11580_ (.A1(_03419_),
    .A2(_04719_),
    .B(_04212_),
    .C(_03736_),
    .Y(_04720_));
 OAI22x1_ASAP7_75t_R _11581_ (.A1(_04716_),
    .A2(_04218_),
    .B1(_04720_),
    .B2(_04214_),
    .Y(_04721_));
 OA211x2_ASAP7_75t_R _11582_ (.A1(_04712_),
    .A2(_04715_),
    .B(_03698_),
    .C(_04721_),
    .Y(_04722_));
 INVx1_ASAP7_75t_R _11583_ (.A(_00208_),
    .Y(_04723_));
 INVx1_ASAP7_75t_R _11584_ (.A(_00209_),
    .Y(_04724_));
 AOI22x1_ASAP7_75t_R _11585_ (.A1(_04723_),
    .A2(_03671_),
    .B1(_03813_),
    .B2(_04724_),
    .Y(_04725_));
 AND4x1_ASAP7_75t_R _11586_ (.A(_04244_),
    .B(_03794_),
    .C(_03652_),
    .D(_04725_),
    .Y(_04726_));
 BUFx10_ASAP7_75t_R _11587_ (.A(_03720_),
    .Y(_04727_));
 AND3x1_ASAP7_75t_R _11588_ (.A(_03374_),
    .B(_03672_),
    .C(_00207_),
    .Y(_04728_));
 AO21x1_ASAP7_75t_R _11589_ (.A1(_00206_),
    .A2(_03612_),
    .B(_04728_),
    .Y(_04729_));
 AND3x1_ASAP7_75t_R _11590_ (.A(_03677_),
    .B(_04727_),
    .C(_04729_),
    .Y(_04730_));
 INVx1_ASAP7_75t_R _11591_ (.A(_00204_),
    .Y(_04731_));
 INVx1_ASAP7_75t_R _11592_ (.A(_00203_),
    .Y(_04732_));
 NAND2x1_ASAP7_75t_R _11593_ (.A(_03591_),
    .B(_00205_),
    .Y(_04733_));
 OA211x2_ASAP7_75t_R _11594_ (.A1(_03619_),
    .A2(_04732_),
    .B(_04733_),
    .C(_03613_),
    .Y(_04734_));
 AOI21x1_ASAP7_75t_R _11595_ (.A1(_04731_),
    .A2(_04185_),
    .B(_04734_),
    .Y(_04735_));
 OA211x2_ASAP7_75t_R _11596_ (.A1(_03628_),
    .A2(_04735_),
    .B(_03771_),
    .C(_03645_),
    .Y(_04736_));
 OA22x2_ASAP7_75t_R _11597_ (.A1(_00202_),
    .A2(_03758_),
    .B1(_04736_),
    .B2(_03539_),
    .Y(_04737_));
 OR4x1_ASAP7_75t_R _11598_ (.A(_04195_),
    .B(_04726_),
    .C(_04730_),
    .D(_04737_),
    .Y(_04738_));
 OA22x2_ASAP7_75t_R _11599_ (.A1(_04698_),
    .A2(_04710_),
    .B1(_04722_),
    .B2(_04738_),
    .Y(_04739_));
 BUFx4f_ASAP7_75t_R _11600_ (.A(_04739_),
    .Y(_09977_));
 INVx3_ASAP7_75t_R _11601_ (.A(_09977_),
    .Y(_09979_));
 AND3x1_ASAP7_75t_R _11602_ (.A(net89),
    .B(net16),
    .C(_03600_),
    .Y(_04740_));
 OA21x2_ASAP7_75t_R _11603_ (.A1(_04251_),
    .A2(_04740_),
    .B(_04253_),
    .Y(_10158_));
 AND2x2_ASAP7_75t_R _11604_ (.A(_04033_),
    .B(_00238_),
    .Y(_04741_));
 AO21x1_ASAP7_75t_R _11605_ (.A1(_03950_),
    .A2(_00237_),
    .B(_04741_),
    .Y(_04742_));
 AO21x1_ASAP7_75t_R _11606_ (.A1(_03975_),
    .A2(_04742_),
    .B(_04130_),
    .Y(_04743_));
 AO22x1_ASAP7_75t_R _11607_ (.A1(_03986_),
    .A2(_00235_),
    .B1(_00236_),
    .B2(_04101_),
    .Y(_04744_));
 AO22x1_ASAP7_75t_R _11608_ (.A1(_03984_),
    .A2(_00235_),
    .B1(_04744_),
    .B2(_03992_),
    .Y(_04745_));
 AO21x1_ASAP7_75t_R _11609_ (.A1(_03381_),
    .A2(_04743_),
    .B(_04745_),
    .Y(_04746_));
 AND2x2_ASAP7_75t_R _11610_ (.A(_03933_),
    .B(_00242_),
    .Y(_04747_));
 AO21x1_ASAP7_75t_R _11611_ (.A1(_04125_),
    .A2(_00241_),
    .B(_04747_),
    .Y(_04748_));
 AND3x1_ASAP7_75t_R _11612_ (.A(_04137_),
    .B(_03943_),
    .C(_00240_),
    .Y(_04749_));
 AO21x1_ASAP7_75t_R _11613_ (.A1(_00239_),
    .A2(_03939_),
    .B(_04749_),
    .Y(_04750_));
 AO221x1_ASAP7_75t_R _11614_ (.A1(_04255_),
    .A2(_04748_),
    .B1(_04750_),
    .B2(_03938_),
    .C(_03947_),
    .Y(_04751_));
 AND2x2_ASAP7_75t_R _11615_ (.A(_04256_),
    .B(_00250_),
    .Y(_04752_));
 AO21x1_ASAP7_75t_R _11616_ (.A1(_04125_),
    .A2(_00249_),
    .B(_04752_),
    .Y(_04753_));
 AND3x1_ASAP7_75t_R _11617_ (.A(_03933_),
    .B(_03379_),
    .C(_00248_),
    .Y(_04754_));
 AO21x1_ASAP7_75t_R _11618_ (.A1(_00247_),
    .A2(_03939_),
    .B(_04754_),
    .Y(_04755_));
 AO221x2_ASAP7_75t_R _11619_ (.A1(_04255_),
    .A2(_04753_),
    .B1(_04755_),
    .B2(_03938_),
    .C(_03947_),
    .Y(_04756_));
 AND2x2_ASAP7_75t_R _11620_ (.A(_04043_),
    .B(_00245_),
    .Y(_04757_));
 AO21x1_ASAP7_75t_R _11621_ (.A1(_04520_),
    .A2(_00243_),
    .B(_04757_),
    .Y(_04758_));
 AO22x1_ASAP7_75t_R _11622_ (.A1(_00246_),
    .A2(_04090_),
    .B1(_04758_),
    .B2(_04663_),
    .Y(_04759_));
 AO21x1_ASAP7_75t_R _11623_ (.A1(_00244_),
    .A2(_03964_),
    .B(_03981_),
    .Y(_04760_));
 OA21x2_ASAP7_75t_R _11624_ (.A1(_04759_),
    .A2(_04760_),
    .B(_04280_),
    .Y(_04761_));
 AO32x2_ASAP7_75t_R _11625_ (.A1(_04514_),
    .A2(_04746_),
    .A3(_04751_),
    .B1(_04756_),
    .B2(_04761_),
    .Y(_04762_));
 BUFx10_ASAP7_75t_R _11626_ (.A(_04051_),
    .Y(_04763_));
 AND2x2_ASAP7_75t_R _11627_ (.A(_03942_),
    .B(_00258_),
    .Y(_04764_));
 AO21x1_ASAP7_75t_R _11628_ (.A1(_04671_),
    .A2(_00257_),
    .B(_04764_),
    .Y(_04765_));
 AND3x1_ASAP7_75t_R _11629_ (.A(_04666_),
    .B(_04559_),
    .C(_00256_),
    .Y(_04766_));
 AO21x1_ASAP7_75t_R _11630_ (.A1(_00255_),
    .A2(_04292_),
    .B(_04766_),
    .Y(_04767_));
 AO221x1_ASAP7_75t_R _11631_ (.A1(_04289_),
    .A2(_04765_),
    .B1(_04767_),
    .B2(_04295_),
    .C(_04298_),
    .Y(_04768_));
 AND2x2_ASAP7_75t_R _11632_ (.A(_03942_),
    .B(_00266_),
    .Y(_04769_));
 AO21x1_ASAP7_75t_R _11633_ (.A1(_04663_),
    .A2(_00265_),
    .B(_04769_),
    .Y(_04770_));
 AND3x1_ASAP7_75t_R _11634_ (.A(_04666_),
    .B(_04559_),
    .C(_00264_),
    .Y(_04771_));
 AO21x1_ASAP7_75t_R _11635_ (.A1(_00263_),
    .A2(_04292_),
    .B(_04771_),
    .Y(_04772_));
 AO221x1_ASAP7_75t_R _11636_ (.A1(_04289_),
    .A2(_04770_),
    .B1(_04772_),
    .B2(_04295_),
    .C(_04304_),
    .Y(_04773_));
 AND3x1_ASAP7_75t_R _11637_ (.A(_04763_),
    .B(_04768_),
    .C(_04773_),
    .Y(_04774_));
 AO22x1_ASAP7_75t_R _11638_ (.A1(_04529_),
    .A2(_00254_),
    .B1(_04068_),
    .B2(_00252_),
    .Y(_04775_));
 AO221x1_ASAP7_75t_R _11639_ (.A1(_04018_),
    .A2(_00262_),
    .B1(_04068_),
    .B2(_00260_),
    .C(_03996_),
    .Y(_04776_));
 OA211x2_ASAP7_75t_R _11640_ (.A1(_04156_),
    .A2(_04775_),
    .B(_04776_),
    .C(_04308_),
    .Y(_04777_));
 AND2x2_ASAP7_75t_R _11641_ (.A(_03974_),
    .B(_00261_),
    .Y(_04778_));
 AO21x1_ASAP7_75t_R _11642_ (.A1(_04276_),
    .A2(_00259_),
    .B(_04778_),
    .Y(_04779_));
 AND2x2_ASAP7_75t_R _11643_ (.A(_04105_),
    .B(_00253_),
    .Y(_04780_));
 AO221x1_ASAP7_75t_R _11644_ (.A1(_04111_),
    .A2(_04315_),
    .B1(_00251_),
    .B2(_04103_),
    .C(_04780_),
    .Y(_04781_));
 OA211x2_ASAP7_75t_R _11645_ (.A1(_03997_),
    .A2(_04779_),
    .B(_04781_),
    .C(_04265_),
    .Y(_04782_));
 OR3x1_ASAP7_75t_R _11646_ (.A(_04131_),
    .B(_04777_),
    .C(_04782_),
    .Y(_04783_));
 AO221x2_ASAP7_75t_R _11647_ (.A1(_03917_),
    .A2(_04762_),
    .B1(_04774_),
    .B2(_04783_),
    .C(_04055_),
    .Y(_04784_));
 NOR2x1_ASAP7_75t_R _11648_ (.A(_04254_),
    .B(_04784_),
    .Y(_04785_));
 AOI21x1_ASAP7_75t_R _11649_ (.A1(_04250_),
    .A2(_10158_),
    .B(_04785_),
    .Y(_04786_));
 XNOR2x1_ASAP7_75t_R _11650_ (.B(_04786_),
    .Y(_09985_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _11651_ (.A(_09985_),
    .Y(_09983_));
 AND3x1_ASAP7_75t_R _11652_ (.A(_03639_),
    .B(_03762_),
    .C(_00240_),
    .Y(_04787_));
 AO22x1_ASAP7_75t_R _11653_ (.A1(_00239_),
    .A2(_03878_),
    .B1(_04787_),
    .B2(_03677_),
    .Y(_04788_));
 OA222x2_ASAP7_75t_R _11654_ (.A1(_00241_),
    .A2(_03886_),
    .B1(_03585_),
    .B2(_00242_),
    .C1(_03765_),
    .C2(_03667_),
    .Y(_04789_));
 AO21x1_ASAP7_75t_R _11655_ (.A1(_03825_),
    .A2(_04788_),
    .B(_04789_),
    .Y(_04790_));
 AO21x2_ASAP7_75t_R _11656_ (.A1(_03791_),
    .A2(_04790_),
    .B(_03907_),
    .Y(_04791_));
 BUFx12_ASAP7_75t_R _11657_ (.A(_03825_),
    .Y(_04792_));
 AND3x1_ASAP7_75t_R _11658_ (.A(_03663_),
    .B(_03665_),
    .C(_00262_),
    .Y(_04793_));
 AO21x1_ASAP7_75t_R _11659_ (.A1(_00261_),
    .A2(_03711_),
    .B(_04793_),
    .Y(_04794_));
 AND3x1_ASAP7_75t_R _11660_ (.A(_03715_),
    .B(_03717_),
    .C(_00266_),
    .Y(_04795_));
 AO221x1_ASAP7_75t_R _11661_ (.A1(_00265_),
    .A2(_03805_),
    .B1(_03735_),
    .B2(_04478_),
    .C(_04795_),
    .Y(_04796_));
 OA21x2_ASAP7_75t_R _11662_ (.A1(_04602_),
    .A2(_04794_),
    .B(_04796_),
    .Y(_04797_));
 INVx2_ASAP7_75t_R _11663_ (.A(_00259_),
    .Y(_04798_));
 BUFx16f_ASAP7_75t_R _11664_ (.A(_04218_),
    .Y(_04799_));
 BUFx12f_ASAP7_75t_R _11665_ (.A(_04456_),
    .Y(_04800_));
 AND2x2_ASAP7_75t_R _11666_ (.A(_03610_),
    .B(_00264_),
    .Y(_04801_));
 AO21x1_ASAP7_75t_R _11667_ (.A1(_04609_),
    .A2(_00260_),
    .B(_04801_),
    .Y(_04802_));
 AOI22x1_ASAP7_75t_R _11668_ (.A1(_00263_),
    .A2(_04800_),
    .B1(_04802_),
    .B2(_04597_),
    .Y(_04803_));
 BUFx10_ASAP7_75t_R _11669_ (.A(_03607_),
    .Y(_04804_));
 OA211x2_ASAP7_75t_R _11670_ (.A1(_03481_),
    .A2(_04803_),
    .B(_04804_),
    .C(_03861_),
    .Y(_04805_));
 BUFx12_ASAP7_75t_R _11671_ (.A(_04163_),
    .Y(_04806_));
 OAI22x1_ASAP7_75t_R _11672_ (.A1(_04798_),
    .A2(_04799_),
    .B1(_04805_),
    .B2(_04806_),
    .Y(_04807_));
 OA211x2_ASAP7_75t_R _11673_ (.A1(_04792_),
    .A2(_04797_),
    .B(_04807_),
    .C(_03850_),
    .Y(_04808_));
 NAND2x2_ASAP7_75t_R _11674_ (.A(_04791_),
    .B(_04808_),
    .Y(_04809_));
 AND3x1_ASAP7_75t_R _11675_ (.A(_00256_),
    .B(_04591_),
    .C(_04727_),
    .Y(_04810_));
 BUFx12_ASAP7_75t_R _11676_ (.A(_03628_),
    .Y(_04811_));
 INVx2_ASAP7_75t_R _11677_ (.A(_00253_),
    .Y(_04812_));
 INVx1_ASAP7_75t_R _11678_ (.A(_00252_),
    .Y(_04813_));
 NAND2x1_ASAP7_75t_R _11679_ (.A(_03619_),
    .B(_00254_),
    .Y(_04814_));
 OA211x2_ASAP7_75t_R _11680_ (.A1(_03636_),
    .A2(_04813_),
    .B(_04814_),
    .C(_03614_),
    .Y(_04815_));
 AOI21x1_ASAP7_75t_R _11681_ (.A1(_04812_),
    .A2(_04442_),
    .B(_04815_),
    .Y(_04816_));
 OA211x2_ASAP7_75t_R _11682_ (.A1(_04811_),
    .A2(_04816_),
    .B(_03771_),
    .C(_03860_),
    .Y(_04817_));
 OA22x2_ASAP7_75t_R _11683_ (.A1(_00251_),
    .A2(_03759_),
    .B1(_04817_),
    .B2(_03785_),
    .Y(_04818_));
 AND3x1_ASAP7_75t_R _11684_ (.A(_03395_),
    .B(_03672_),
    .C(_00258_),
    .Y(_04819_));
 AO21x1_ASAP7_75t_R _11685_ (.A1(_00257_),
    .A2(_03671_),
    .B(_04819_),
    .Y(_04820_));
 OA21x2_ASAP7_75t_R _11686_ (.A1(_03606_),
    .A2(_03681_),
    .B(_04820_),
    .Y(_04821_));
 AND3x1_ASAP7_75t_R _11687_ (.A(_00255_),
    .B(_03646_),
    .C(_03648_),
    .Y(_04822_));
 OA211x2_ASAP7_75t_R _11688_ (.A1(_04821_),
    .A2(_04822_),
    .B(_04244_),
    .C(_03653_),
    .Y(_04823_));
 OR4x2_ASAP7_75t_R _11689_ (.A(_03723_),
    .B(_04810_),
    .C(_04818_),
    .D(_04823_),
    .Y(_04824_));
 AND4x1_ASAP7_75t_R _11690_ (.A(_00238_),
    .B(_03677_),
    .C(_03678_),
    .D(_04587_),
    .Y(_04825_));
 AO21x1_ASAP7_75t_R _11691_ (.A1(_00236_),
    .A2(_04583_),
    .B(_04825_),
    .Y(_04826_));
 OA21x2_ASAP7_75t_R _11692_ (.A1(_00237_),
    .A2(_03866_),
    .B(_04627_),
    .Y(_04827_));
 OA22x2_ASAP7_75t_R _11693_ (.A1(_03587_),
    .A2(_04826_),
    .B1(_04827_),
    .B2(_04165_),
    .Y(_04828_));
 AND2x2_ASAP7_75t_R _11694_ (.A(_03624_),
    .B(_00250_),
    .Y(_04829_));
 AO21x1_ASAP7_75t_R _11695_ (.A1(_03629_),
    .A2(_00249_),
    .B(_04829_),
    .Y(_04830_));
 BUFx12f_ASAP7_75t_R _11696_ (.A(_03744_),
    .Y(_04831_));
 AO22x2_ASAP7_75t_R _11697_ (.A1(_03510_),
    .A2(_03490_),
    .B1(_03394_),
    .B2(_03613_),
    .Y(_04832_));
 OA222x2_ASAP7_75t_R _11698_ (.A1(_03480_),
    .A2(_04831_),
    .B1(_00246_),
    .B2(_03710_),
    .C1(_04832_),
    .C2(_00245_),
    .Y(_04833_));
 AO21x1_ASAP7_75t_R _11699_ (.A1(_03670_),
    .A2(_04830_),
    .B(_04833_),
    .Y(_04834_));
 OR3x1_ASAP7_75t_R _11700_ (.A(_00245_),
    .B(_03657_),
    .C(_04204_),
    .Y(_04835_));
 OR4x2_ASAP7_75t_R _11701_ (.A(_03511_),
    .B(_03512_),
    .C(_03513_),
    .D(_03514_),
    .Y(_04836_));
 OR4x1_ASAP7_75t_R _11702_ (.A(_00249_),
    .B(_04836_),
    .C(_03642_),
    .D(_03728_),
    .Y(_04837_));
 AND3x1_ASAP7_75t_R _11703_ (.A(_04834_),
    .B(_04835_),
    .C(_04837_),
    .Y(_04838_));
 AND2x6_ASAP7_75t_R _11704_ (.A(_03898_),
    .B(_03698_),
    .Y(_04839_));
 INVx1_ASAP7_75t_R _11705_ (.A(_00243_),
    .Y(_04840_));
 AND2x2_ASAP7_75t_R _11706_ (.A(_04610_),
    .B(_00248_),
    .Y(_04841_));
 AO21x1_ASAP7_75t_R _11707_ (.A1(_04609_),
    .A2(_00244_),
    .B(_04841_),
    .Y(_04842_));
 AOI22x1_ASAP7_75t_R _11708_ (.A1(_00247_),
    .A2(_04800_),
    .B1(_04842_),
    .B2(_03853_),
    .Y(_04843_));
 OA211x2_ASAP7_75t_R _11709_ (.A1(_03481_),
    .A2(_04843_),
    .B(_03802_),
    .C(_03836_),
    .Y(_04844_));
 OAI22x1_ASAP7_75t_R _11710_ (.A1(_04840_),
    .A2(_04799_),
    .B1(_04844_),
    .B2(_04164_),
    .Y(_04845_));
 OA211x2_ASAP7_75t_R _11711_ (.A1(_04583_),
    .A2(_04838_),
    .B(_04839_),
    .C(_04845_),
    .Y(_04846_));
 AOI211x1_ASAP7_75t_R _11712_ (.A1(_04791_),
    .A2(_04824_),
    .B(_04828_),
    .C(_04846_),
    .Y(_04847_));
 AND2x2_ASAP7_75t_R _11713_ (.A(_04809_),
    .B(_04847_),
    .Y(_09984_));
 BUFx3_ASAP7_75t_R _11714_ (.A(_04165_),
    .Y(_04848_));
 BUFx4f_ASAP7_75t_R _11715_ (.A(_04848_),
    .Y(_04849_));
 AO21x1_ASAP7_75t_R _11716_ (.A1(_04124_),
    .A2(_04849_),
    .B(_04251_),
    .Y(_04850_));
 AND2x2_ASAP7_75t_R _11717_ (.A(_04253_),
    .B(_04850_),
    .Y(_10156_));
 AND2x2_ASAP7_75t_R _11718_ (.A(_04033_),
    .B(_00271_),
    .Y(_04851_));
 AO21x1_ASAP7_75t_R _11719_ (.A1(_03976_),
    .A2(_00270_),
    .B(_04851_),
    .Y(_04852_));
 AO21x1_ASAP7_75t_R _11720_ (.A1(_03975_),
    .A2(_04852_),
    .B(_03981_),
    .Y(_04853_));
 AO22x1_ASAP7_75t_R _11721_ (.A1(_03986_),
    .A2(_00268_),
    .B1(_00269_),
    .B2(_03989_),
    .Y(_04854_));
 AO22x1_ASAP7_75t_R _11722_ (.A1(_03984_),
    .A2(_00268_),
    .B1(_04854_),
    .B2(_03992_),
    .Y(_04855_));
 AO21x1_ASAP7_75t_R _11723_ (.A1(_03381_),
    .A2(_04853_),
    .B(_04855_),
    .Y(_04856_));
 AND2x2_ASAP7_75t_R _11724_ (.A(_04256_),
    .B(_00275_),
    .Y(_04857_));
 AO21x1_ASAP7_75t_R _11725_ (.A1(_04125_),
    .A2(_00274_),
    .B(_04857_),
    .Y(_04858_));
 AND3x1_ASAP7_75t_R _11726_ (.A(_04137_),
    .B(_03379_),
    .C(_00273_),
    .Y(_04859_));
 AO21x1_ASAP7_75t_R _11727_ (.A1(_00272_),
    .A2(_03939_),
    .B(_04859_),
    .Y(_04860_));
 AO221x1_ASAP7_75t_R _11728_ (.A1(_04255_),
    .A2(_04858_),
    .B1(_04860_),
    .B2(_03938_),
    .C(_03947_),
    .Y(_04861_));
 AND2x2_ASAP7_75t_R _11729_ (.A(_04256_),
    .B(_00283_),
    .Y(_04862_));
 AO21x1_ASAP7_75t_R _11730_ (.A1(_04125_),
    .A2(_00282_),
    .B(_04862_),
    .Y(_04863_));
 AND3x1_ASAP7_75t_R _11731_ (.A(_03933_),
    .B(_03379_),
    .C(_00281_),
    .Y(_04864_));
 AO21x1_ASAP7_75t_R _11732_ (.A1(_00280_),
    .A2(_03939_),
    .B(_04864_),
    .Y(_04865_));
 AO221x1_ASAP7_75t_R _11733_ (.A1(_04255_),
    .A2(_04863_),
    .B1(_04865_),
    .B2(_03938_),
    .C(_03947_),
    .Y(_04866_));
 AND2x2_ASAP7_75t_R _11734_ (.A(_04043_),
    .B(_00278_),
    .Y(_04867_));
 AO21x1_ASAP7_75t_R _11735_ (.A1(_03991_),
    .A2(_00276_),
    .B(_04867_),
    .Y(_04868_));
 AO22x1_ASAP7_75t_R _11736_ (.A1(_00279_),
    .A2(_04090_),
    .B1(_04868_),
    .B2(_04663_),
    .Y(_04869_));
 AO21x1_ASAP7_75t_R _11737_ (.A1(_00277_),
    .A2(_03964_),
    .B(_03981_),
    .Y(_04870_));
 OA21x2_ASAP7_75t_R _11738_ (.A1(_04869_),
    .A2(_04870_),
    .B(_04280_),
    .Y(_04871_));
 AO32x1_ASAP7_75t_R _11739_ (.A1(_04514_),
    .A2(_04856_),
    .A3(_04861_),
    .B1(_04866_),
    .B2(_04871_),
    .Y(_04872_));
 AND2x2_ASAP7_75t_R _11740_ (.A(_03942_),
    .B(_00291_),
    .Y(_04873_));
 AO21x1_ASAP7_75t_R _11741_ (.A1(_04663_),
    .A2(_00290_),
    .B(_04873_),
    .Y(_04874_));
 AND3x1_ASAP7_75t_R _11742_ (.A(_04666_),
    .B(_03943_),
    .C(_00289_),
    .Y(_04875_));
 AO21x1_ASAP7_75t_R _11743_ (.A1(_00288_),
    .A2(_04292_),
    .B(_04875_),
    .Y(_04876_));
 AO221x1_ASAP7_75t_R _11744_ (.A1(_04289_),
    .A2(_04874_),
    .B1(_04876_),
    .B2(_04295_),
    .C(_04298_),
    .Y(_04877_));
 AND2x2_ASAP7_75t_R _11745_ (.A(_04137_),
    .B(_00299_),
    .Y(_04878_));
 AO21x2_ASAP7_75t_R _11746_ (.A1(_04663_),
    .A2(_00298_),
    .B(_04878_),
    .Y(_04879_));
 AND3x1_ASAP7_75t_R _11747_ (.A(_04666_),
    .B(_03943_),
    .C(_00297_),
    .Y(_04880_));
 AO21x1_ASAP7_75t_R _11748_ (.A1(_00296_),
    .A2(_04292_),
    .B(_04880_),
    .Y(_04881_));
 AO221x1_ASAP7_75t_R _11749_ (.A1(_04289_),
    .A2(_04879_),
    .B1(_04881_),
    .B2(_04295_),
    .C(_04304_),
    .Y(_04882_));
 AND3x1_ASAP7_75t_R _11750_ (.A(_04051_),
    .B(_04877_),
    .C(_04882_),
    .Y(_04883_));
 AO221x1_ASAP7_75t_R _11751_ (.A1(_04270_),
    .A2(_00295_),
    .B1(_04632_),
    .B2(_00293_),
    .C(_04097_),
    .Y(_04884_));
 AO221x1_ASAP7_75t_R _11752_ (.A1(_04270_),
    .A2(_00287_),
    .B1(_04632_),
    .B2(_00285_),
    .C(_03920_),
    .Y(_04885_));
 AO21x1_ASAP7_75t_R _11753_ (.A1(_04884_),
    .A2(_04885_),
    .B(_04080_),
    .Y(_04886_));
 INVx1_ASAP7_75t_R _11754_ (.A(_00286_),
    .Y(_04887_));
 NAND2x1_ASAP7_75t_R _11755_ (.A(_04276_),
    .B(_00284_),
    .Y(_04888_));
 OA211x2_ASAP7_75t_R _11756_ (.A1(_04114_),
    .A2(_04887_),
    .B(_04097_),
    .C(_04888_),
    .Y(_04889_));
 INVx1_ASAP7_75t_R _11757_ (.A(_00294_),
    .Y(_04890_));
 NAND2x1_ASAP7_75t_R _11758_ (.A(_04276_),
    .B(_00292_),
    .Y(_04891_));
 OA211x2_ASAP7_75t_R _11759_ (.A1(_04114_),
    .A2(_04890_),
    .B(_03920_),
    .C(_04891_),
    .Y(_04892_));
 OAI21x1_ASAP7_75t_R _11760_ (.A1(_04889_),
    .A2(_04892_),
    .B(_04089_),
    .Y(_04893_));
 AO21x1_ASAP7_75t_R _11761_ (.A1(_04886_),
    .A2(_04893_),
    .B(_04131_),
    .Y(_04894_));
 AO221x2_ASAP7_75t_R _11762_ (.A1(_03917_),
    .A2(_04872_),
    .B1(_04883_),
    .B2(_04894_),
    .C(_04055_),
    .Y(_04895_));
 NOR2x1_ASAP7_75t_R _11763_ (.A(_04254_),
    .B(_04895_),
    .Y(_04896_));
 AOI21x1_ASAP7_75t_R _11764_ (.A1(_04250_),
    .A2(_10156_),
    .B(_04896_),
    .Y(_04897_));
 XNOR2x1_ASAP7_75t_R _11765_ (.B(_04897_),
    .Y(_09988_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _11766_ (.A(_09988_),
    .Y(_09990_));
 INVx1_ASAP7_75t_R _11767_ (.A(_00295_),
    .Y(_04898_));
 OR3x1_ASAP7_75t_R _11768_ (.A(_03839_),
    .B(_03840_),
    .C(_04898_),
    .Y(_04899_));
 INVx1_ASAP7_75t_R _11769_ (.A(_00298_),
    .Y(_04900_));
 AO21x1_ASAP7_75t_R _11770_ (.A1(_03639_),
    .A2(_03717_),
    .B(_04900_),
    .Y(_04901_));
 INVx1_ASAP7_75t_R _11771_ (.A(_00299_),
    .Y(_04902_));
 OR3x1_ASAP7_75t_R _11772_ (.A(_03480_),
    .B(_03629_),
    .C(_04902_),
    .Y(_04903_));
 AO22x2_ASAP7_75t_R _11773_ (.A1(_03836_),
    .A2(_03735_),
    .B1(_04901_),
    .B2(_04903_),
    .Y(_04904_));
 AO21x1_ASAP7_75t_R _11774_ (.A1(_00294_),
    .A2(_03830_),
    .B(_03775_),
    .Y(_04905_));
 NAND2x1_ASAP7_75t_R _11775_ (.A(_03705_),
    .B(_04905_),
    .Y(_04906_));
 OA211x2_ASAP7_75t_R _11776_ (.A1(_04602_),
    .A2(_04899_),
    .B(_04904_),
    .C(_04906_),
    .Y(_04907_));
 INVx1_ASAP7_75t_R _11777_ (.A(_00292_),
    .Y(_04908_));
 AND2x2_ASAP7_75t_R _11778_ (.A(_04610_),
    .B(_00297_),
    .Y(_04909_));
 AO21x1_ASAP7_75t_R _11779_ (.A1(_04609_),
    .A2(_00293_),
    .B(_04909_),
    .Y(_04910_));
 AOI22x1_ASAP7_75t_R _11780_ (.A1(_00296_),
    .A2(_04576_),
    .B1(_04910_),
    .B2(_03665_),
    .Y(_04911_));
 OA211x2_ASAP7_75t_R _11781_ (.A1(_03839_),
    .A2(_04911_),
    .B(_03802_),
    .C(_03836_),
    .Y(_04912_));
 OA22x2_ASAP7_75t_R _11782_ (.A1(_04908_),
    .A2(_04575_),
    .B1(_04912_),
    .B2(_04164_),
    .Y(_04913_));
 OR3x4_ASAP7_75t_R _11783_ (.A(_04468_),
    .B(_04907_),
    .C(_04913_),
    .Y(_04914_));
 BUFx6f_ASAP7_75t_R _11784_ (.A(_03701_),
    .Y(_04915_));
 BUFx12_ASAP7_75t_R _11785_ (.A(_03623_),
    .Y(_04916_));
 AND3x1_ASAP7_75t_R _11786_ (.A(_04916_),
    .B(_04584_),
    .C(_00287_),
    .Y(_04917_));
 AO21x1_ASAP7_75t_R _11787_ (.A1(_00286_),
    .A2(_03891_),
    .B(_04917_),
    .Y(_04918_));
 AO32x1_ASAP7_75t_R _11788_ (.A1(_03655_),
    .A2(_04587_),
    .A3(_04918_),
    .B1(_03703_),
    .B2(_00284_),
    .Y(_04919_));
 BUFx10_ASAP7_75t_R _11789_ (.A(_03653_),
    .Y(_04920_));
 BUFx12f_ASAP7_75t_R _11790_ (.A(_03881_),
    .Y(_04921_));
 AND2x2_ASAP7_75t_R _11791_ (.A(_00290_),
    .B(_03710_),
    .Y(_04922_));
 AO221x1_ASAP7_75t_R _11792_ (.A1(_00291_),
    .A2(_04921_),
    .B1(_04804_),
    .B2(_04478_),
    .C(_04922_),
    .Y(_04923_));
 OA33x2_ASAP7_75t_R _11793_ (.A1(_03816_),
    .A2(_00289_),
    .A3(_03805_),
    .B1(_04344_),
    .B2(_03667_),
    .B3(_00288_),
    .Y(_04924_));
 AND4x1_ASAP7_75t_R _11794_ (.A(_03655_),
    .B(_04920_),
    .C(_04923_),
    .D(_04924_),
    .Y(_04925_));
 AND3x1_ASAP7_75t_R _11795_ (.A(_00285_),
    .B(_04591_),
    .C(_03776_),
    .Y(_04926_));
 AO21x1_ASAP7_75t_R _11796_ (.A1(_04915_),
    .A2(_04926_),
    .B(_04499_),
    .Y(_04927_));
 AOI211x1_ASAP7_75t_R _11797_ (.A1(_04915_),
    .A2(_04919_),
    .B(_04925_),
    .C(_04927_),
    .Y(_04928_));
 BUFx10_ASAP7_75t_R _11798_ (.A(_03714_),
    .Y(_04929_));
 BUFx12f_ASAP7_75t_R _11799_ (.A(_03665_),
    .Y(_04930_));
 AND3x1_ASAP7_75t_R _11800_ (.A(_03815_),
    .B(_04930_),
    .C(_00275_),
    .Y(_04931_));
 AO21x1_ASAP7_75t_R _11801_ (.A1(_00274_),
    .A2(_04929_),
    .B(_04931_),
    .Y(_04932_));
 INVx2_ASAP7_75t_R _11802_ (.A(_00276_),
    .Y(_04933_));
 BUFx16f_ASAP7_75t_R _11803_ (.A(_04575_),
    .Y(_04934_));
 BUFx10_ASAP7_75t_R _11804_ (.A(_03839_),
    .Y(_04935_));
 BUFx16f_ASAP7_75t_R _11805_ (.A(_04576_),
    .Y(_04936_));
 BUFx12f_ASAP7_75t_R _11806_ (.A(_04457_),
    .Y(_04937_));
 BUFx10_ASAP7_75t_R _11807_ (.A(_03609_),
    .Y(_04938_));
 AND2x2_ASAP7_75t_R _11808_ (.A(_04938_),
    .B(_00281_),
    .Y(_04939_));
 AO21x1_ASAP7_75t_R _11809_ (.A1(_04937_),
    .A2(_00277_),
    .B(_04939_),
    .Y(_04940_));
 AOI22x1_ASAP7_75t_R _11810_ (.A1(_00280_),
    .A2(_04936_),
    .B1(_04940_),
    .B2(_03845_),
    .Y(_04941_));
 OA211x2_ASAP7_75t_R _11811_ (.A1(_04935_),
    .A2(_04941_),
    .B(_03776_),
    .C(_03829_),
    .Y(_04942_));
 OAI22x1_ASAP7_75t_R _11812_ (.A1(_04933_),
    .A2(_04934_),
    .B1(_04942_),
    .B2(_03786_),
    .Y(_04943_));
 AO21x1_ASAP7_75t_R _11813_ (.A1(_03860_),
    .A2(_03707_),
    .B(_03881_),
    .Y(_04944_));
 NAND2x2_ASAP7_75t_R _11814_ (.A(_03614_),
    .B(_03609_),
    .Y(_04945_));
 OA22x2_ASAP7_75t_R _11815_ (.A1(_00278_),
    .A2(_03690_),
    .B1(_04945_),
    .B2(_00283_),
    .Y(_04946_));
 OR3x1_ASAP7_75t_R _11816_ (.A(_03414_),
    .B(_03631_),
    .C(_03608_),
    .Y(_04947_));
 BUFx10_ASAP7_75t_R _11817_ (.A(_04947_),
    .Y(_04948_));
 OR2x2_ASAP7_75t_R _11818_ (.A(_03709_),
    .B(_04948_),
    .Y(_04949_));
 OA22x2_ASAP7_75t_R _11819_ (.A1(_04592_),
    .A2(_04946_),
    .B1(_04949_),
    .B2(_00279_),
    .Y(_04950_));
 OA211x2_ASAP7_75t_R _11820_ (.A1(_00282_),
    .A2(_04944_),
    .B(_04950_),
    .C(_03868_),
    .Y(_04951_));
 BUFx12_ASAP7_75t_R _11821_ (.A(_03620_),
    .Y(_04952_));
 OR2x2_ASAP7_75t_R _11822_ (.A(_00269_),
    .B(_04952_),
    .Y(_04953_));
 AND3x1_ASAP7_75t_R _11823_ (.A(_03623_),
    .B(_04435_),
    .C(_00271_),
    .Y(_04954_));
 AO21x1_ASAP7_75t_R _11824_ (.A1(_00270_),
    .A2(_03890_),
    .B(_04954_),
    .Y(_04955_));
 OA211x2_ASAP7_75t_R _11825_ (.A1(_04804_),
    .A2(_04955_),
    .B(_04192_),
    .C(_04478_),
    .Y(_04956_));
 AND3x1_ASAP7_75t_R _11826_ (.A(_04455_),
    .B(_04584_),
    .C(_00273_),
    .Y(_04957_));
 AO21x1_ASAP7_75t_R _11827_ (.A1(_00272_),
    .A2(_03782_),
    .B(_04957_),
    .Y(_04958_));
 BUFx6f_ASAP7_75t_R _11828_ (.A(_04194_),
    .Y(_04959_));
 AO221x1_ASAP7_75t_R _11829_ (.A1(_04953_),
    .A2(_04956_),
    .B1(_04958_),
    .B2(_04727_),
    .C(_04959_),
    .Y(_04960_));
 AOI221x1_ASAP7_75t_R _11830_ (.A1(_04440_),
    .A2(_04932_),
    .B1(_04943_),
    .B2(_04951_),
    .C(_04960_),
    .Y(_04961_));
 AO21x1_ASAP7_75t_R _11831_ (.A1(_04914_),
    .A2(_04928_),
    .B(_04961_),
    .Y(_04962_));
 BUFx4f_ASAP7_75t_R _11832_ (.A(_04962_),
    .Y(_09987_));
 INVx3_ASAP7_75t_R _11833_ (.A(_09987_),
    .Y(_09989_));
 AO21x1_ASAP7_75t_R _11834_ (.A1(_04157_),
    .A2(_04849_),
    .B(_04251_),
    .Y(_04963_));
 AND2x2_ASAP7_75t_R _11835_ (.A(_04253_),
    .B(_04963_),
    .Y(_10154_));
 AND2x2_ASAP7_75t_R _11836_ (.A(_04256_),
    .B(_00304_),
    .Y(_04964_));
 AO21x1_ASAP7_75t_R _11837_ (.A1(_04125_),
    .A2(_00303_),
    .B(_04964_),
    .Y(_04965_));
 AO21x1_ASAP7_75t_R _11838_ (.A1(_03927_),
    .A2(_04965_),
    .B(_04130_),
    .Y(_04966_));
 AO22x1_ASAP7_75t_R _11839_ (.A1(_03950_),
    .A2(_00301_),
    .B1(_00302_),
    .B2(_04101_),
    .Y(_04967_));
 AO22x1_ASAP7_75t_R _11840_ (.A1(_04071_),
    .A2(_00301_),
    .B1(_04967_),
    .B2(_04521_),
    .Y(_04968_));
 AO21x1_ASAP7_75t_R _11841_ (.A1(_03381_),
    .A2(_04966_),
    .B(_04968_),
    .Y(_04969_));
 AND2x2_ASAP7_75t_R _11842_ (.A(_04015_),
    .B(_00308_),
    .Y(_04970_));
 AO21x1_ASAP7_75t_R _11843_ (.A1(_04556_),
    .A2(_00307_),
    .B(_04970_),
    .Y(_04971_));
 AND3x1_ASAP7_75t_R _11844_ (.A(_04015_),
    .B(_04559_),
    .C(_00306_),
    .Y(_04972_));
 AO21x1_ASAP7_75t_R _11845_ (.A1(_00305_),
    .A2(_04535_),
    .B(_04972_),
    .Y(_04973_));
 AO221x1_ASAP7_75t_R _11846_ (.A1(_04502_),
    .A2(_04971_),
    .B1(_04973_),
    .B2(_04540_),
    .C(_04094_),
    .Y(_04974_));
 AND2x2_ASAP7_75t_R _11847_ (.A(_04666_),
    .B(_00316_),
    .Y(_04975_));
 AO21x1_ASAP7_75t_R _11848_ (.A1(_04671_),
    .A2(_00315_),
    .B(_04975_),
    .Y(_04976_));
 AND3x1_ASAP7_75t_R _11849_ (.A(_04015_),
    .B(_04559_),
    .C(_00314_),
    .Y(_04977_));
 AO21x1_ASAP7_75t_R _11850_ (.A1(_00313_),
    .A2(_04535_),
    .B(_04977_),
    .Y(_04978_));
 AO221x1_ASAP7_75t_R _11851_ (.A1(_04502_),
    .A2(_04976_),
    .B1(_04978_),
    .B2(_04540_),
    .C(_04094_),
    .Y(_04979_));
 AND2x2_ASAP7_75t_R _11852_ (.A(_03925_),
    .B(_00311_),
    .Y(_04980_));
 AO21x1_ASAP7_75t_R _11853_ (.A1(_04113_),
    .A2(_00309_),
    .B(_04980_),
    .Y(_04981_));
 AO22x1_ASAP7_75t_R _11854_ (.A1(_00312_),
    .A2(_04090_),
    .B1(_04981_),
    .B2(_04647_),
    .Y(_04982_));
 BUFx10_ASAP7_75t_R _11855_ (.A(_04266_),
    .Y(_04983_));
 AO21x1_ASAP7_75t_R _11856_ (.A1(_00310_),
    .A2(_04983_),
    .B(_04130_),
    .Y(_04984_));
 OA21x2_ASAP7_75t_R _11857_ (.A1(_04982_),
    .A2(_04984_),
    .B(_04280_),
    .Y(_04985_));
 AO32x1_ASAP7_75t_R _11858_ (.A1(_04099_),
    .A2(_04969_),
    .A3(_04974_),
    .B1(_04979_),
    .B2(_04985_),
    .Y(_04986_));
 BUFx12_ASAP7_75t_R _11859_ (.A(_04269_),
    .Y(_04987_));
 BUFx6f_ASAP7_75t_R _11860_ (.A(_04987_),
    .Y(_04988_));
 AND2x2_ASAP7_75t_R _11861_ (.A(_04537_),
    .B(_00324_),
    .Y(_04989_));
 AO21x1_ASAP7_75t_R _11862_ (.A1(_04647_),
    .A2(_00323_),
    .B(_04989_),
    .Y(_04990_));
 BUFx10_ASAP7_75t_R _11863_ (.A(_04001_),
    .Y(_04991_));
 BUFx10_ASAP7_75t_R _11864_ (.A(_04536_),
    .Y(_04992_));
 AND3x1_ASAP7_75t_R _11865_ (.A(_04992_),
    .B(_03971_),
    .C(_00322_),
    .Y(_04993_));
 AO21x1_ASAP7_75t_R _11866_ (.A1(_00321_),
    .A2(_04991_),
    .B(_04993_),
    .Y(_04994_));
 BUFx6f_ASAP7_75t_R _11867_ (.A(_03937_),
    .Y(_04995_));
 BUFx10_ASAP7_75t_R _11868_ (.A(_04995_),
    .Y(_04996_));
 AO221x1_ASAP7_75t_R _11869_ (.A1(_04988_),
    .A2(_04990_),
    .B1(_04994_),
    .B2(_04996_),
    .C(_04298_),
    .Y(_04997_));
 AND2x2_ASAP7_75t_R _11870_ (.A(_04537_),
    .B(_00332_),
    .Y(_04998_));
 AO21x1_ASAP7_75t_R _11871_ (.A1(_04647_),
    .A2(_00331_),
    .B(_04998_),
    .Y(_04999_));
 AND3x1_ASAP7_75t_R _11872_ (.A(_04537_),
    .B(_03971_),
    .C(_00330_),
    .Y(_05000_));
 AO21x1_ASAP7_75t_R _11873_ (.A1(_00329_),
    .A2(_04991_),
    .B(_05000_),
    .Y(_05001_));
 AO221x1_ASAP7_75t_R _11874_ (.A1(_04530_),
    .A2(_04999_),
    .B1(_05001_),
    .B2(_04996_),
    .C(_04304_),
    .Y(_05002_));
 AND3x1_ASAP7_75t_R _11875_ (.A(_04763_),
    .B(_04997_),
    .C(_05002_),
    .Y(_05003_));
 AO221x1_ASAP7_75t_R _11876_ (.A1(_04987_),
    .A2(_00328_),
    .B1(_04632_),
    .B2(_00326_),
    .C(_04097_),
    .Y(_05004_));
 AO221x1_ASAP7_75t_R _11877_ (.A1(_04987_),
    .A2(_00320_),
    .B1(_04068_),
    .B2(_00318_),
    .C(_04279_),
    .Y(_05005_));
 AND3x1_ASAP7_75t_R _11878_ (.A(_04308_),
    .B(_05004_),
    .C(_05005_),
    .Y(_05006_));
 AND2x2_ASAP7_75t_R _11879_ (.A(_04018_),
    .B(_00327_),
    .Y(_05007_));
 AO21x1_ASAP7_75t_R _11880_ (.A1(_04521_),
    .A2(_00325_),
    .B(_05007_),
    .Y(_05008_));
 AND2x2_ASAP7_75t_R _11881_ (.A(_04269_),
    .B(_00319_),
    .Y(_05009_));
 AO221x1_ASAP7_75t_R _11882_ (.A1(_04111_),
    .A2(_04315_),
    .B1(_00317_),
    .B2(_04276_),
    .C(_05009_),
    .Y(_05010_));
 OA211x2_ASAP7_75t_R _11883_ (.A1(_04098_),
    .A2(_05008_),
    .B(_05010_),
    .C(_04136_),
    .Y(_05011_));
 OR3x1_ASAP7_75t_R _11884_ (.A(_04131_),
    .B(_05006_),
    .C(_05011_),
    .Y(_05012_));
 AO221x2_ASAP7_75t_R _11885_ (.A1(_03917_),
    .A2(_04986_),
    .B1(_05003_),
    .B2(_05012_),
    .C(_04055_),
    .Y(_05013_));
 BUFx3_ASAP7_75t_R _11886_ (.A(_05013_),
    .Y(_05014_));
 NOR2x1_ASAP7_75t_R _11887_ (.A(_04254_),
    .B(_05014_),
    .Y(_05015_));
 AOI21x1_ASAP7_75t_R _11888_ (.A1(_04250_),
    .A2(_10154_),
    .B(_05015_),
    .Y(_05016_));
 XNOR2x1_ASAP7_75t_R _11889_ (.B(_05016_),
    .Y(_09993_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _11890_ (.A(_09993_),
    .Y(_09995_));
 INVx1_ASAP7_75t_R _11891_ (.A(_00325_),
    .Y(_05017_));
 AND2x2_ASAP7_75t_R _11892_ (.A(_03685_),
    .B(_00330_),
    .Y(_05018_));
 AO21x1_ASAP7_75t_R _11893_ (.A1(_03683_),
    .A2(_00326_),
    .B(_05018_),
    .Y(_05019_));
 AOI22x1_ASAP7_75t_R _11894_ (.A1(_00329_),
    .A2(_04210_),
    .B1(_05019_),
    .B2(_03664_),
    .Y(_05020_));
 OA211x2_ASAP7_75t_R _11895_ (.A1(_03419_),
    .A2(_05020_),
    .B(_04212_),
    .C(_03736_),
    .Y(_05021_));
 OA22x2_ASAP7_75t_R _11896_ (.A1(_05017_),
    .A2(_04218_),
    .B1(_05021_),
    .B2(_04214_),
    .Y(_05022_));
 AND3x1_ASAP7_75t_R _11897_ (.A(_03374_),
    .B(_03672_),
    .C(_00328_),
    .Y(_05023_));
 AO21x1_ASAP7_75t_R _11898_ (.A1(_00327_),
    .A2(_03612_),
    .B(_05023_),
    .Y(_05024_));
 OR3x1_ASAP7_75t_R _11899_ (.A(_03606_),
    .B(_03670_),
    .C(_05024_),
    .Y(_05025_));
 AND2x2_ASAP7_75t_R _11900_ (.A(_00331_),
    .B(_03612_),
    .Y(_05026_));
 AO221x1_ASAP7_75t_R _11901_ (.A1(_00332_),
    .A2(_03881_),
    .B1(_03661_),
    .B2(_03860_),
    .C(_05026_),
    .Y(_05027_));
 AOI21x1_ASAP7_75t_R _11902_ (.A1(_05025_),
    .A2(_05027_),
    .B(_04454_),
    .Y(_05028_));
 OR3x1_ASAP7_75t_R _11903_ (.A(_03740_),
    .B(_05022_),
    .C(_05028_),
    .Y(_05029_));
 AND3x1_ASAP7_75t_R _11904_ (.A(_03549_),
    .B(_03624_),
    .C(_00320_),
    .Y(_05030_));
 AO21x1_ASAP7_75t_R _11905_ (.A1(_00319_),
    .A2(_03890_),
    .B(_05030_),
    .Y(_05031_));
 AO32x1_ASAP7_75t_R _11906_ (.A1(_04244_),
    .A2(_03731_),
    .A3(_05031_),
    .B1(_03702_),
    .B2(_00317_),
    .Y(_05032_));
 AND2x2_ASAP7_75t_R _11907_ (.A(_00323_),
    .B(_03709_),
    .Y(_05033_));
 AO221x1_ASAP7_75t_R _11908_ (.A1(_00324_),
    .A2(_03885_),
    .B1(_03801_),
    .B2(_03660_),
    .C(_05033_),
    .Y(_05034_));
 OA33x2_ASAP7_75t_R _11909_ (.A1(_03897_),
    .A2(_00322_),
    .A3(_03671_),
    .B1(_04344_),
    .B2(_03679_),
    .B3(_00321_),
    .Y(_05035_));
 AND4x1_ASAP7_75t_R _11910_ (.A(_03518_),
    .B(_03653_),
    .C(_05034_),
    .D(_05035_),
    .Y(_05036_));
 AND3x1_ASAP7_75t_R _11911_ (.A(_00318_),
    .B(_03813_),
    .C(_03775_),
    .Y(_05037_));
 AO21x1_ASAP7_75t_R _11912_ (.A1(_03701_),
    .A2(_05037_),
    .B(_03723_),
    .Y(_05038_));
 AOI211x1_ASAP7_75t_R _11913_ (.A1(_03701_),
    .A2(_05032_),
    .B(_05036_),
    .C(_05038_),
    .Y(_05039_));
 AND3x1_ASAP7_75t_R _11914_ (.A(_03663_),
    .B(_03853_),
    .C(_00308_),
    .Y(_05040_));
 AO21x1_ASAP7_75t_R _11915_ (.A1(_00307_),
    .A2(_03711_),
    .B(_05040_),
    .Y(_05041_));
 INVx1_ASAP7_75t_R _11916_ (.A(_00309_),
    .Y(_05042_));
 AND2x2_ASAP7_75t_R _11917_ (.A(_03609_),
    .B(_00314_),
    .Y(_05043_));
 AO21x1_ASAP7_75t_R _11918_ (.A1(_04457_),
    .A2(_00310_),
    .B(_05043_),
    .Y(_05044_));
 AOI22x1_ASAP7_75t_R _11919_ (.A1(_00313_),
    .A2(_04576_),
    .B1(_05044_),
    .B2(_03762_),
    .Y(_05045_));
 OA211x2_ASAP7_75t_R _11920_ (.A1(_04811_),
    .A2(_05045_),
    .B(_03607_),
    .C(_03646_),
    .Y(_05046_));
 OAI22x1_ASAP7_75t_R _11921_ (.A1(_05042_),
    .A2(_04575_),
    .B1(_05046_),
    .B2(_03785_),
    .Y(_05047_));
 OA22x2_ASAP7_75t_R _11922_ (.A1(_00311_),
    .A2(_03690_),
    .B1(_04945_),
    .B2(_00316_),
    .Y(_05048_));
 OA22x2_ASAP7_75t_R _11923_ (.A1(_00312_),
    .A2(_04949_),
    .B1(_05048_),
    .B2(_03607_),
    .Y(_05049_));
 OA211x2_ASAP7_75t_R _11924_ (.A1(_00315_),
    .A2(_04944_),
    .B(_05049_),
    .C(_03697_),
    .Y(_05050_));
 OR2x2_ASAP7_75t_R _11925_ (.A(_00302_),
    .B(_03620_),
    .Y(_05051_));
 AND3x1_ASAP7_75t_R _11926_ (.A(_03402_),
    .B(_03633_),
    .C(_00304_),
    .Y(_05052_));
 AO21x1_ASAP7_75t_R _11927_ (.A1(_00303_),
    .A2(_03709_),
    .B(_05052_),
    .Y(_05053_));
 OA211x2_ASAP7_75t_R _11928_ (.A1(_03801_),
    .A2(_05053_),
    .B(_04192_),
    .C(_04350_),
    .Y(_05054_));
 AND3x1_ASAP7_75t_R _11929_ (.A(_03549_),
    .B(_03624_),
    .C(_00306_),
    .Y(_05055_));
 AO21x1_ASAP7_75t_R _11930_ (.A1(_00305_),
    .A2(_03890_),
    .B(_05055_),
    .Y(_05056_));
 AO221x1_ASAP7_75t_R _11931_ (.A1(_05051_),
    .A2(_05054_),
    .B1(_05056_),
    .B2(_04727_),
    .C(_04194_),
    .Y(_05057_));
 AOI221x1_ASAP7_75t_R _11932_ (.A1(_04440_),
    .A2(_05041_),
    .B1(_05047_),
    .B2(_05050_),
    .C(_05057_),
    .Y(_05058_));
 AO21x2_ASAP7_75t_R _11933_ (.A1(_05029_),
    .A2(_05039_),
    .B(_05058_),
    .Y(_05059_));
 BUFx6f_ASAP7_75t_R _11934_ (.A(_05059_),
    .Y(_09992_));
 INVx4_ASAP7_75t_R _11935_ (.A(_09992_),
    .Y(_09994_));
 AO21x1_ASAP7_75t_R _11936_ (.A1(_04406_),
    .A2(_04849_),
    .B(_04251_),
    .Y(_05060_));
 AND2x2_ASAP7_75t_R _11937_ (.A(_04253_),
    .B(_05060_),
    .Y(_10152_));
 AND2x2_ASAP7_75t_R _11938_ (.A(_04034_),
    .B(_00350_),
    .Y(_05061_));
 AO21x1_ASAP7_75t_R _11939_ (.A1(_04265_),
    .A2(_00349_),
    .B(_05061_),
    .Y(_05062_));
 AND3x1_ASAP7_75t_R _11940_ (.A(_04127_),
    .B(_03380_),
    .C(_00348_),
    .Y(_05063_));
 AO21x1_ASAP7_75t_R _11941_ (.A1(_00347_),
    .A2(_04141_),
    .B(_05063_),
    .Y(_05064_));
 AO221x1_ASAP7_75t_R _11942_ (.A1(_04656_),
    .A2(_05062_),
    .B1(_05064_),
    .B2(_04145_),
    .C(_04008_),
    .Y(_05065_));
 AND2x2_ASAP7_75t_R _11943_ (.A(_04076_),
    .B(_00345_),
    .Y(_05066_));
 AO21x1_ASAP7_75t_R _11944_ (.A1(_04074_),
    .A2(_00343_),
    .B(_05066_),
    .Y(_05067_));
 AO21x1_ASAP7_75t_R _11945_ (.A1(_00344_),
    .A2(_04983_),
    .B(_04032_),
    .Y(_05068_));
 AO221x1_ASAP7_75t_R _11946_ (.A1(_00346_),
    .A2(_04091_),
    .B1(_05067_),
    .B2(_04080_),
    .C(_05068_),
    .Y(_05069_));
 AND2x2_ASAP7_75t_R _11947_ (.A(_04992_),
    .B(_00338_),
    .Y(_05070_));
 AO21x1_ASAP7_75t_R _11948_ (.A1(_04079_),
    .A2(_00337_),
    .B(_05070_),
    .Y(_05071_));
 AO21x1_ASAP7_75t_R _11949_ (.A1(_04988_),
    .A2(_05071_),
    .B(_04119_),
    .Y(_05072_));
 BUFx6f_ASAP7_75t_R _11950_ (.A(_03988_),
    .Y(_05073_));
 AO22x1_ASAP7_75t_R _11951_ (.A1(_04671_),
    .A2(_00335_),
    .B1(_00336_),
    .B2(_05073_),
    .Y(_05074_));
 AO22x1_ASAP7_75t_R _11952_ (.A1(_04504_),
    .A2(_00335_),
    .B1(_05074_),
    .B2(_04074_),
    .Y(_05075_));
 AO21x1_ASAP7_75t_R _11953_ (.A1(_04060_),
    .A2(_05072_),
    .B(_05075_),
    .Y(_05076_));
 AND2x2_ASAP7_75t_R _11954_ (.A(_04034_),
    .B(_00342_),
    .Y(_05077_));
 AO21x1_ASAP7_75t_R _11955_ (.A1(_04265_),
    .A2(_00341_),
    .B(_05077_),
    .Y(_05078_));
 AND3x1_ASAP7_75t_R _11956_ (.A(_04034_),
    .B(_03380_),
    .C(_00340_),
    .Y(_05079_));
 AO21x1_ASAP7_75t_R _11957_ (.A1(_00339_),
    .A2(_04141_),
    .B(_05079_),
    .Y(_05080_));
 AOI221x1_ASAP7_75t_R _11958_ (.A1(_04656_),
    .A2(_05078_),
    .B1(_05080_),
    .B2(_04145_),
    .C(_04008_),
    .Y(_05081_));
 NOR2x1_ASAP7_75t_R _11959_ (.A(_04157_),
    .B(_05081_),
    .Y(_05082_));
 AO32x1_ASAP7_75t_R _11960_ (.A1(_04157_),
    .A2(_05065_),
    .A3(_05069_),
    .B1(_05076_),
    .B2(_05082_),
    .Y(_05083_));
 AND2x2_ASAP7_75t_R _11961_ (.A(_04127_),
    .B(_00358_),
    .Y(_05084_));
 AO21x1_ASAP7_75t_R _11962_ (.A1(_04126_),
    .A2(_00357_),
    .B(_05084_),
    .Y(_05085_));
 AND3x1_ASAP7_75t_R _11963_ (.A(_04138_),
    .B(_03380_),
    .C(_00356_),
    .Y(_05086_));
 AO21x1_ASAP7_75t_R _11964_ (.A1(_00355_),
    .A2(_04141_),
    .B(_05086_),
    .Y(_05087_));
 AO221x1_ASAP7_75t_R _11965_ (.A1(_04067_),
    .A2(_05085_),
    .B1(_05087_),
    .B2(_04145_),
    .C(_04298_),
    .Y(_05088_));
 AND2x2_ASAP7_75t_R _11966_ (.A(_04127_),
    .B(_00366_),
    .Y(_05089_));
 AO21x1_ASAP7_75t_R _11967_ (.A1(_04126_),
    .A2(_00365_),
    .B(_05089_),
    .Y(_05090_));
 AND3x1_ASAP7_75t_R _11968_ (.A(_04138_),
    .B(_03380_),
    .C(_00364_),
    .Y(_05091_));
 AO21x1_ASAP7_75t_R _11969_ (.A1(_00363_),
    .A2(_04141_),
    .B(_05091_),
    .Y(_05092_));
 AO221x1_ASAP7_75t_R _11970_ (.A1(_04067_),
    .A2(_05090_),
    .B1(_05092_),
    .B2(_04145_),
    .C(_04304_),
    .Y(_05093_));
 AND3x1_ASAP7_75t_R _11971_ (.A(_04124_),
    .B(_05088_),
    .C(_05093_),
    .Y(_05094_));
 AO221x1_ASAP7_75t_R _11972_ (.A1(_04289_),
    .A2(_00362_),
    .B1(_04069_),
    .B2(_00360_),
    .C(_03997_),
    .Y(_05095_));
 AO221x1_ASAP7_75t_R _11973_ (.A1(_03927_),
    .A2(_00354_),
    .B1(_04069_),
    .B2(_00352_),
    .C(_04156_),
    .Y(_05096_));
 AND3x1_ASAP7_75t_R _11974_ (.A(_04066_),
    .B(_05095_),
    .C(_05096_),
    .Y(_05097_));
 AND2x2_ASAP7_75t_R _11975_ (.A(_04987_),
    .B(_00361_),
    .Y(_05098_));
 AO21x1_ASAP7_75t_R _11976_ (.A1(_04074_),
    .A2(_00359_),
    .B(_05098_),
    .Y(_05099_));
 AND2x2_ASAP7_75t_R _11977_ (.A(_03926_),
    .B(_00353_),
    .Y(_05100_));
 AO221x1_ASAP7_75t_R _11978_ (.A1(_04112_),
    .A2(_03972_),
    .B1(_00351_),
    .B2(_04114_),
    .C(_05100_),
    .Y(_05101_));
 OA211x2_ASAP7_75t_R _11979_ (.A1(_04514_),
    .A2(_05099_),
    .B(_05101_),
    .C(_04089_),
    .Y(_05102_));
 OR3x1_ASAP7_75t_R _11980_ (.A(_04120_),
    .B(_05097_),
    .C(_05102_),
    .Y(_05103_));
 AO221x2_ASAP7_75t_R _11981_ (.A1(_04122_),
    .A2(_05083_),
    .B1(_05094_),
    .B2(_05103_),
    .C(_04565_),
    .Y(_05104_));
 NOR2x1_ASAP7_75t_R _11982_ (.A(_04254_),
    .B(_05104_),
    .Y(_05105_));
 AOI21x1_ASAP7_75t_R _11983_ (.A1(_04250_),
    .A2(_10152_),
    .B(_05105_),
    .Y(_05106_));
 XNOR2x1_ASAP7_75t_R _11984_ (.B(_05106_),
    .Y(_10000_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _11985_ (.A(_10000_),
    .Y(_09998_));
 INVx2_ASAP7_75t_R _11986_ (.A(_00359_),
    .Y(_05107_));
 AND2x2_ASAP7_75t_R _11987_ (.A(_03685_),
    .B(_00364_),
    .Y(_05108_));
 AO21x1_ASAP7_75t_R _11988_ (.A1(_03744_),
    .A2(_00360_),
    .B(_05108_),
    .Y(_05109_));
 AOI22x1_ASAP7_75t_R _11989_ (.A1(_00363_),
    .A2(_04456_),
    .B1(_05109_),
    .B2(_04435_),
    .Y(_05110_));
 OA211x2_ASAP7_75t_R _11990_ (.A1(_03480_),
    .A2(_05110_),
    .B(_03607_),
    .C(_03860_),
    .Y(_05111_));
 OAI22x1_ASAP7_75t_R _11991_ (.A1(_05107_),
    .A2(_04218_),
    .B1(_05111_),
    .B2(_04163_),
    .Y(_05112_));
 AND3x1_ASAP7_75t_R _11992_ (.A(_03402_),
    .B(_03633_),
    .C(_00362_),
    .Y(_05113_));
 AO21x1_ASAP7_75t_R _11993_ (.A1(_00361_),
    .A2(_03612_),
    .B(_05113_),
    .Y(_05114_));
 OR3x1_ASAP7_75t_R _11994_ (.A(_03679_),
    .B(_03669_),
    .C(_05114_),
    .Y(_05115_));
 AND2x2_ASAP7_75t_R _11995_ (.A(_00365_),
    .B(_03709_),
    .Y(_05116_));
 AO221x1_ASAP7_75t_R _11996_ (.A1(_00366_),
    .A2(_03885_),
    .B1(_03661_),
    .B2(_04350_),
    .C(_05116_),
    .Y(_05117_));
 AO21x1_ASAP7_75t_R _11997_ (.A1(_05115_),
    .A2(_05117_),
    .B(_04229_),
    .Y(_05118_));
 OA211x2_ASAP7_75t_R _11998_ (.A1(_03723_),
    .A2(_05112_),
    .B(_05118_),
    .C(_04231_),
    .Y(_05119_));
 OR3x1_ASAP7_75t_R _11999_ (.A(_00352_),
    .B(_03679_),
    .C(_03681_),
    .Y(_05120_));
 AO21x1_ASAP7_75t_R _12000_ (.A1(_03646_),
    .A2(_03607_),
    .B(_00354_),
    .Y(_05121_));
 AO21x1_ASAP7_75t_R _12001_ (.A1(_05120_),
    .A2(_05121_),
    .B(_03714_),
    .Y(_05122_));
 OR2x2_ASAP7_75t_R _12002_ (.A(_00353_),
    .B(_03865_),
    .Y(_05123_));
 OA21x2_ASAP7_75t_R _12003_ (.A1(_00351_),
    .A2(_03759_),
    .B(_03701_),
    .Y(_05124_));
 OR3x1_ASAP7_75t_R _12004_ (.A(_00356_),
    .B(_03679_),
    .C(_03681_),
    .Y(_05125_));
 AO21x1_ASAP7_75t_R _12005_ (.A1(_03646_),
    .A2(_03607_),
    .B(_00358_),
    .Y(_05126_));
 AO21x1_ASAP7_75t_R _12006_ (.A1(_05125_),
    .A2(_05126_),
    .B(_03714_),
    .Y(_05127_));
 OR3x1_ASAP7_75t_R _12007_ (.A(_00355_),
    .B(_04233_),
    .C(_04344_),
    .Y(_05128_));
 AO221x1_ASAP7_75t_R _12008_ (.A1(_03549_),
    .A2(_03624_),
    .B1(_03827_),
    .B2(_03593_),
    .C(_00357_),
    .Y(_05129_));
 AND4x1_ASAP7_75t_R _12009_ (.A(_04244_),
    .B(_03653_),
    .C(_05128_),
    .D(_05129_),
    .Y(_05130_));
 AO32x2_ASAP7_75t_R _12010_ (.A1(_05122_),
    .A2(_05123_),
    .A3(_05124_),
    .B1(_05127_),
    .B2(_05130_),
    .Y(_05131_));
 INVx1_ASAP7_75t_R _12011_ (.A(_00343_),
    .Y(_05132_));
 AND2x2_ASAP7_75t_R _12012_ (.A(_03609_),
    .B(_00348_),
    .Y(_05133_));
 AO21x1_ASAP7_75t_R _12013_ (.A1(_04457_),
    .A2(_00344_),
    .B(_05133_),
    .Y(_05134_));
 AOI22x1_ASAP7_75t_R _12014_ (.A1(_00347_),
    .A2(_04456_),
    .B1(_05134_),
    .B2(_04460_),
    .Y(_05135_));
 OA211x2_ASAP7_75t_R _12015_ (.A1(_04811_),
    .A2(_05135_),
    .B(_03607_),
    .C(_03860_),
    .Y(_05136_));
 OAI22x1_ASAP7_75t_R _12016_ (.A1(_05132_),
    .A2(_04218_),
    .B1(_05136_),
    .B2(_03785_),
    .Y(_05137_));
 AND3x1_ASAP7_75t_R _12017_ (.A(_00346_),
    .B(_04350_),
    .C(_03661_),
    .Y(_05138_));
 OA21x2_ASAP7_75t_R _12018_ (.A1(_03679_),
    .A2(_03669_),
    .B(_00350_),
    .Y(_05139_));
 AND3x1_ASAP7_75t_R _12019_ (.A(_00345_),
    .B(_03660_),
    .C(_03661_),
    .Y(_05140_));
 OA21x2_ASAP7_75t_R _12020_ (.A1(_03679_),
    .A2(_03669_),
    .B(_00349_),
    .Y(_05141_));
 OA33x2_ASAP7_75t_R _12021_ (.A1(_03869_),
    .A2(_05138_),
    .A3(_05139_),
    .B1(_05140_),
    .B2(_05141_),
    .B3(_03865_),
    .Y(_05142_));
 AND3x1_ASAP7_75t_R _12022_ (.A(_03698_),
    .B(_05137_),
    .C(_05142_),
    .Y(_05143_));
 OA211x2_ASAP7_75t_R _12023_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03727_),
    .C(_00340_),
    .Y(_05144_));
 AO21x1_ASAP7_75t_R _12024_ (.A1(_00339_),
    .A2(_03585_),
    .B(_05144_),
    .Y(_05145_));
 OA222x2_ASAP7_75t_R _12025_ (.A1(_00341_),
    .A2(_03885_),
    .B1(_03584_),
    .B2(_00342_),
    .C1(_03681_),
    .C2(_03679_),
    .Y(_05146_));
 AO21x1_ASAP7_75t_R _12026_ (.A1(_04454_),
    .A2(_05145_),
    .B(_05146_),
    .Y(_05147_));
 INVx1_ASAP7_75t_R _12027_ (.A(_00337_),
    .Y(_05148_));
 INVx2_ASAP7_75t_R _12028_ (.A(_00336_),
    .Y(_05149_));
 NAND2x1_ASAP7_75t_R _12029_ (.A(_03619_),
    .B(_00338_),
    .Y(_05150_));
 OA211x2_ASAP7_75t_R _12030_ (.A1(_03636_),
    .A2(_05149_),
    .B(_05150_),
    .C(_03633_),
    .Y(_05151_));
 AOI21x1_ASAP7_75t_R _12031_ (.A1(_05148_),
    .A2(_04185_),
    .B(_05151_),
    .Y(_05152_));
 OA211x2_ASAP7_75t_R _12032_ (.A1(_03480_),
    .A2(_05152_),
    .B(_03771_),
    .C(_04350_),
    .Y(_05153_));
 OA22x2_ASAP7_75t_R _12033_ (.A1(_00335_),
    .A2(_03759_),
    .B1(_05153_),
    .B2(_04163_),
    .Y(_05154_));
 AO211x2_ASAP7_75t_R _12034_ (.A1(_03791_),
    .A2(_05147_),
    .B(_05154_),
    .C(_04195_),
    .Y(_05155_));
 OA22x2_ASAP7_75t_R _12035_ (.A1(_05119_),
    .A2(_05131_),
    .B1(_05143_),
    .B2(_05155_),
    .Y(_05156_));
 BUFx3_ASAP7_75t_R _12036_ (.A(_05156_),
    .Y(_09997_));
 INVx6_ASAP7_75t_R _12037_ (.A(_09997_),
    .Y(_09999_));
 AO21x1_ASAP7_75t_R _12038_ (.A1(_04849_),
    .A2(_04412_),
    .B(_04251_),
    .Y(_05157_));
 AND2x2_ASAP7_75t_R _12039_ (.A(_04253_),
    .B(_05157_),
    .Y(_10150_));
 AO221x1_ASAP7_75t_R _12040_ (.A1(_04643_),
    .A2(_00391_),
    .B1(_04069_),
    .B2(_00389_),
    .C(_04265_),
    .Y(_05158_));
 AND2x2_ASAP7_75t_R _12041_ (.A(_04529_),
    .B(_00390_),
    .Y(_05159_));
 AO211x2_ASAP7_75t_R _12042_ (.A1(_04074_),
    .A2(_00388_),
    .B(_05159_),
    .C(_04308_),
    .Y(_05160_));
 AO221x1_ASAP7_75t_R _12043_ (.A1(_04072_),
    .A2(_00388_),
    .B1(_05158_),
    .B2(_05160_),
    .C(_03921_),
    .Y(_05161_));
 AND2x2_ASAP7_75t_R _12044_ (.A(_04270_),
    .B(_00398_),
    .Y(_05162_));
 AO21x1_ASAP7_75t_R _12045_ (.A1(_04074_),
    .A2(_00396_),
    .B(_05162_),
    .Y(_05163_));
 AO21x1_ASAP7_75t_R _12046_ (.A1(_00399_),
    .A2(_03962_),
    .B(_04009_),
    .Y(_05164_));
 AO221x1_ASAP7_75t_R _12047_ (.A1(_00397_),
    .A2(_04083_),
    .B1(_05163_),
    .B2(_04089_),
    .C(_05164_),
    .Y(_05165_));
 AOI21x1_ASAP7_75t_R _12048_ (.A1(_05161_),
    .A2(_05165_),
    .B(_04095_),
    .Y(_05166_));
 INVx1_ASAP7_75t_R _12049_ (.A(_00392_),
    .Y(_05167_));
 NAND2x1_ASAP7_75t_R _12050_ (.A(_04076_),
    .B(_00394_),
    .Y(_05168_));
 OA211x2_ASAP7_75t_R _12051_ (.A1(_04643_),
    .A2(_05167_),
    .B(_05168_),
    .C(_04079_),
    .Y(_05169_));
 INVx1_ASAP7_75t_R _12052_ (.A(_00395_),
    .Y(_05170_));
 OA21x2_ASAP7_75t_R _12053_ (.A1(_04104_),
    .A2(_05170_),
    .B(_04016_),
    .Y(_05171_));
 INVx1_ASAP7_75t_R _12054_ (.A(_00393_),
    .Y(_05172_));
 OR4x1_ASAP7_75t_R _12055_ (.A(_04531_),
    .B(_04270_),
    .C(_03984_),
    .D(_05172_),
    .Y(_05173_));
 OA211x2_ASAP7_75t_R _12056_ (.A1(_05169_),
    .A2(_05171_),
    .B(_03921_),
    .C(_05173_),
    .Y(_05174_));
 INVx1_ASAP7_75t_R _12057_ (.A(_00384_),
    .Y(_05175_));
 NAND2x1_ASAP7_75t_R _12058_ (.A(_04076_),
    .B(_00386_),
    .Y(_05176_));
 OA211x2_ASAP7_75t_R _12059_ (.A1(_04643_),
    .A2(_05175_),
    .B(_05176_),
    .C(_04647_),
    .Y(_05177_));
 INVx1_ASAP7_75t_R _12060_ (.A(_00387_),
    .Y(_05178_));
 OA21x2_ASAP7_75t_R _12061_ (.A1(_04104_),
    .A2(_05178_),
    .B(_04016_),
    .Y(_05179_));
 INVx1_ASAP7_75t_R _12062_ (.A(_00385_),
    .Y(_05180_));
 OR4x1_ASAP7_75t_R _12063_ (.A(_04556_),
    .B(_04270_),
    .C(_03984_),
    .D(_05180_),
    .Y(_05181_));
 OA211x2_ASAP7_75t_R _12064_ (.A1(_05177_),
    .A2(_05179_),
    .B(_04098_),
    .C(_05181_),
    .Y(_05182_));
 OA21x2_ASAP7_75t_R _12065_ (.A1(_05174_),
    .A2(_05182_),
    .B(_04296_),
    .Y(_05183_));
 OAI21x1_ASAP7_75t_R _12066_ (.A1(_05166_),
    .A2(_05183_),
    .B(_04124_),
    .Y(_05184_));
 AND2x2_ASAP7_75t_R _12067_ (.A(_04034_),
    .B(_00383_),
    .Y(_05185_));
 AO21x1_ASAP7_75t_R _12068_ (.A1(_04126_),
    .A2(_00382_),
    .B(_05185_),
    .Y(_05186_));
 AND3x1_ASAP7_75t_R _12069_ (.A(_04127_),
    .B(_03380_),
    .C(_00381_),
    .Y(_05187_));
 AO21x1_ASAP7_75t_R _12070_ (.A1(_00380_),
    .A2(_04141_),
    .B(_05187_),
    .Y(_05188_));
 AO221x1_ASAP7_75t_R _12071_ (.A1(_04656_),
    .A2(_05186_),
    .B1(_05188_),
    .B2(_04145_),
    .C(_04008_),
    .Y(_05189_));
 AND2x2_ASAP7_75t_R _12072_ (.A(_04544_),
    .B(_00378_),
    .Y(_05190_));
 AO21x1_ASAP7_75t_R _12073_ (.A1(_04084_),
    .A2(_00376_),
    .B(_05190_),
    .Y(_05191_));
 AO22x1_ASAP7_75t_R _12074_ (.A1(_00379_),
    .A2(_03962_),
    .B1(_05191_),
    .B2(_04126_),
    .Y(_05192_));
 AO21x1_ASAP7_75t_R _12075_ (.A1(_00377_),
    .A2(_04083_),
    .B(_04119_),
    .Y(_05193_));
 OA21x2_ASAP7_75t_R _12076_ (.A1(_05192_),
    .A2(_05193_),
    .B(_04157_),
    .Y(_05194_));
 AO22x1_ASAP7_75t_R _12077_ (.A1(_04265_),
    .A2(_00368_),
    .B1(_00369_),
    .B2(_04102_),
    .Y(_05195_));
 AND2x2_ASAP7_75t_R _12078_ (.A(_04015_),
    .B(_00371_),
    .Y(_05196_));
 AO21x1_ASAP7_75t_R _12079_ (.A1(_04556_),
    .A2(_00370_),
    .B(_05196_),
    .Y(_05197_));
 AO21x1_ASAP7_75t_R _12080_ (.A1(_04530_),
    .A2(_05197_),
    .B(_04032_),
    .Y(_05198_));
 AND2x2_ASAP7_75t_R _12081_ (.A(_04504_),
    .B(_00368_),
    .Y(_05199_));
 AO221x1_ASAP7_75t_R _12082_ (.A1(_04085_),
    .A2(_05195_),
    .B1(_05198_),
    .B2(_04060_),
    .C(_05199_),
    .Y(_05200_));
 AND2x2_ASAP7_75t_R _12083_ (.A(_04307_),
    .B(_00375_),
    .Y(_05201_));
 AO21x1_ASAP7_75t_R _12084_ (.A1(_04088_),
    .A2(_00374_),
    .B(_05201_),
    .Y(_05202_));
 AO21x1_ASAP7_75t_R _12085_ (.A1(_04656_),
    .A2(_05202_),
    .B(_04542_),
    .Y(_05203_));
 AND3x1_ASAP7_75t_R _12086_ (.A(_04138_),
    .B(_04142_),
    .C(_00373_),
    .Y(_05204_));
 OA21x2_ASAP7_75t_R _12087_ (.A1(_04531_),
    .A2(_04071_),
    .B(_00372_),
    .Y(_05205_));
 OA21x2_ASAP7_75t_R _12088_ (.A1(_05204_),
    .A2(_05205_),
    .B(_04996_),
    .Y(_05206_));
 OA21x2_ASAP7_75t_R _12089_ (.A1(_05203_),
    .A2(_05206_),
    .B(_04514_),
    .Y(_05207_));
 AO221x1_ASAP7_75t_R _12090_ (.A1(_05189_),
    .A2(_05194_),
    .B1(_05200_),
    .B2(_05207_),
    .C(_04124_),
    .Y(_05208_));
 AOI21x1_ASAP7_75t_R _12091_ (.A1(_05184_),
    .A2(_05208_),
    .B(_04565_),
    .Y(_05209_));
 AND2x2_ASAP7_75t_R _12092_ (.A(_04059_),
    .B(_05209_),
    .Y(_05210_));
 AO21x1_ASAP7_75t_R _12093_ (.A1(_04250_),
    .A2(_10150_),
    .B(_05210_),
    .Y(_05211_));
 XNOR2x1_ASAP7_75t_R _12094_ (.B(_05211_),
    .Y(_10005_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _12095_ (.A(_10005_),
    .Y(_10003_));
 AND3x1_ASAP7_75t_R _12096_ (.A(_04596_),
    .B(_04436_),
    .C(_00387_),
    .Y(_05212_));
 AO21x1_ASAP7_75t_R _12097_ (.A1(_00386_),
    .A2(_04595_),
    .B(_05212_),
    .Y(_05213_));
 AO222x2_ASAP7_75t_R _12098_ (.A1(_00384_),
    .A2(_03703_),
    .B1(_04628_),
    .B2(_00385_),
    .C1(_05213_),
    .C2(_03733_),
    .Y(_05214_));
 BUFx12_ASAP7_75t_R _12099_ (.A(_04460_),
    .Y(_05215_));
 AND3x1_ASAP7_75t_R _12100_ (.A(_03376_),
    .B(_05215_),
    .C(_00391_),
    .Y(_05216_));
 AO21x1_ASAP7_75t_R _12101_ (.A1(_00390_),
    .A2(_04434_),
    .B(_05216_),
    .Y(_05217_));
 BUFx10_ASAP7_75t_R _12102_ (.A(_03825_),
    .Y(_05218_));
 OA222x2_ASAP7_75t_R _12103_ (.A1(_00389_),
    .A2(_04952_),
    .B1(_05217_),
    .B2(_05218_),
    .C1(_04492_),
    .C2(_00388_),
    .Y(_05219_));
 AOI221x1_ASAP7_75t_R _12104_ (.A1(_04915_),
    .A2(_05214_),
    .B1(_05219_),
    .B2(_03792_),
    .C(_03809_),
    .Y(_05220_));
 BUFx12f_ASAP7_75t_R _12105_ (.A(_04576_),
    .Y(_05221_));
 AND2x2_ASAP7_75t_R _12106_ (.A(_04938_),
    .B(_00397_),
    .Y(_05222_));
 AO21x1_ASAP7_75t_R _12107_ (.A1(_04937_),
    .A2(_00393_),
    .B(_05222_),
    .Y(_05223_));
 BUFx12_ASAP7_75t_R _12108_ (.A(_04460_),
    .Y(_05224_));
 AO22x1_ASAP7_75t_R _12109_ (.A1(_00396_),
    .A2(_05221_),
    .B1(_05223_),
    .B2(_05224_),
    .Y(_05225_));
 NAND2x1_ASAP7_75t_R _12110_ (.A(_03377_),
    .B(_05225_),
    .Y(_05226_));
 BUFx16f_ASAP7_75t_R _12111_ (.A(_03785_),
    .Y(_05227_));
 AO21x1_ASAP7_75t_R _12112_ (.A1(_05218_),
    .A2(_05226_),
    .B(_05227_),
    .Y(_05228_));
 NAND2x1_ASAP7_75t_R _12113_ (.A(_00392_),
    .B(_03811_),
    .Y(_05229_));
 BUFx10_ASAP7_75t_R _12114_ (.A(_04198_),
    .Y(_05230_));
 AND3x1_ASAP7_75t_R _12115_ (.A(_00394_),
    .B(_03804_),
    .C(_03831_),
    .Y(_05231_));
 AOI221x1_ASAP7_75t_R _12116_ (.A1(_00399_),
    .A2(_05230_),
    .B1(_04476_),
    .B2(_00398_),
    .C(_05231_),
    .Y(_05232_));
 BUFx10_ASAP7_75t_R _12117_ (.A(_03834_),
    .Y(_05233_));
 AOI21x1_ASAP7_75t_R _12118_ (.A1(_00395_),
    .A2(_05233_),
    .B(_04792_),
    .Y(_05234_));
 BUFx6f_ASAP7_75t_R _12119_ (.A(_04468_),
    .Y(_05235_));
 AO221x2_ASAP7_75t_R _12120_ (.A1(_05228_),
    .A2(_05229_),
    .B1(_05232_),
    .B2(_05234_),
    .C(_05235_),
    .Y(_05236_));
 AND3x1_ASAP7_75t_R _12121_ (.A(_00379_),
    .B(_03777_),
    .C(_03838_),
    .Y(_05237_));
 AOI211x1_ASAP7_75t_R _12122_ (.A1(_00383_),
    .A2(_03872_),
    .B(_03869_),
    .C(_05237_),
    .Y(_05238_));
 INVx1_ASAP7_75t_R _12123_ (.A(_00376_),
    .Y(_05239_));
 AND2x2_ASAP7_75t_R _12124_ (.A(_03610_),
    .B(_00381_),
    .Y(_05240_));
 AO21x1_ASAP7_75t_R _12125_ (.A1(_04609_),
    .A2(_00377_),
    .B(_05240_),
    .Y(_05241_));
 AOI22x1_ASAP7_75t_R _12126_ (.A1(_00380_),
    .A2(_04800_),
    .B1(_05241_),
    .B2(_04584_),
    .Y(_05242_));
 OA211x2_ASAP7_75t_R _12127_ (.A1(_03481_),
    .A2(_05242_),
    .B(_04804_),
    .C(_04478_),
    .Y(_05243_));
 OA22x2_ASAP7_75t_R _12128_ (.A1(_05239_),
    .A2(_04575_),
    .B1(_05243_),
    .B2(_04164_),
    .Y(_05244_));
 AND3x1_ASAP7_75t_R _12129_ (.A(_00378_),
    .B(_03777_),
    .C(_03874_),
    .Y(_05245_));
 AOI211x1_ASAP7_75t_R _12130_ (.A1(_00382_),
    .A2(_03872_),
    .B(_03866_),
    .C(_05245_),
    .Y(_05246_));
 OR4x2_ASAP7_75t_R _12131_ (.A(_04468_),
    .B(_05238_),
    .C(_05244_),
    .D(_05246_),
    .Y(_05247_));
 AND3x1_ASAP7_75t_R _12132_ (.A(_04053_),
    .B(_04624_),
    .C(_00375_),
    .Y(_05248_));
 AO21x1_ASAP7_75t_R _12133_ (.A1(_00374_),
    .A2(_04623_),
    .B(_05248_),
    .Y(_05249_));
 AND2x2_ASAP7_75t_R _12134_ (.A(_00370_),
    .B(_04242_),
    .Y(_05250_));
 AO221x1_ASAP7_75t_R _12135_ (.A1(_00371_),
    .A2(_03882_),
    .B1(_04592_),
    .B2(_03829_),
    .C(_05250_),
    .Y(_05251_));
 OA211x2_ASAP7_75t_R _12136_ (.A1(_00369_),
    .A2(_04952_),
    .B(_04627_),
    .C(_05251_),
    .Y(_05252_));
 AND3x1_ASAP7_75t_R _12137_ (.A(_03797_),
    .B(_03798_),
    .C(_00373_),
    .Y(_05253_));
 AO21x1_ASAP7_75t_R _12138_ (.A1(_00372_),
    .A2(_04929_),
    .B(_05253_),
    .Y(_05254_));
 AO21x1_ASAP7_75t_R _12139_ (.A1(_04727_),
    .A2(_05254_),
    .B(_04959_),
    .Y(_05255_));
 AOI211x1_ASAP7_75t_R _12140_ (.A1(_04440_),
    .A2(_05249_),
    .B(_05252_),
    .C(_05255_),
    .Y(_05256_));
 AOI22x1_ASAP7_75t_R _12141_ (.A1(_05220_),
    .A2(_05236_),
    .B1(_05247_),
    .B2(_05256_),
    .Y(_10002_));
 INVx4_ASAP7_75t_R _12142_ (.A(_10002_),
    .Y(_10004_));
 AND2x2_ASAP7_75t_R _12143_ (.A(_04138_),
    .B(_00424_),
    .Y(_05257_));
 AO21x1_ASAP7_75t_R _12144_ (.A1(_04126_),
    .A2(_00423_),
    .B(_05257_),
    .Y(_05258_));
 AO21x1_ASAP7_75t_R _12145_ (.A1(_04067_),
    .A2(_05258_),
    .B(_04298_),
    .Y(_05259_));
 AND3x1_ASAP7_75t_R _12146_ (.A(_04127_),
    .B(_03380_),
    .C(_00422_),
    .Y(_05260_));
 AO21x1_ASAP7_75t_R _12147_ (.A1(_00421_),
    .A2(_04141_),
    .B(_05260_),
    .Y(_05261_));
 AND2x2_ASAP7_75t_R _12148_ (.A(_04145_),
    .B(_05261_),
    .Y(_05262_));
 AND2x2_ASAP7_75t_R _12149_ (.A(_04307_),
    .B(_00432_),
    .Y(_05263_));
 AO21x1_ASAP7_75t_R _12150_ (.A1(_04088_),
    .A2(_00431_),
    .B(_05263_),
    .Y(_05264_));
 AND3x1_ASAP7_75t_R _12151_ (.A(_04307_),
    .B(_04315_),
    .C(_00430_),
    .Y(_05265_));
 AO21x1_ASAP7_75t_R _12152_ (.A1(_00429_),
    .A2(_04991_),
    .B(_05265_),
    .Y(_05266_));
 AO221x1_ASAP7_75t_R _12153_ (.A1(_04988_),
    .A2(_05264_),
    .B1(_05266_),
    .B2(_04996_),
    .C(_04304_),
    .Y(_05267_));
 OA211x2_ASAP7_75t_R _12154_ (.A1(_05259_),
    .A2(_05262_),
    .B(_05267_),
    .C(_04763_),
    .Y(_05268_));
 AO221x1_ASAP7_75t_R _12155_ (.A1(_03975_),
    .A2(_00428_),
    .B1(_04632_),
    .B2(_00426_),
    .C(_04414_),
    .Y(_05269_));
 AO221x1_ASAP7_75t_R _12156_ (.A1(_03975_),
    .A2(_00420_),
    .B1(_04632_),
    .B2(_00418_),
    .C(_03920_),
    .Y(_05270_));
 AND3x1_ASAP7_75t_R _12157_ (.A(_04066_),
    .B(_05269_),
    .C(_05270_),
    .Y(_05271_));
 AND2x2_ASAP7_75t_R _12158_ (.A(_04106_),
    .B(_00427_),
    .Y(_05272_));
 AO21x1_ASAP7_75t_R _12159_ (.A1(_04104_),
    .A2(_00425_),
    .B(_05272_),
    .Y(_05273_));
 AND2x2_ASAP7_75t_R _12160_ (.A(_04544_),
    .B(_00419_),
    .Y(_05274_));
 AO221x1_ASAP7_75t_R _12161_ (.A1(_04111_),
    .A2(_04142_),
    .B1(_00417_),
    .B2(_04084_),
    .C(_05274_),
    .Y(_05275_));
 OA211x2_ASAP7_75t_R _12162_ (.A1(_04098_),
    .A2(_05273_),
    .B(_05275_),
    .C(_04080_),
    .Y(_05276_));
 OR3x1_ASAP7_75t_R _12163_ (.A(_04120_),
    .B(_05271_),
    .C(_05276_),
    .Y(_05277_));
 AND2x2_ASAP7_75t_R _12164_ (.A(_03974_),
    .B(_00411_),
    .Y(_05278_));
 AO21x1_ASAP7_75t_R _12165_ (.A1(_03992_),
    .A2(_00409_),
    .B(_05278_),
    .Y(_05279_));
 AO221x1_ASAP7_75t_R _12166_ (.A1(_04106_),
    .A2(_00412_),
    .B1(_04068_),
    .B2(_00410_),
    .C(_03930_),
    .Y(_05280_));
 OA21x2_ASAP7_75t_R _12167_ (.A1(_04308_),
    .A2(_05279_),
    .B(_05280_),
    .Y(_05281_));
 AND2x2_ASAP7_75t_R _12168_ (.A(_04033_),
    .B(_00416_),
    .Y(_05282_));
 AO21x1_ASAP7_75t_R _12169_ (.A1(_04281_),
    .A2(_00415_),
    .B(_05282_),
    .Y(_05283_));
 AND3x1_ASAP7_75t_R _12170_ (.A(_04256_),
    .B(_03379_),
    .C(_00414_),
    .Y(_05284_));
 AO21x1_ASAP7_75t_R _12171_ (.A1(_00413_),
    .A2(_03939_),
    .B(_05284_),
    .Y(_05285_));
 AO221x1_ASAP7_75t_R _12172_ (.A1(_04643_),
    .A2(_05283_),
    .B1(_05285_),
    .B2(_04995_),
    .C(_03947_),
    .Y(_05286_));
 OA211x2_ASAP7_75t_R _12173_ (.A1(_04131_),
    .A2(_05281_),
    .B(_05286_),
    .C(_03921_),
    .Y(_05287_));
 AND2x2_ASAP7_75t_R _12174_ (.A(_04137_),
    .B(_00408_),
    .Y(_05288_));
 AO21x1_ASAP7_75t_R _12175_ (.A1(_03930_),
    .A2(_00407_),
    .B(_05288_),
    .Y(_05289_));
 AND3x1_ASAP7_75t_R _12176_ (.A(_03942_),
    .B(_03943_),
    .C(_00406_),
    .Y(_05290_));
 AO21x1_ASAP7_75t_R _12177_ (.A1(_00405_),
    .A2(_04292_),
    .B(_05290_),
    .Y(_05291_));
 AO221x1_ASAP7_75t_R _12178_ (.A1(_04289_),
    .A2(_05289_),
    .B1(_05291_),
    .B2(_04295_),
    .C(_04094_),
    .Y(_05292_));
 AO22x1_ASAP7_75t_R _12179_ (.A1(_04556_),
    .A2(_00401_),
    .B1(_00402_),
    .B2(_04522_),
    .Y(_05293_));
 AND2x2_ASAP7_75t_R _12180_ (.A(_04536_),
    .B(_00404_),
    .Y(_05294_));
 AO21x1_ASAP7_75t_R _12181_ (.A1(_04028_),
    .A2(_00403_),
    .B(_05294_),
    .Y(_05295_));
 AO221x1_ASAP7_75t_R _12182_ (.A1(_03984_),
    .A2(_00401_),
    .B1(_04412_),
    .B2(_05295_),
    .C(_04406_),
    .Y(_05296_));
 AO21x1_ASAP7_75t_R _12183_ (.A1(_04074_),
    .A2(_05293_),
    .B(_05296_),
    .Y(_05297_));
 AND3x1_ASAP7_75t_R _12184_ (.A(_04514_),
    .B(_05292_),
    .C(_05297_),
    .Y(_05298_));
 OA21x2_ASAP7_75t_R _12185_ (.A1(_05287_),
    .A2(_05298_),
    .B(_03917_),
    .Y(_05299_));
 AOI211x1_ASAP7_75t_R _12186_ (.A1(_05268_),
    .A2(_05277_),
    .B(_05299_),
    .C(_04565_),
    .Y(_05300_));
 AO21x1_ASAP7_75t_R _12187_ (.A1(_04849_),
    .A2(_04102_),
    .B(_04251_),
    .Y(_05301_));
 AND3x1_ASAP7_75t_R _12188_ (.A(_04162_),
    .B(_04253_),
    .C(_05301_),
    .Y(_05302_));
 AOI21x1_ASAP7_75t_R _12189_ (.A1(_04065_),
    .A2(_05300_),
    .B(_05302_),
    .Y(_05303_));
 XNOR2x1_ASAP7_75t_R _12190_ (.B(_05303_),
    .Y(_10008_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _12191_ (.A(_10008_),
    .Y(_10010_));
 OA211x2_ASAP7_75t_R _12192_ (.A1(_03524_),
    .A2(_03880_),
    .B(_04921_),
    .C(_00422_),
    .Y(_05304_));
 AO21x1_ASAP7_75t_R _12193_ (.A1(_00421_),
    .A2(_03879_),
    .B(_05304_),
    .Y(_05305_));
 AND2x2_ASAP7_75t_R _12194_ (.A(_00423_),
    .B(_03805_),
    .Y(_05306_));
 AO221x1_ASAP7_75t_R _12195_ (.A1(_00424_),
    .A2(_03774_),
    .B1(_03803_),
    .B2(_03804_),
    .C(_05306_),
    .Y(_05307_));
 OA21x2_ASAP7_75t_R _12196_ (.A1(_03795_),
    .A2(_05305_),
    .B(_05307_),
    .Y(_05308_));
 AO21x1_ASAP7_75t_R _12197_ (.A1(_03792_),
    .A2(_05308_),
    .B(_03809_),
    .Y(_05309_));
 AND3x1_ASAP7_75t_R _12198_ (.A(_03376_),
    .B(_05215_),
    .C(_00420_),
    .Y(_05310_));
 AO21x1_ASAP7_75t_R _12199_ (.A1(_00419_),
    .A2(_04434_),
    .B(_05310_),
    .Y(_05311_));
 AO32x1_ASAP7_75t_R _12200_ (.A1(_03822_),
    .A2(_04587_),
    .A3(_05311_),
    .B1(_03703_),
    .B2(_00417_),
    .Y(_05312_));
 AND3x1_ASAP7_75t_R _12201_ (.A(_00418_),
    .B(_03814_),
    .C(_03889_),
    .Y(_05313_));
 OA21x2_ASAP7_75t_R _12202_ (.A1(_05312_),
    .A2(_05313_),
    .B(_04915_),
    .Y(_05314_));
 AND2x2_ASAP7_75t_R _12203_ (.A(_04938_),
    .B(_00430_),
    .Y(_05315_));
 AO21x1_ASAP7_75t_R _12204_ (.A1(_04937_),
    .A2(_00426_),
    .B(_05315_),
    .Y(_05316_));
 AO22x1_ASAP7_75t_R _12205_ (.A1(_00429_),
    .A2(_05221_),
    .B1(_05316_),
    .B2(_03845_),
    .Y(_05317_));
 NAND2x1_ASAP7_75t_R _12206_ (.A(_04053_),
    .B(_05317_),
    .Y(_05318_));
 AO21x1_ASAP7_75t_R _12207_ (.A1(_05218_),
    .A2(_05318_),
    .B(_05227_),
    .Y(_05319_));
 NAND2x1_ASAP7_75t_R _12208_ (.A(_00425_),
    .B(_03811_),
    .Y(_05320_));
 AND3x1_ASAP7_75t_R _12209_ (.A(_00427_),
    .B(_03804_),
    .C(_03831_),
    .Y(_05321_));
 AOI221x1_ASAP7_75t_R _12210_ (.A1(_00432_),
    .A2(_05230_),
    .B1(_04476_),
    .B2(_00431_),
    .C(_05321_),
    .Y(_05322_));
 AOI21x1_ASAP7_75t_R _12211_ (.A1(_00428_),
    .A2(_05233_),
    .B(_04792_),
    .Y(_05323_));
 AOI221x1_ASAP7_75t_R _12212_ (.A1(_05319_),
    .A2(_05320_),
    .B1(_05322_),
    .B2(_05323_),
    .C(_05235_),
    .Y(_05324_));
 AND3x1_ASAP7_75t_R _12213_ (.A(_03797_),
    .B(_03798_),
    .C(_00408_),
    .Y(_05325_));
 AO21x1_ASAP7_75t_R _12214_ (.A1(_00407_),
    .A2(_03796_),
    .B(_05325_),
    .Y(_05326_));
 AND3x1_ASAP7_75t_R _12215_ (.A(_03797_),
    .B(_03798_),
    .C(_00406_),
    .Y(_05327_));
 AO21x1_ASAP7_75t_R _12216_ (.A1(_00405_),
    .A2(_03796_),
    .B(_05327_),
    .Y(_05328_));
 AO32x2_ASAP7_75t_R _12217_ (.A1(_03852_),
    .A2(_04920_),
    .A3(_05326_),
    .B1(_05328_),
    .B2(_03721_),
    .Y(_05329_));
 INVx2_ASAP7_75t_R _12218_ (.A(_00409_),
    .Y(_05330_));
 BUFx10_ASAP7_75t_R _12219_ (.A(_04609_),
    .Y(_05331_));
 BUFx10_ASAP7_75t_R _12220_ (.A(_04610_),
    .Y(_05332_));
 AND2x2_ASAP7_75t_R _12221_ (.A(_05332_),
    .B(_00414_),
    .Y(_05333_));
 AO21x1_ASAP7_75t_R _12222_ (.A1(_05331_),
    .A2(_00410_),
    .B(_05333_),
    .Y(_05334_));
 AOI22x1_ASAP7_75t_R _12223_ (.A1(_00413_),
    .A2(_04936_),
    .B1(_05334_),
    .B2(_04930_),
    .Y(_05335_));
 OA211x2_ASAP7_75t_R _12224_ (.A1(_04935_),
    .A2(_05335_),
    .B(_03803_),
    .C(_03804_),
    .Y(_05336_));
 OAI22x1_ASAP7_75t_R _12225_ (.A1(_05330_),
    .A2(_04934_),
    .B1(_05336_),
    .B2(_04165_),
    .Y(_05337_));
 OA22x2_ASAP7_75t_R _12226_ (.A1(_00411_),
    .A2(_03690_),
    .B1(_04945_),
    .B2(_00416_),
    .Y(_05338_));
 OA22x2_ASAP7_75t_R _12227_ (.A1(_00412_),
    .A2(_04949_),
    .B1(_05338_),
    .B2(_03776_),
    .Y(_05339_));
 OA211x2_ASAP7_75t_R _12228_ (.A1(_00415_),
    .A2(_04944_),
    .B(_05339_),
    .C(_03868_),
    .Y(_05340_));
 AND2x2_ASAP7_75t_R _12229_ (.A(_05337_),
    .B(_05340_),
    .Y(_05341_));
 OA33x2_ASAP7_75t_R _12230_ (.A1(_05309_),
    .A2(_05314_),
    .A3(_05324_),
    .B1(_05329_),
    .B2(_05341_),
    .B3(_04452_),
    .Y(_05342_));
 AND3x1_ASAP7_75t_R _12231_ (.A(_03377_),
    .B(_04624_),
    .C(_00404_),
    .Y(_05343_));
 AO21x1_ASAP7_75t_R _12232_ (.A1(_00403_),
    .A2(_04623_),
    .B(_05343_),
    .Y(_05344_));
 AO222x2_ASAP7_75t_R _12233_ (.A1(_00401_),
    .A2(_04622_),
    .B1(_03901_),
    .B2(_05344_),
    .C1(_04629_),
    .C2(_00402_),
    .Y(_05345_));
 NOR2x2_ASAP7_75t_R _12234_ (.A(_05342_),
    .B(_05345_),
    .Y(_10007_));
 INVx3_ASAP7_75t_R _12235_ (.A(_10007_),
    .Y(_10009_));
 BUFx4f_ASAP7_75t_R _12236_ (.A(_03542_),
    .Y(_05346_));
 BUFx3_ASAP7_75t_R _12237_ (.A(_04175_),
    .Y(_05347_));
 AO32x1_ASAP7_75t_R _12238_ (.A1(_04171_),
    .A2(_04172_),
    .A3(_03905_),
    .B1(_03651_),
    .B2(_04848_),
    .Y(_05348_));
 OA21x2_ASAP7_75t_R _12239_ (.A1(_05347_),
    .A2(_05348_),
    .B(_04168_),
    .Y(_05349_));
 AO21x1_ASAP7_75t_R _12240_ (.A1(_04848_),
    .A2(_03905_),
    .B(_04176_),
    .Y(_05350_));
 AND3x1_ASAP7_75t_R _12241_ (.A(_04174_),
    .B(_04168_),
    .C(_05350_),
    .Y(_05351_));
 AO21x2_ASAP7_75t_R _12242_ (.A1(_05346_),
    .A2(_05349_),
    .B(_05351_),
    .Y(_10146_));
 AO22x1_ASAP7_75t_R _12243_ (.A1(_04656_),
    .A2(_00457_),
    .B1(_04069_),
    .B2(_00455_),
    .Y(_05352_));
 AND2x2_ASAP7_75t_R _12244_ (.A(_03926_),
    .B(_00456_),
    .Y(_05353_));
 AO21x1_ASAP7_75t_R _12245_ (.A1(_04114_),
    .A2(_00454_),
    .B(_05353_),
    .Y(_05354_));
 AO221x1_ASAP7_75t_R _12246_ (.A1(_04504_),
    .A2(_00454_),
    .B1(_05354_),
    .B2(_04080_),
    .C(_04280_),
    .Y(_05355_));
 AO21x1_ASAP7_75t_R _12247_ (.A1(_04066_),
    .A2(_05352_),
    .B(_05355_),
    .Y(_05356_));
 AND2x2_ASAP7_75t_R _12248_ (.A(_03975_),
    .B(_00464_),
    .Y(_05357_));
 AO21x1_ASAP7_75t_R _12249_ (.A1(_04085_),
    .A2(_00462_),
    .B(_05357_),
    .Y(_05358_));
 AO21x1_ASAP7_75t_R _12250_ (.A1(_00465_),
    .A2(_04091_),
    .B(_04009_),
    .Y(_05359_));
 AO221x1_ASAP7_75t_R _12251_ (.A1(_00463_),
    .A2(_04083_),
    .B1(_05358_),
    .B2(_04089_),
    .C(_05359_),
    .Y(_05360_));
 AO21x1_ASAP7_75t_R _12252_ (.A1(_05356_),
    .A2(_05360_),
    .B(_04095_),
    .Y(_05361_));
 AND3x1_ASAP7_75t_R _12253_ (.A(_04308_),
    .B(_04656_),
    .C(_00461_),
    .Y(_05362_));
 AND2x2_ASAP7_75t_R _12254_ (.A(_04018_),
    .B(_00460_),
    .Y(_05363_));
 AO21x1_ASAP7_75t_R _12255_ (.A1(_04521_),
    .A2(_00458_),
    .B(_05363_),
    .Y(_05364_));
 AO32x1_ASAP7_75t_R _12256_ (.A1(_04085_),
    .A2(_00459_),
    .A3(_04102_),
    .B1(_05364_),
    .B2(_04136_),
    .Y(_05365_));
 OR3x1_ASAP7_75t_R _12257_ (.A(_04099_),
    .B(_05362_),
    .C(_05365_),
    .Y(_05366_));
 AND2x2_ASAP7_75t_R _12258_ (.A(_04544_),
    .B(_00452_),
    .Y(_05367_));
 AO21x1_ASAP7_75t_R _12259_ (.A1(_04084_),
    .A2(_00450_),
    .B(_05367_),
    .Y(_05368_));
 AO32x1_ASAP7_75t_R _12260_ (.A1(_04074_),
    .A2(_00451_),
    .A3(_04102_),
    .B1(_05368_),
    .B2(_04136_),
    .Y(_05369_));
 AO221x1_ASAP7_75t_R _12261_ (.A1(_04112_),
    .A2(_04060_),
    .B1(_00453_),
    .B2(_04091_),
    .C(_05369_),
    .Y(_05370_));
 AO21x1_ASAP7_75t_R _12262_ (.A1(_05366_),
    .A2(_05370_),
    .B(_04120_),
    .Y(_05371_));
 AO21x2_ASAP7_75t_R _12263_ (.A1(_05361_),
    .A2(_05371_),
    .B(_04122_),
    .Y(_05372_));
 AND2x2_ASAP7_75t_R _12264_ (.A(_04127_),
    .B(_00449_),
    .Y(_05373_));
 AO21x1_ASAP7_75t_R _12265_ (.A1(_04126_),
    .A2(_00448_),
    .B(_05373_),
    .Y(_05374_));
 AND3x1_ASAP7_75t_R _12266_ (.A(_04138_),
    .B(_03380_),
    .C(_00447_),
    .Y(_05375_));
 AO21x1_ASAP7_75t_R _12267_ (.A1(_00446_),
    .A2(_04141_),
    .B(_05375_),
    .Y(_05376_));
 AO221x1_ASAP7_75t_R _12268_ (.A1(_04067_),
    .A2(_05374_),
    .B1(_05376_),
    .B2(_04145_),
    .C(_04008_),
    .Y(_05377_));
 AND2x2_ASAP7_75t_R _12269_ (.A(_04987_),
    .B(_00444_),
    .Y(_05378_));
 AO21x1_ASAP7_75t_R _12270_ (.A1(_04074_),
    .A2(_00442_),
    .B(_05378_),
    .Y(_05379_));
 AO21x1_ASAP7_75t_R _12271_ (.A1(_00443_),
    .A2(_04083_),
    .B(_04032_),
    .Y(_05380_));
 AO221x1_ASAP7_75t_R _12272_ (.A1(_00445_),
    .A2(_04091_),
    .B1(_05379_),
    .B2(_04089_),
    .C(_05380_),
    .Y(_05381_));
 AND3x1_ASAP7_75t_R _12273_ (.A(_04157_),
    .B(_05377_),
    .C(_05381_),
    .Y(_05382_));
 AND2x2_ASAP7_75t_R _12274_ (.A(_04307_),
    .B(_00437_),
    .Y(_05383_));
 AO21x1_ASAP7_75t_R _12275_ (.A1(_03951_),
    .A2(_00436_),
    .B(_05383_),
    .Y(_05384_));
 AO21x1_ASAP7_75t_R _12276_ (.A1(_04656_),
    .A2(_05384_),
    .B(_04119_),
    .Y(_05385_));
 AO22x1_ASAP7_75t_R _12277_ (.A1(_04531_),
    .A2(_00434_),
    .B1(_00435_),
    .B2(_04522_),
    .Y(_05386_));
 AO22x1_ASAP7_75t_R _12278_ (.A1(_04504_),
    .A2(_00434_),
    .B1(_05386_),
    .B2(_04085_),
    .Y(_05387_));
 AO21x1_ASAP7_75t_R _12279_ (.A1(_04060_),
    .A2(_05385_),
    .B(_05387_),
    .Y(_05388_));
 AND2x2_ASAP7_75t_R _12280_ (.A(_04127_),
    .B(_00441_),
    .Y(_05389_));
 AO21x1_ASAP7_75t_R _12281_ (.A1(_04126_),
    .A2(_00440_),
    .B(_05389_),
    .Y(_05390_));
 AND3x1_ASAP7_75t_R _12282_ (.A(_04138_),
    .B(_03380_),
    .C(_00439_),
    .Y(_05391_));
 AO21x1_ASAP7_75t_R _12283_ (.A1(_00438_),
    .A2(_04141_),
    .B(_05391_),
    .Y(_05392_));
 AO221x1_ASAP7_75t_R _12284_ (.A1(_04067_),
    .A2(_05390_),
    .B1(_05392_),
    .B2(_04145_),
    .C(_04008_),
    .Y(_05393_));
 AND3x1_ASAP7_75t_R _12285_ (.A(_04099_),
    .B(_05388_),
    .C(_05393_),
    .Y(_05394_));
 OR3x1_ASAP7_75t_R _12286_ (.A(_04124_),
    .B(_05382_),
    .C(_05394_),
    .Y(_05395_));
 AOI21x1_ASAP7_75t_R _12287_ (.A1(_05372_),
    .A2(_05395_),
    .B(_04565_),
    .Y(_05396_));
 OR2x2_ASAP7_75t_R _12288_ (.A(_04162_),
    .B(_05396_),
    .Y(_05397_));
 OA21x2_ASAP7_75t_R _12289_ (.A1(_04065_),
    .A2(_10146_),
    .B(_05397_),
    .Y(_05398_));
 XNOR2x1_ASAP7_75t_R _12290_ (.B(_05398_),
    .Y(_10013_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _12291_ (.A(_10013_),
    .Y(_10015_));
 AND3x1_ASAP7_75t_R _12292_ (.A(_04455_),
    .B(_04597_),
    .C(_00453_),
    .Y(_05399_));
 AO21x1_ASAP7_75t_R _12293_ (.A1(_00452_),
    .A2(_03782_),
    .B(_05399_),
    .Y(_05400_));
 AO32x1_ASAP7_75t_R _12294_ (.A1(_03655_),
    .A2(_04587_),
    .A3(_05400_),
    .B1(_03703_),
    .B2(_00450_),
    .Y(_05401_));
 AND2x2_ASAP7_75t_R _12295_ (.A(_04915_),
    .B(_05401_),
    .Y(_05402_));
 BUFx10_ASAP7_75t_R _12296_ (.A(_03791_),
    .Y(_05403_));
 AND2x2_ASAP7_75t_R _12297_ (.A(_00455_),
    .B(_04591_),
    .Y(_05404_));
 AND2x2_ASAP7_75t_R _12298_ (.A(_00454_),
    .B(_03878_),
    .Y(_05405_));
 OR3x1_ASAP7_75t_R _12299_ (.A(_03794_),
    .B(_05404_),
    .C(_05405_),
    .Y(_05406_));
 AND2x2_ASAP7_75t_R _12300_ (.A(_00456_),
    .B(_03711_),
    .Y(_05407_));
 AO221x1_ASAP7_75t_R _12301_ (.A1(_00457_),
    .A2(_03887_),
    .B1(_03803_),
    .B2(_03837_),
    .C(_05407_),
    .Y(_05408_));
 AND2x2_ASAP7_75t_R _12302_ (.A(_03701_),
    .B(_04628_),
    .Y(_05409_));
 AO32x1_ASAP7_75t_R _12303_ (.A1(_05403_),
    .A2(_05406_),
    .A3(_05408_),
    .B1(_05409_),
    .B2(_00451_),
    .Y(_05410_));
 AND3x1_ASAP7_75t_R _12304_ (.A(_04916_),
    .B(_04584_),
    .C(_00461_),
    .Y(_05411_));
 AO21x1_ASAP7_75t_R _12305_ (.A1(_00460_),
    .A2(_03891_),
    .B(_05411_),
    .Y(_05412_));
 AND2x2_ASAP7_75t_R _12306_ (.A(_00464_),
    .B(_03890_),
    .Y(_05413_));
 AO221x1_ASAP7_75t_R _12307_ (.A1(_00465_),
    .A2(_04921_),
    .B1(_03874_),
    .B2(_03861_),
    .C(_05413_),
    .Y(_05414_));
 OA21x2_ASAP7_75t_R _12308_ (.A1(_04602_),
    .A2(_05412_),
    .B(_05414_),
    .Y(_05415_));
 INVx1_ASAP7_75t_R _12309_ (.A(_00458_),
    .Y(_05416_));
 BUFx10_ASAP7_75t_R _12310_ (.A(_04811_),
    .Y(_05417_));
 AND2x2_ASAP7_75t_R _12311_ (.A(_03610_),
    .B(_00463_),
    .Y(_05418_));
 AO21x1_ASAP7_75t_R _12312_ (.A1(_04831_),
    .A2(_00459_),
    .B(_05418_),
    .Y(_05419_));
 AOI22x1_ASAP7_75t_R _12313_ (.A1(_00462_),
    .A2(_05221_),
    .B1(_05419_),
    .B2(_05215_),
    .Y(_05420_));
 OA211x2_ASAP7_75t_R _12314_ (.A1(_05417_),
    .A2(_05420_),
    .B(_03888_),
    .C(_03705_),
    .Y(_05421_));
 OAI22x1_ASAP7_75t_R _12315_ (.A1(_05416_),
    .A2(_04799_),
    .B1(_05421_),
    .B2(_05227_),
    .Y(_05422_));
 OA211x2_ASAP7_75t_R _12316_ (.A1(_04792_),
    .A2(_05415_),
    .B(_05422_),
    .C(_03850_),
    .Y(_05423_));
 OR4x2_ASAP7_75t_R _12317_ (.A(_03809_),
    .B(_05402_),
    .C(_05410_),
    .D(_05423_),
    .Y(_05424_));
 AND3x1_ASAP7_75t_R _12318_ (.A(_03797_),
    .B(_04930_),
    .C(_00437_),
    .Y(_05425_));
 AO21x1_ASAP7_75t_R _12319_ (.A1(_00436_),
    .A2(_04929_),
    .B(_05425_),
    .Y(_05426_));
 AO222x2_ASAP7_75t_R _12320_ (.A1(_00434_),
    .A2(_04622_),
    .B1(_03901_),
    .B2(_05426_),
    .C1(_04629_),
    .C2(_00435_),
    .Y(_05427_));
 OR3x1_ASAP7_75t_R _12321_ (.A(_00438_),
    .B(_03814_),
    .C(_03794_),
    .Y(_05428_));
 OR2x2_ASAP7_75t_R _12322_ (.A(_00440_),
    .B(_03866_),
    .Y(_05429_));
 OR3x1_ASAP7_75t_R _12323_ (.A(_00439_),
    .B(_03780_),
    .C(_03765_),
    .Y(_05430_));
 AO21x1_ASAP7_75t_R _12324_ (.A1(_03829_),
    .A2(_04592_),
    .B(_00441_),
    .Y(_05431_));
 AO21x1_ASAP7_75t_R _12325_ (.A1(_05430_),
    .A2(_05431_),
    .B(_03879_),
    .Y(_05432_));
 AND4x1_ASAP7_75t_R _12326_ (.A(_05403_),
    .B(_05428_),
    .C(_05429_),
    .D(_05432_),
    .Y(_05433_));
 AO21x1_ASAP7_75t_R _12327_ (.A1(_03639_),
    .A2(_03717_),
    .B(_00448_),
    .Y(_05434_));
 OA21x2_ASAP7_75t_R _12328_ (.A1(_00449_),
    .A2(_03714_),
    .B(_05434_),
    .Y(_05435_));
 OR3x1_ASAP7_75t_R _12329_ (.A(_00444_),
    .B(_03881_),
    .C(_04948_),
    .Y(_05436_));
 OA21x2_ASAP7_75t_R _12330_ (.A1(_03836_),
    .A2(_05434_),
    .B(_05436_),
    .Y(_05437_));
 OA211x2_ASAP7_75t_R _12331_ (.A1(_03707_),
    .A2(_05435_),
    .B(_05437_),
    .C(_03698_),
    .Y(_05438_));
 INVx2_ASAP7_75t_R _12332_ (.A(_00442_),
    .Y(_05439_));
 AND2x2_ASAP7_75t_R _12333_ (.A(_03610_),
    .B(_00447_),
    .Y(_05440_));
 AO21x1_ASAP7_75t_R _12334_ (.A1(_04831_),
    .A2(_00443_),
    .B(_05440_),
    .Y(_05441_));
 AOI22x1_ASAP7_75t_R _12335_ (.A1(_00446_),
    .A2(_05221_),
    .B1(_05441_),
    .B2(_05215_),
    .Y(_05442_));
 OA211x2_ASAP7_75t_R _12336_ (.A1(_05417_),
    .A2(_05442_),
    .B(_03888_),
    .C(_03705_),
    .Y(_05443_));
 OAI22x1_ASAP7_75t_R _12337_ (.A1(_05439_),
    .A2(_04799_),
    .B1(_05443_),
    .B2(_05227_),
    .Y(_05444_));
 OA211x2_ASAP7_75t_R _12338_ (.A1(_00445_),
    .A2(_04949_),
    .B(_05438_),
    .C(_05444_),
    .Y(_05445_));
 OR4x2_ASAP7_75t_R _12339_ (.A(_04452_),
    .B(_05427_),
    .C(_05433_),
    .D(_05445_),
    .Y(_05446_));
 NAND2x2_ASAP7_75t_R _12340_ (.A(_05424_),
    .B(_05446_),
    .Y(_10012_));
 INVx4_ASAP7_75t_R _12341_ (.A(_10012_),
    .Y(_10014_));
 AO32x1_ASAP7_75t_R _12342_ (.A1(_04171_),
    .A2(_04172_),
    .A3(_03651_),
    .B1(_03872_),
    .B2(_04848_),
    .Y(_05447_));
 OA21x2_ASAP7_75t_R _12343_ (.A1(_05347_),
    .A2(_05447_),
    .B(_04167_),
    .Y(_05448_));
 AND2x2_ASAP7_75t_R _12344_ (.A(_05346_),
    .B(_05448_),
    .Y(_05449_));
 AO21x2_ASAP7_75t_R _12345_ (.A1(_04174_),
    .A2(_05349_),
    .B(_05449_),
    .Y(_10144_));
 AO22x1_ASAP7_75t_R _12346_ (.A1(_04255_),
    .A2(_00490_),
    .B1(_04632_),
    .B2(_00488_),
    .Y(_05450_));
 AND2x2_ASAP7_75t_R _12347_ (.A(_03925_),
    .B(_00489_),
    .Y(_05451_));
 AO21x1_ASAP7_75t_R _12348_ (.A1(_04103_),
    .A2(_00487_),
    .B(_05451_),
    .Y(_05452_));
 AO221x1_ASAP7_75t_R _12349_ (.A1(_04071_),
    .A2(_00487_),
    .B1(_05452_),
    .B2(_04079_),
    .C(_03920_),
    .Y(_05453_));
 AO21x1_ASAP7_75t_R _12350_ (.A1(_04066_),
    .A2(_05450_),
    .B(_05453_),
    .Y(_05454_));
 AND2x2_ASAP7_75t_R _12351_ (.A(_04544_),
    .B(_00497_),
    .Y(_05455_));
 AO21x1_ASAP7_75t_R _12352_ (.A1(_04521_),
    .A2(_00495_),
    .B(_05455_),
    .Y(_05456_));
 AO21x1_ASAP7_75t_R _12353_ (.A1(_00498_),
    .A2(_04262_),
    .B(_04009_),
    .Y(_05457_));
 AO221x1_ASAP7_75t_R _12354_ (.A1(_00496_),
    .A2(_04083_),
    .B1(_05456_),
    .B2(_04136_),
    .C(_05457_),
    .Y(_05458_));
 AO21x1_ASAP7_75t_R _12355_ (.A1(_05454_),
    .A2(_05458_),
    .B(_04095_),
    .Y(_05459_));
 AND3x1_ASAP7_75t_R _12356_ (.A(_04016_),
    .B(_03975_),
    .C(_00494_),
    .Y(_05460_));
 AND2x2_ASAP7_75t_R _12357_ (.A(_03925_),
    .B(_00493_),
    .Y(_05461_));
 AO21x1_ASAP7_75t_R _12358_ (.A1(_04113_),
    .A2(_00491_),
    .B(_05461_),
    .Y(_05462_));
 AO32x1_ASAP7_75t_R _12359_ (.A1(_04084_),
    .A2(_00492_),
    .A3(_04522_),
    .B1(_05462_),
    .B2(_04531_),
    .Y(_05463_));
 OR3x1_ASAP7_75t_R _12360_ (.A(_04098_),
    .B(_05460_),
    .C(_05463_),
    .Y(_05464_));
 AND2x2_ASAP7_75t_R _12361_ (.A(_04017_),
    .B(_00485_),
    .Y(_05465_));
 AO21x1_ASAP7_75t_R _12362_ (.A1(_04520_),
    .A2(_00483_),
    .B(_05465_),
    .Y(_05466_));
 AO32x1_ASAP7_75t_R _12363_ (.A1(_04084_),
    .A2(_00484_),
    .A3(_04522_),
    .B1(_05466_),
    .B2(_04556_),
    .Y(_05467_));
 AO221x1_ASAP7_75t_R _12364_ (.A1(_04112_),
    .A2(_03381_),
    .B1(_00486_),
    .B2(_03962_),
    .C(_05467_),
    .Y(_05468_));
 AO21x1_ASAP7_75t_R _12365_ (.A1(_05464_),
    .A2(_05468_),
    .B(_04120_),
    .Y(_05469_));
 AOI21x1_ASAP7_75t_R _12366_ (.A1(_05459_),
    .A2(_05469_),
    .B(_04122_),
    .Y(_05470_));
 AND2x2_ASAP7_75t_R _12367_ (.A(_04034_),
    .B(_00470_),
    .Y(_05471_));
 AO21x1_ASAP7_75t_R _12368_ (.A1(_03951_),
    .A2(_00469_),
    .B(_05471_),
    .Y(_05472_));
 AO21x1_ASAP7_75t_R _12369_ (.A1(_04656_),
    .A2(_05472_),
    .B(_04119_),
    .Y(_05473_));
 AO22x1_ASAP7_75t_R _12370_ (.A1(_04647_),
    .A2(_00467_),
    .B1(_00468_),
    .B2(_04522_),
    .Y(_05474_));
 AO22x1_ASAP7_75t_R _12371_ (.A1(_04072_),
    .A2(_00467_),
    .B1(_05474_),
    .B2(_04085_),
    .Y(_05475_));
 AO21x1_ASAP7_75t_R _12372_ (.A1(_04060_),
    .A2(_05473_),
    .B(_05475_),
    .Y(_05476_));
 AND2x2_ASAP7_75t_R _12373_ (.A(_03942_),
    .B(_00474_),
    .Y(_05477_));
 AO21x1_ASAP7_75t_R _12374_ (.A1(_04671_),
    .A2(_00473_),
    .B(_05477_),
    .Y(_05478_));
 AND3x1_ASAP7_75t_R _12375_ (.A(_04666_),
    .B(_04559_),
    .C(_00472_),
    .Y(_05479_));
 AO21x1_ASAP7_75t_R _12376_ (.A1(_00471_),
    .A2(_04292_),
    .B(_05479_),
    .Y(_05480_));
 AO221x1_ASAP7_75t_R _12377_ (.A1(_04289_),
    .A2(_05478_),
    .B1(_05480_),
    .B2(_04295_),
    .C(_04094_),
    .Y(_05481_));
 AND2x2_ASAP7_75t_R _12378_ (.A(_04514_),
    .B(_05481_),
    .Y(_05482_));
 AND2x2_ASAP7_75t_R _12379_ (.A(_04666_),
    .B(_00482_),
    .Y(_05483_));
 AO21x1_ASAP7_75t_R _12380_ (.A1(_04671_),
    .A2(_00481_),
    .B(_05483_),
    .Y(_05484_));
 AND3x1_ASAP7_75t_R _12381_ (.A(_04015_),
    .B(_04559_),
    .C(_00480_),
    .Y(_05485_));
 AO21x1_ASAP7_75t_R _12382_ (.A1(_00479_),
    .A2(_04535_),
    .B(_05485_),
    .Y(_05486_));
 AO221x1_ASAP7_75t_R _12383_ (.A1(_04502_),
    .A2(_05484_),
    .B1(_05486_),
    .B2(_04295_),
    .C(_04094_),
    .Y(_05487_));
 AND2x2_ASAP7_75t_R _12384_ (.A(_03974_),
    .B(_00477_),
    .Y(_05488_));
 AO21x1_ASAP7_75t_R _12385_ (.A1(_03992_),
    .A2(_00475_),
    .B(_05488_),
    .Y(_05489_));
 AO21x1_ASAP7_75t_R _12386_ (.A1(_00476_),
    .A2(_03964_),
    .B(_03981_),
    .Y(_05490_));
 AO221x1_ASAP7_75t_R _12387_ (.A1(_00478_),
    .A2(_03962_),
    .B1(_05489_),
    .B2(_04126_),
    .C(_05490_),
    .Y(_05491_));
 AND3x1_ASAP7_75t_R _12388_ (.A(_04157_),
    .B(_05487_),
    .C(_05491_),
    .Y(_05492_));
 AOI211x1_ASAP7_75t_R _12389_ (.A1(_05476_),
    .A2(_05482_),
    .B(_04124_),
    .C(_05492_),
    .Y(_05493_));
 OA21x2_ASAP7_75t_R _12390_ (.A1(_05470_),
    .A2(_05493_),
    .B(_03447_),
    .Y(_05494_));
 OR2x2_ASAP7_75t_R _12391_ (.A(_04162_),
    .B(_05494_),
    .Y(_05495_));
 OA21x2_ASAP7_75t_R _12392_ (.A1(_04065_),
    .A2(_10144_),
    .B(_05495_),
    .Y(_05496_));
 XNOR2x1_ASAP7_75t_R _12393_ (.B(_05496_),
    .Y(_10018_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _12394_ (.A(_10018_),
    .Y(_10020_));
 AND2x2_ASAP7_75t_R _12395_ (.A(_04591_),
    .B(_04727_),
    .Y(_05497_));
 AO21x1_ASAP7_75t_R _12396_ (.A1(_00488_),
    .A2(_05497_),
    .B(_04499_),
    .Y(_05498_));
 AND3x1_ASAP7_75t_R _12397_ (.A(_03843_),
    .B(_04460_),
    .C(_00490_),
    .Y(_05499_));
 AO21x1_ASAP7_75t_R _12398_ (.A1(_00489_),
    .A2(_04236_),
    .B(_05499_),
    .Y(_05500_));
 AO32x1_ASAP7_75t_R _12399_ (.A1(_00487_),
    .A2(_03829_),
    .A3(_03648_),
    .B1(_05500_),
    .B2(_03794_),
    .Y(_05501_));
 INVx2_ASAP7_75t_R _12400_ (.A(_00485_),
    .Y(_05502_));
 INVx1_ASAP7_75t_R _12401_ (.A(_00484_),
    .Y(_05503_));
 NAND2x1_ASAP7_75t_R _12402_ (.A(_03636_),
    .B(_00486_),
    .Y(_05504_));
 OA211x2_ASAP7_75t_R _12403_ (.A1(_03897_),
    .A2(_05503_),
    .B(_05504_),
    .C(_03672_),
    .Y(_05505_));
 AOI21x1_ASAP7_75t_R _12404_ (.A1(_05502_),
    .A2(_04442_),
    .B(_05505_),
    .Y(_05506_));
 OA211x2_ASAP7_75t_R _12405_ (.A1(_04811_),
    .A2(_05506_),
    .B(_03771_),
    .C(_03828_),
    .Y(_05507_));
 OA22x2_ASAP7_75t_R _12406_ (.A1(_00483_),
    .A2(_03759_),
    .B1(_05507_),
    .B2(_03785_),
    .Y(_05508_));
 AO21x1_ASAP7_75t_R _12407_ (.A1(_03791_),
    .A2(_05501_),
    .B(_05508_),
    .Y(_05509_));
 AND2x2_ASAP7_75t_R _12408_ (.A(_04592_),
    .B(_03698_),
    .Y(_05510_));
 AND3x1_ASAP7_75t_R _12409_ (.A(_03375_),
    .B(_04435_),
    .C(_00494_),
    .Y(_05511_));
 AO21x1_ASAP7_75t_R _12410_ (.A1(_00493_),
    .A2(_03781_),
    .B(_05511_),
    .Y(_05512_));
 AND2x2_ASAP7_75t_R _12411_ (.A(_00497_),
    .B(_03612_),
    .Y(_05513_));
 AO221x1_ASAP7_75t_R _12412_ (.A1(_00498_),
    .A2(_03881_),
    .B1(_03661_),
    .B2(_03860_),
    .C(_05513_),
    .Y(_05514_));
 OA211x2_ASAP7_75t_R _12413_ (.A1(_03871_),
    .A2(_05512_),
    .B(_05514_),
    .C(_03697_),
    .Y(_05515_));
 INVx1_ASAP7_75t_R _12414_ (.A(_00491_),
    .Y(_05516_));
 AND2x2_ASAP7_75t_R _12415_ (.A(_04610_),
    .B(_00496_),
    .Y(_05517_));
 AO21x1_ASAP7_75t_R _12416_ (.A1(_04457_),
    .A2(_00492_),
    .B(_05517_),
    .Y(_05518_));
 AOI22x1_ASAP7_75t_R _12417_ (.A1(_00495_),
    .A2(_04576_),
    .B1(_05518_),
    .B2(_03665_),
    .Y(_05519_));
 OA211x2_ASAP7_75t_R _12418_ (.A1(_03839_),
    .A2(_05519_),
    .B(_03775_),
    .C(_03737_),
    .Y(_05520_));
 OAI22x1_ASAP7_75t_R _12419_ (.A1(_05516_),
    .A2(_04575_),
    .B1(_05520_),
    .B2(_04164_),
    .Y(_05521_));
 OA21x2_ASAP7_75t_R _12420_ (.A1(_05510_),
    .A2(_05515_),
    .B(_05521_),
    .Y(_05522_));
 OR3x1_ASAP7_75t_R _12421_ (.A(_00471_),
    .B(_04591_),
    .C(_03794_),
    .Y(_05523_));
 OA211x2_ASAP7_75t_R _12422_ (.A1(_00473_),
    .A2(_03865_),
    .B(_03653_),
    .C(_04244_),
    .Y(_05524_));
 OR3x1_ASAP7_75t_R _12423_ (.A(_00472_),
    .B(_03606_),
    .C(_03765_),
    .Y(_05525_));
 AO21x1_ASAP7_75t_R _12424_ (.A1(_03737_),
    .A2(_03775_),
    .B(_00474_),
    .Y(_05526_));
 AO21x1_ASAP7_75t_R _12425_ (.A1(_05525_),
    .A2(_05526_),
    .B(_03586_),
    .Y(_05527_));
 AO32x2_ASAP7_75t_R _12426_ (.A1(_05523_),
    .A2(_05524_),
    .A3(_05527_),
    .B1(_03905_),
    .B2(_03742_),
    .Y(_05528_));
 OA31x2_ASAP7_75t_R _12427_ (.A1(_05498_),
    .A2(_05509_),
    .A3(_05522_),
    .B1(_05528_),
    .Y(_05529_));
 INVx2_ASAP7_75t_R _12428_ (.A(_00475_),
    .Y(_05530_));
 AND2x2_ASAP7_75t_R _12429_ (.A(_04938_),
    .B(_00480_),
    .Y(_05531_));
 AO21x1_ASAP7_75t_R _12430_ (.A1(_04937_),
    .A2(_00476_),
    .B(_05531_),
    .Y(_05532_));
 AOI22x1_ASAP7_75t_R _12431_ (.A1(_00479_),
    .A2(_05221_),
    .B1(_05532_),
    .B2(_03845_),
    .Y(_05533_));
 OA21x2_ASAP7_75t_R _12432_ (.A1(_04935_),
    .A2(_05533_),
    .B(_03825_),
    .Y(_05534_));
 OAI22x1_ASAP7_75t_R _12433_ (.A1(_05530_),
    .A2(_04934_),
    .B1(_05534_),
    .B2(_03786_),
    .Y(_05535_));
 AND3x1_ASAP7_75t_R _12434_ (.A(_00477_),
    .B(_03737_),
    .C(_03735_),
    .Y(_05536_));
 AO21x1_ASAP7_75t_R _12435_ (.A1(_00481_),
    .A2(_03871_),
    .B(_05536_),
    .Y(_05537_));
 AO221x1_ASAP7_75t_R _12436_ (.A1(_00482_),
    .A2(_04198_),
    .B1(_03833_),
    .B2(_00478_),
    .C(_03659_),
    .Y(_05538_));
 AO21x1_ASAP7_75t_R _12437_ (.A1(_04929_),
    .A2(_05537_),
    .B(_05538_),
    .Y(_05539_));
 OA21x2_ASAP7_75t_R _12438_ (.A1(_00469_),
    .A2(_03865_),
    .B(_04193_),
    .Y(_05540_));
 OR2x2_ASAP7_75t_R _12439_ (.A(_03785_),
    .B(_05540_),
    .Y(_05541_));
 AND2x2_ASAP7_75t_R _12440_ (.A(_00468_),
    .B(_03659_),
    .Y(_05542_));
 AND2x2_ASAP7_75t_R _12441_ (.A(_00470_),
    .B(_03733_),
    .Y(_05543_));
 OR3x1_ASAP7_75t_R _12442_ (.A(_03879_),
    .B(_05542_),
    .C(_05543_),
    .Y(_05544_));
 AO32x2_ASAP7_75t_R _12443_ (.A1(_04839_),
    .A2(_05535_),
    .A3(_05539_),
    .B1(_05541_),
    .B2(_05544_),
    .Y(_05545_));
 OR2x2_ASAP7_75t_R _12444_ (.A(_05529_),
    .B(_05545_),
    .Y(_05546_));
 BUFx4f_ASAP7_75t_R _12445_ (.A(_05546_),
    .Y(_10019_));
 BUFx4f_ASAP7_75t_R _12446_ (.A(_04059_),
    .Y(_05547_));
 AO32x1_ASAP7_75t_R _12447_ (.A1(_04171_),
    .A2(_04172_),
    .A3(_03872_),
    .B1(_03852_),
    .B2(_04848_),
    .Y(_05548_));
 OA21x2_ASAP7_75t_R _12448_ (.A1(_04175_),
    .A2(_05548_),
    .B(_04167_),
    .Y(_05549_));
 AND2x2_ASAP7_75t_R _12449_ (.A(_05346_),
    .B(_05549_),
    .Y(_05550_));
 AO21x2_ASAP7_75t_R _12450_ (.A1(_04174_),
    .A2(_05448_),
    .B(_05550_),
    .Y(_10142_));
 AO22x1_ASAP7_75t_R _12451_ (.A1(_04643_),
    .A2(_00523_),
    .B1(_04632_),
    .B2(_00521_),
    .Y(_05551_));
 AND2x2_ASAP7_75t_R _12452_ (.A(_03925_),
    .B(_00522_),
    .Y(_05552_));
 AO21x1_ASAP7_75t_R _12453_ (.A1(_04113_),
    .A2(_00520_),
    .B(_05552_),
    .Y(_05553_));
 AO221x1_ASAP7_75t_R _12454_ (.A1(_03984_),
    .A2(_00520_),
    .B1(_05553_),
    .B2(_04531_),
    .C(_03920_),
    .Y(_05554_));
 AO21x1_ASAP7_75t_R _12455_ (.A1(_04066_),
    .A2(_05551_),
    .B(_05554_),
    .Y(_05555_));
 AND2x2_ASAP7_75t_R _12456_ (.A(_04544_),
    .B(_00530_),
    .Y(_05556_));
 AO21x1_ASAP7_75t_R _12457_ (.A1(_04084_),
    .A2(_00528_),
    .B(_05556_),
    .Y(_05557_));
 AO21x1_ASAP7_75t_R _12458_ (.A1(_00531_),
    .A2(_04090_),
    .B(_04009_),
    .Y(_05558_));
 AO221x1_ASAP7_75t_R _12459_ (.A1(_00529_),
    .A2(_04983_),
    .B1(_05557_),
    .B2(_04136_),
    .C(_05558_),
    .Y(_05559_));
 AO21x1_ASAP7_75t_R _12460_ (.A1(_05555_),
    .A2(_05559_),
    .B(_04095_),
    .Y(_05560_));
 AND3x1_ASAP7_75t_R _12461_ (.A(_04138_),
    .B(_04270_),
    .C(_00527_),
    .Y(_05561_));
 AND2x2_ASAP7_75t_R _12462_ (.A(_04017_),
    .B(_00526_),
    .Y(_05562_));
 AO21x1_ASAP7_75t_R _12463_ (.A1(_04520_),
    .A2(_00524_),
    .B(_05562_),
    .Y(_05563_));
 AO32x1_ASAP7_75t_R _12464_ (.A1(_03992_),
    .A2(_00525_),
    .A3(_05073_),
    .B1(_05563_),
    .B2(_04671_),
    .Y(_05564_));
 OR3x1_ASAP7_75t_R _12465_ (.A(_04098_),
    .B(_05561_),
    .C(_05564_),
    .Y(_05565_));
 AND2x2_ASAP7_75t_R _12466_ (.A(_04043_),
    .B(_00518_),
    .Y(_05566_));
 AO21x1_ASAP7_75t_R _12467_ (.A1(_04520_),
    .A2(_00516_),
    .B(_05566_),
    .Y(_05567_));
 AO32x1_ASAP7_75t_R _12468_ (.A1(_04276_),
    .A2(_00517_),
    .A3(_05073_),
    .B1(_05567_),
    .B2(_04671_),
    .Y(_05568_));
 AO221x1_ASAP7_75t_R _12469_ (.A1(_04112_),
    .A2(_03972_),
    .B1(_00519_),
    .B2(_03962_),
    .C(_05568_),
    .Y(_05569_));
 AO21x1_ASAP7_75t_R _12470_ (.A1(_05565_),
    .A2(_05569_),
    .B(_04131_),
    .Y(_05570_));
 AO21x2_ASAP7_75t_R _12471_ (.A1(_05560_),
    .A2(_05570_),
    .B(_03917_),
    .Y(_05571_));
 AND2x2_ASAP7_75t_R _12472_ (.A(_03933_),
    .B(_00515_),
    .Y(_05572_));
 AO21x1_ASAP7_75t_R _12473_ (.A1(_03930_),
    .A2(_00514_),
    .B(_05572_),
    .Y(_05573_));
 AND3x1_ASAP7_75t_R _12474_ (.A(_04137_),
    .B(_03943_),
    .C(_00513_),
    .Y(_05574_));
 AO21x1_ASAP7_75t_R _12475_ (.A1(_00512_),
    .A2(_03939_),
    .B(_05574_),
    .Y(_05575_));
 AO221x1_ASAP7_75t_R _12476_ (.A1(_03927_),
    .A2(_05573_),
    .B1(_05575_),
    .B2(_03938_),
    .C(_03947_),
    .Y(_05576_));
 AND2x2_ASAP7_75t_R _12477_ (.A(_03957_),
    .B(_00510_),
    .Y(_05577_));
 AO21x1_ASAP7_75t_R _12478_ (.A1(_04276_),
    .A2(_00508_),
    .B(_05577_),
    .Y(_05578_));
 AO21x1_ASAP7_75t_R _12479_ (.A1(_00509_),
    .A2(_03964_),
    .B(_03966_),
    .Y(_05579_));
 AO221x1_ASAP7_75t_R _12480_ (.A1(_00511_),
    .A2(_04262_),
    .B1(_05578_),
    .B2(_04265_),
    .C(_05579_),
    .Y(_05580_));
 AND3x1_ASAP7_75t_R _12481_ (.A(_04157_),
    .B(_05576_),
    .C(_05580_),
    .Y(_05581_));
 AND2x2_ASAP7_75t_R _12482_ (.A(_04403_),
    .B(_00503_),
    .Y(_05582_));
 AO21x1_ASAP7_75t_R _12483_ (.A1(_03986_),
    .A2(_00502_),
    .B(_05582_),
    .Y(_05583_));
 AO21x1_ASAP7_75t_R _12484_ (.A1(_04529_),
    .A2(_05583_),
    .B(_03966_),
    .Y(_05584_));
 AND2x2_ASAP7_75t_R _12485_ (.A(_03972_),
    .B(_05584_),
    .Y(_05585_));
 AO22x1_ASAP7_75t_R _12486_ (.A1(_04125_),
    .A2(_00500_),
    .B1(_00501_),
    .B2(_05073_),
    .Y(_05586_));
 AO22x2_ASAP7_75t_R _12487_ (.A1(_04504_),
    .A2(_00500_),
    .B1(_05586_),
    .B2(_04104_),
    .Y(_05587_));
 AND2x2_ASAP7_75t_R _12488_ (.A(_04033_),
    .B(_00507_),
    .Y(_05588_));
 AO21x1_ASAP7_75t_R _12489_ (.A1(_03950_),
    .A2(_00506_),
    .B(_05588_),
    .Y(_05589_));
 BUFx6f_ASAP7_75t_R _12490_ (.A(_03548_),
    .Y(_05590_));
 AND3x1_ASAP7_75t_R _12491_ (.A(_04033_),
    .B(_04314_),
    .C(_00505_),
    .Y(_05591_));
 AO21x1_ASAP7_75t_R _12492_ (.A1(_00504_),
    .A2(_05590_),
    .B(_05591_),
    .Y(_05592_));
 AO221x1_ASAP7_75t_R _12493_ (.A1(_03975_),
    .A2(_05589_),
    .B1(_05592_),
    .B2(_04995_),
    .C(_04541_),
    .Y(_05593_));
 OA211x2_ASAP7_75t_R _12494_ (.A1(_05585_),
    .A2(_05587_),
    .B(_05593_),
    .C(_04514_),
    .Y(_05594_));
 OR3x1_ASAP7_75t_R _12495_ (.A(_04763_),
    .B(_05581_),
    .C(_05594_),
    .Y(_05595_));
 AOI21x1_ASAP7_75t_R _12496_ (.A1(_05571_),
    .A2(_05595_),
    .B(_04565_),
    .Y(_05596_));
 OR2x2_ASAP7_75t_R _12497_ (.A(_04162_),
    .B(_05596_),
    .Y(_05597_));
 OA21x2_ASAP7_75t_R _12498_ (.A1(_05547_),
    .A2(_10142_),
    .B(_05597_),
    .Y(_05598_));
 XNOR2x1_ASAP7_75t_R _12499_ (.B(_05598_),
    .Y(_10023_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _12500_ (.A(_10023_),
    .Y(_10025_));
 AND3x1_ASAP7_75t_R _12501_ (.A(_00510_),
    .B(_03828_),
    .C(_03661_),
    .Y(_05599_));
 OA21x2_ASAP7_75t_R _12502_ (.A1(_03606_),
    .A2(_03670_),
    .B(_00514_),
    .Y(_05600_));
 AND3x1_ASAP7_75t_R _12503_ (.A(_00511_),
    .B(_03828_),
    .C(_03661_),
    .Y(_05601_));
 OA21x2_ASAP7_75t_R _12504_ (.A1(_03667_),
    .A2(_03670_),
    .B(_00515_),
    .Y(_05602_));
 OA33x2_ASAP7_75t_R _12505_ (.A1(_03866_),
    .A2(_05599_),
    .A3(_05600_),
    .B1(_05601_),
    .B2(_05602_),
    .B3(_03869_),
    .Y(_05603_));
 INVx1_ASAP7_75t_R _12506_ (.A(_00508_),
    .Y(_05604_));
 AND2x2_ASAP7_75t_R _12507_ (.A(_04610_),
    .B(_00513_),
    .Y(_05605_));
 AO21x1_ASAP7_75t_R _12508_ (.A1(_04609_),
    .A2(_00509_),
    .B(_05605_),
    .Y(_05606_));
 AOI22x1_ASAP7_75t_R _12509_ (.A1(_00512_),
    .A2(_04576_),
    .B1(_05606_),
    .B2(_03665_),
    .Y(_05607_));
 OA211x2_ASAP7_75t_R _12510_ (.A1(_03839_),
    .A2(_05607_),
    .B(_03802_),
    .C(_03737_),
    .Y(_05608_));
 OAI22x1_ASAP7_75t_R _12511_ (.A1(_05604_),
    .A2(_04575_),
    .B1(_05608_),
    .B2(_04164_),
    .Y(_05609_));
 AND3x1_ASAP7_75t_R _12512_ (.A(_03868_),
    .B(_05603_),
    .C(_05609_),
    .Y(_05610_));
 AND2x2_ASAP7_75t_R _12513_ (.A(_00502_),
    .B(_03890_),
    .Y(_05611_));
 AO221x1_ASAP7_75t_R _12514_ (.A1(_00503_),
    .A2(_04921_),
    .B1(_04804_),
    .B2(_03861_),
    .C(_05611_),
    .Y(_05612_));
 OA211x2_ASAP7_75t_R _12515_ (.A1(_00501_),
    .A2(_04952_),
    .B(_04627_),
    .C(_05612_),
    .Y(_05613_));
 AND3x1_ASAP7_75t_R _12516_ (.A(_04455_),
    .B(_04584_),
    .C(_00507_),
    .Y(_05614_));
 AO21x1_ASAP7_75t_R _12517_ (.A1(_00506_),
    .A2(_03782_),
    .B(_05614_),
    .Y(_05615_));
 AND3x1_ASAP7_75t_R _12518_ (.A(_04455_),
    .B(_04597_),
    .C(_00505_),
    .Y(_05616_));
 AO21x1_ASAP7_75t_R _12519_ (.A1(_00504_),
    .A2(_03782_),
    .B(_05616_),
    .Y(_05617_));
 AO221x2_ASAP7_75t_R _12520_ (.A1(_04440_),
    .A2(_05615_),
    .B1(_05617_),
    .B2(_04727_),
    .C(_04959_),
    .Y(_05618_));
 AND3x1_ASAP7_75t_R _12521_ (.A(_03843_),
    .B(_03762_),
    .C(_00527_),
    .Y(_05619_));
 AO21x1_ASAP7_75t_R _12522_ (.A1(_00526_),
    .A2(_03761_),
    .B(_05619_),
    .Y(_05620_));
 AND2x2_ASAP7_75t_R _12523_ (.A(_00530_),
    .B(_03671_),
    .Y(_05621_));
 AO221x1_ASAP7_75t_R _12524_ (.A1(_00531_),
    .A2(_03728_),
    .B1(_03735_),
    .B2(_03828_),
    .C(_05621_),
    .Y(_05622_));
 OA21x2_ASAP7_75t_R _12525_ (.A1(_04602_),
    .A2(_05620_),
    .B(_05622_),
    .Y(_05623_));
 INVx1_ASAP7_75t_R _12526_ (.A(_00524_),
    .Y(_05624_));
 AND2x2_ASAP7_75t_R _12527_ (.A(_03609_),
    .B(_00529_),
    .Y(_05625_));
 AO21x1_ASAP7_75t_R _12528_ (.A1(_04457_),
    .A2(_00525_),
    .B(_05625_),
    .Y(_05626_));
 AOI22x1_ASAP7_75t_R _12529_ (.A1(_00528_),
    .A2(_04576_),
    .B1(_05626_),
    .B2(_03717_),
    .Y(_05627_));
 OA211x2_ASAP7_75t_R _12530_ (.A1(_03839_),
    .A2(_05627_),
    .B(_03775_),
    .C(_03737_),
    .Y(_05628_));
 OAI22x1_ASAP7_75t_R _12531_ (.A1(_05624_),
    .A2(_04575_),
    .B1(_05628_),
    .B2(_04164_),
    .Y(_05629_));
 OA211x2_ASAP7_75t_R _12532_ (.A1(_05218_),
    .A2(_05623_),
    .B(_05629_),
    .C(_03868_),
    .Y(_05630_));
 AO21x2_ASAP7_75t_R _12533_ (.A1(_00517_),
    .A2(_05409_),
    .B(_04499_),
    .Y(_05631_));
 AND3x1_ASAP7_75t_R _12534_ (.A(_03375_),
    .B(_04435_),
    .C(_00523_),
    .Y(_05632_));
 AO21x1_ASAP7_75t_R _12535_ (.A1(_00522_),
    .A2(_04242_),
    .B(_05632_),
    .Y(_05633_));
 OA222x2_ASAP7_75t_R _12536_ (.A1(_00521_),
    .A2(_04952_),
    .B1(_05633_),
    .B2(_04454_),
    .C1(_04492_),
    .C2(_00520_),
    .Y(_05634_));
 AND3x1_ASAP7_75t_R _12537_ (.A(_03843_),
    .B(_04460_),
    .C(_00519_),
    .Y(_05635_));
 AO21x1_ASAP7_75t_R _12538_ (.A1(_00518_),
    .A2(_04236_),
    .B(_05635_),
    .Y(_05636_));
 AO32x1_ASAP7_75t_R _12539_ (.A1(_03518_),
    .A2(_04587_),
    .A3(_05636_),
    .B1(_03702_),
    .B2(_00516_),
    .Y(_05637_));
 AO32x2_ASAP7_75t_R _12540_ (.A1(_03655_),
    .A2(_04920_),
    .A3(_05634_),
    .B1(_05637_),
    .B2(_03701_),
    .Y(_05638_));
 OA33x2_ASAP7_75t_R _12541_ (.A1(_05610_),
    .A2(_05613_),
    .A3(_05618_),
    .B1(_05630_),
    .B2(_05631_),
    .B3(_05638_),
    .Y(_05639_));
 BUFx6f_ASAP7_75t_R _12542_ (.A(_05639_),
    .Y(_10024_));
 BUFx12f_ASAP7_75t_R _12543_ (.A(_04921_),
    .Y(_05640_));
 AO32x1_ASAP7_75t_R _12544_ (.A1(_04171_),
    .A2(_04172_),
    .A3(_03852_),
    .B1(_05640_),
    .B2(_04848_),
    .Y(_05641_));
 OA21x2_ASAP7_75t_R _12545_ (.A1(_05347_),
    .A2(_05641_),
    .B(_05346_),
    .Y(_05642_));
 AO21x2_ASAP7_75t_R _12546_ (.A1(_04174_),
    .A2(_05549_),
    .B(_05642_),
    .Y(_10140_));
 AO221x1_ASAP7_75t_R _12547_ (.A1(_03974_),
    .A2(_00556_),
    .B1(_04021_),
    .B2(_00554_),
    .C(_04028_),
    .Y(_05643_));
 AND2x2_ASAP7_75t_R _12548_ (.A(_03925_),
    .B(_00555_),
    .Y(_05644_));
 AO211x2_ASAP7_75t_R _12549_ (.A1(_04113_),
    .A2(_00553_),
    .B(_05644_),
    .C(_04992_),
    .Y(_05645_));
 AO221x1_ASAP7_75t_R _12550_ (.A1(_04071_),
    .A2(_00553_),
    .B1(_05643_),
    .B2(_05645_),
    .C(_03920_),
    .Y(_05646_));
 AND2x2_ASAP7_75t_R _12551_ (.A(_04105_),
    .B(_00563_),
    .Y(_05647_));
 AO21x1_ASAP7_75t_R _12552_ (.A1(_04073_),
    .A2(_00561_),
    .B(_05647_),
    .Y(_05648_));
 AO21x1_ASAP7_75t_R _12553_ (.A1(_00564_),
    .A2(_03961_),
    .B(_03413_),
    .Y(_05649_));
 AO221x1_ASAP7_75t_R _12554_ (.A1(_00562_),
    .A2(_04983_),
    .B1(_05648_),
    .B2(_04088_),
    .C(_05649_),
    .Y(_05650_));
 AOI21x1_ASAP7_75t_R _12555_ (.A1(_05646_),
    .A2(_05650_),
    .B(_04008_),
    .Y(_05651_));
 INVx2_ASAP7_75t_R _12556_ (.A(_00557_),
    .Y(_05652_));
 NAND2x1_ASAP7_75t_R _12557_ (.A(_04017_),
    .B(_00559_),
    .Y(_05653_));
 OA211x2_ASAP7_75t_R _12558_ (.A1(_04269_),
    .A2(_05652_),
    .B(_05653_),
    .C(_03998_),
    .Y(_05654_));
 INVx3_ASAP7_75t_R _12559_ (.A(_00560_),
    .Y(_05655_));
 OA21x2_ASAP7_75t_R _12560_ (.A1(_04520_),
    .A2(_05655_),
    .B(_04532_),
    .Y(_05656_));
 INVx1_ASAP7_75t_R _12561_ (.A(_00558_),
    .Y(_05657_));
 OR4x1_ASAP7_75t_R _12562_ (.A(_03929_),
    .B(_04105_),
    .C(_03983_),
    .D(_05657_),
    .Y(_05658_));
 OA211x2_ASAP7_75t_R _12563_ (.A1(_05654_),
    .A2(_05656_),
    .B(_04279_),
    .C(_05658_),
    .Y(_05659_));
 INVx2_ASAP7_75t_R _12564_ (.A(_00549_),
    .Y(_05660_));
 NAND2x1_ASAP7_75t_R _12565_ (.A(_04017_),
    .B(_00551_),
    .Y(_05661_));
 OA211x2_ASAP7_75t_R _12566_ (.A1(_04269_),
    .A2(_05660_),
    .B(_05661_),
    .C(_03998_),
    .Y(_05662_));
 INVx1_ASAP7_75t_R _12567_ (.A(_00552_),
    .Y(_05663_));
 OA21x2_ASAP7_75t_R _12568_ (.A1(_03991_),
    .A2(_05663_),
    .B(_04532_),
    .Y(_05664_));
 INVx1_ASAP7_75t_R _12569_ (.A(_00550_),
    .Y(_05665_));
 OR4x1_ASAP7_75t_R _12570_ (.A(_03929_),
    .B(_04105_),
    .C(_03983_),
    .D(_05665_),
    .Y(_05666_));
 OA211x2_ASAP7_75t_R _12571_ (.A1(_05662_),
    .A2(_05664_),
    .B(_04097_),
    .C(_05666_),
    .Y(_05667_));
 OA21x2_ASAP7_75t_R _12572_ (.A1(_05659_),
    .A2(_05667_),
    .B(_04296_),
    .Y(_05668_));
 OAI21x1_ASAP7_75t_R _12573_ (.A1(_05651_),
    .A2(_05668_),
    .B(_04763_),
    .Y(_05669_));
 AND2x2_ASAP7_75t_R _12574_ (.A(_03978_),
    .B(_00548_),
    .Y(_05670_));
 AO21x1_ASAP7_75t_R _12575_ (.A1(_04028_),
    .A2(_00547_),
    .B(_05670_),
    .Y(_05671_));
 AND3x1_ASAP7_75t_R _12576_ (.A(_03978_),
    .B(_04314_),
    .C(_00546_),
    .Y(_05672_));
 AO21x1_ASAP7_75t_R _12577_ (.A1(_00545_),
    .A2(_05590_),
    .B(_05672_),
    .Y(_05673_));
 AO221x1_ASAP7_75t_R _12578_ (.A1(_04270_),
    .A2(_05671_),
    .B1(_05673_),
    .B2(_04995_),
    .C(_04541_),
    .Y(_05674_));
 AND2x2_ASAP7_75t_R _12579_ (.A(_04025_),
    .B(_00543_),
    .Y(_05675_));
 AO21x1_ASAP7_75t_R _12580_ (.A1(_03954_),
    .A2(_00541_),
    .B(_05675_),
    .Y(_05676_));
 AO22x1_ASAP7_75t_R _12581_ (.A1(_00544_),
    .A2(_03961_),
    .B1(_05676_),
    .B2(_03950_),
    .Y(_05677_));
 AO21x1_ASAP7_75t_R _12582_ (.A1(_00542_),
    .A2(_04266_),
    .B(_03966_),
    .Y(_05678_));
 OA21x2_ASAP7_75t_R _12583_ (.A1(_05677_),
    .A2(_05678_),
    .B(_04156_),
    .Y(_05679_));
 AO22x1_ASAP7_75t_R _12584_ (.A1(_04028_),
    .A2(_00533_),
    .B1(_00534_),
    .B2(_04101_),
    .Y(_05680_));
 AND2x2_ASAP7_75t_R _12585_ (.A(_03932_),
    .B(_00536_),
    .Y(_05681_));
 AO21x1_ASAP7_75t_R _12586_ (.A1(_04037_),
    .A2(_00535_),
    .B(_05681_),
    .Y(_05682_));
 AO21x1_ASAP7_75t_R _12587_ (.A1(_04018_),
    .A2(_05682_),
    .B(_03965_),
    .Y(_05683_));
 AND2x2_ASAP7_75t_R _12588_ (.A(_04023_),
    .B(_00533_),
    .Y(_05684_));
 AO221x1_ASAP7_75t_R _12589_ (.A1(_03992_),
    .A2(_05680_),
    .B1(_05683_),
    .B2(_04142_),
    .C(_05684_),
    .Y(_05685_));
 AND2x2_ASAP7_75t_R _12590_ (.A(_03941_),
    .B(_00540_),
    .Y(_05686_));
 AO21x1_ASAP7_75t_R _12591_ (.A1(_03998_),
    .A2(_00539_),
    .B(_05686_),
    .Y(_05687_));
 AO21x1_ASAP7_75t_R _12592_ (.A1(_04106_),
    .A2(_05687_),
    .B(_03946_),
    .Y(_05688_));
 AND3x1_ASAP7_75t_R _12593_ (.A(_04033_),
    .B(_04314_),
    .C(_00538_),
    .Y(_05689_));
 OA21x2_ASAP7_75t_R _12594_ (.A1(_04037_),
    .A2(_03983_),
    .B(_00537_),
    .Y(_05690_));
 OA21x2_ASAP7_75t_R _12595_ (.A1(_05689_),
    .A2(_05690_),
    .B(_03937_),
    .Y(_05691_));
 OA21x2_ASAP7_75t_R _12596_ (.A1(_05688_),
    .A2(_05691_),
    .B(_04414_),
    .Y(_05692_));
 AO221x1_ASAP7_75t_R _12597_ (.A1(_05674_),
    .A2(_05679_),
    .B1(_05685_),
    .B2(_05692_),
    .C(_04051_),
    .Y(_05693_));
 AO21x2_ASAP7_75t_R _12598_ (.A1(_05669_),
    .A2(_05693_),
    .B(_04055_),
    .Y(_05694_));
 NAND2x1_ASAP7_75t_R _12599_ (.A(_05547_),
    .B(_05694_),
    .Y(_05695_));
 OA21x2_ASAP7_75t_R _12600_ (.A1(_05547_),
    .A2(_10140_),
    .B(_05695_),
    .Y(_05696_));
 XNOR2x1_ASAP7_75t_R _12601_ (.B(_05696_),
    .Y(_10028_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _12602_ (.A(_10028_),
    .Y(_10030_));
 AOI21x1_ASAP7_75t_R _12603_ (.A1(_03648_),
    .A2(_04627_),
    .B(_04959_),
    .Y(_05697_));
 AO21x2_ASAP7_75t_R _12604_ (.A1(_03827_),
    .A2(_03650_),
    .B(_03651_),
    .Y(_05698_));
 INVx1_ASAP7_75t_R _12605_ (.A(_00539_),
    .Y(_05699_));
 INVx1_ASAP7_75t_R _12606_ (.A(_00540_),
    .Y(_05700_));
 OR3x1_ASAP7_75t_R _12607_ (.A(_03415_),
    .B(_03618_),
    .C(_05700_),
    .Y(_05701_));
 OA21x2_ASAP7_75t_R _12608_ (.A1(_05699_),
    .A2(_03885_),
    .B(_05701_),
    .Y(_05702_));
 OR4x1_ASAP7_75t_R _12609_ (.A(_03539_),
    .B(_03824_),
    .C(_05698_),
    .D(_05702_),
    .Y(_05703_));
 AND2x2_ASAP7_75t_R _12610_ (.A(_00538_),
    .B(_03813_),
    .Y(_05704_));
 AND2x2_ASAP7_75t_R _12611_ (.A(_00537_),
    .B(_03585_),
    .Y(_05705_));
 OAI21x1_ASAP7_75t_R _12612_ (.A1(_05704_),
    .A2(_05705_),
    .B(_03721_),
    .Y(_05706_));
 INVx1_ASAP7_75t_R _12613_ (.A(_00533_),
    .Y(_01229_));
 AO21x1_ASAP7_75t_R _12614_ (.A1(_03506_),
    .A2(_03508_),
    .B(_03648_),
    .Y(_05707_));
 INVx1_ASAP7_75t_R _12615_ (.A(_00535_),
    .Y(_05708_));
 INVx1_ASAP7_75t_R _12616_ (.A(_00534_),
    .Y(_05709_));
 NAND2x1_ASAP7_75t_R _12617_ (.A(_03619_),
    .B(_00536_),
    .Y(_05710_));
 OA211x2_ASAP7_75t_R _12618_ (.A1(_03636_),
    .A2(_05709_),
    .B(_05710_),
    .C(_03614_),
    .Y(_05711_));
 AO21x1_ASAP7_75t_R _12619_ (.A1(_05708_),
    .A2(_04442_),
    .B(_05711_),
    .Y(_05712_));
 NAND2x2_ASAP7_75t_R _12620_ (.A(_03660_),
    .B(_03771_),
    .Y(_05713_));
 AO221x1_ASAP7_75t_R _12621_ (.A1(_01229_),
    .A2(_05707_),
    .B1(_05712_),
    .B2(_04916_),
    .C(_05713_),
    .Y(_05714_));
 AND4x2_ASAP7_75t_R _12622_ (.A(_05697_),
    .B(_05703_),
    .C(_05706_),
    .D(_05714_),
    .Y(_05715_));
 AND2x2_ASAP7_75t_R _12623_ (.A(_03685_),
    .B(_00546_),
    .Y(_05716_));
 AO21x1_ASAP7_75t_R _12624_ (.A1(_03744_),
    .A2(_00542_),
    .B(_05716_),
    .Y(_05717_));
 AO22x1_ASAP7_75t_R _12625_ (.A1(_00545_),
    .A2(_04456_),
    .B1(_05717_),
    .B2(_03664_),
    .Y(_05718_));
 NAND2x1_ASAP7_75t_R _12626_ (.A(_03715_),
    .B(_05718_),
    .Y(_05719_));
 AO21x1_ASAP7_75t_R _12627_ (.A1(_03824_),
    .A2(_05719_),
    .B(_04214_),
    .Y(_05720_));
 NAND2x1_ASAP7_75t_R _12628_ (.A(_00541_),
    .B(_03750_),
    .Y(_05721_));
 AND3x1_ASAP7_75t_R _12629_ (.A(_00543_),
    .B(_03860_),
    .C(_03830_),
    .Y(_05722_));
 AOI221x1_ASAP7_75t_R _12630_ (.A1(_00548_),
    .A2(_04198_),
    .B1(_04199_),
    .B2(_00547_),
    .C(_05722_),
    .Y(_05723_));
 AOI21x1_ASAP7_75t_R _12631_ (.A1(_00544_),
    .A2(_03834_),
    .B(_04454_),
    .Y(_05724_));
 AO221x2_ASAP7_75t_R _12632_ (.A1(_05720_),
    .A2(_05721_),
    .B1(_05723_),
    .B2(_05724_),
    .C(_03740_),
    .Y(_05725_));
 OR3x1_ASAP7_75t_R _12633_ (.A(_03419_),
    .B(_03629_),
    .C(_05655_),
    .Y(_05726_));
 INVx1_ASAP7_75t_R _12634_ (.A(_00563_),
    .Y(_05727_));
 AO21x1_ASAP7_75t_R _12635_ (.A1(_03443_),
    .A2(_03716_),
    .B(_05727_),
    .Y(_05728_));
 INVx1_ASAP7_75t_R _12636_ (.A(_00564_),
    .Y(_05729_));
 OR3x1_ASAP7_75t_R _12637_ (.A(_03415_),
    .B(_03618_),
    .C(_05729_),
    .Y(_05730_));
 AO22x1_ASAP7_75t_R _12638_ (.A1(_04350_),
    .A2(_03734_),
    .B1(_05728_),
    .B2(_05730_),
    .Y(_05731_));
 INVx2_ASAP7_75t_R _12639_ (.A(_00559_),
    .Y(_05732_));
 AO21x1_ASAP7_75t_R _12640_ (.A1(_03443_),
    .A2(_03690_),
    .B(_05732_),
    .Y(_05733_));
 AO21x1_ASAP7_75t_R _12641_ (.A1(_03681_),
    .A2(_05733_),
    .B(_03679_),
    .Y(_05734_));
 OA211x2_ASAP7_75t_R _12642_ (.A1(_03871_),
    .A2(_05726_),
    .B(_05731_),
    .C(_05734_),
    .Y(_05735_));
 AND2x2_ASAP7_75t_R _12643_ (.A(_03685_),
    .B(_00562_),
    .Y(_05736_));
 AO21x1_ASAP7_75t_R _12644_ (.A1(_03744_),
    .A2(_00558_),
    .B(_05736_),
    .Y(_05737_));
 AOI22x1_ASAP7_75t_R _12645_ (.A1(_00561_),
    .A2(_04456_),
    .B1(_05737_),
    .B2(_03664_),
    .Y(_05738_));
 OA211x2_ASAP7_75t_R _12646_ (.A1(_03480_),
    .A2(_05738_),
    .B(_04212_),
    .C(_03736_),
    .Y(_05739_));
 OA22x2_ASAP7_75t_R _12647_ (.A1(_05652_),
    .A2(_04218_),
    .B1(_05739_),
    .B2(_04214_),
    .Y(_05740_));
 OR3x1_ASAP7_75t_R _12648_ (.A(_04468_),
    .B(_05735_),
    .C(_05740_),
    .Y(_05741_));
 INVx1_ASAP7_75t_R _12649_ (.A(_00555_),
    .Y(_05742_));
 OA211x2_ASAP7_75t_R _12650_ (.A1(_03606_),
    .A2(_03681_),
    .B(_03710_),
    .C(_05742_),
    .Y(_05743_));
 INVx1_ASAP7_75t_R _12651_ (.A(_00556_),
    .Y(_05744_));
 NAND2x1_ASAP7_75t_R _12652_ (.A(_03632_),
    .B(_00554_),
    .Y(_05745_));
 OA211x2_ASAP7_75t_R _12653_ (.A1(_03632_),
    .A2(_05744_),
    .B(_03881_),
    .C(_05745_),
    .Y(_05746_));
 NOR2x1_ASAP7_75t_R _12654_ (.A(_05743_),
    .B(_05746_),
    .Y(_05747_));
 OA211x2_ASAP7_75t_R _12655_ (.A1(_00553_),
    .A2(_04492_),
    .B(_03653_),
    .C(_04244_),
    .Y(_05748_));
 AND2x2_ASAP7_75t_R _12656_ (.A(_03897_),
    .B(_00552_),
    .Y(_05749_));
 AO21x1_ASAP7_75t_R _12657_ (.A1(_03632_),
    .A2(_00550_),
    .B(_05749_),
    .Y(_05750_));
 OA222x2_ASAP7_75t_R _12658_ (.A1(_04163_),
    .A2(_03772_),
    .B1(_05750_),
    .B2(_03805_),
    .C1(_03865_),
    .C2(_00551_),
    .Y(_05751_));
 NAND2x1_ASAP7_75t_R _12659_ (.A(_05660_),
    .B(_03702_),
    .Y(_05752_));
 AOI221x1_ASAP7_75t_R _12660_ (.A1(_05747_),
    .A2(_05748_),
    .B1(_05751_),
    .B2(_05752_),
    .C(_03723_),
    .Y(_05753_));
 AO22x2_ASAP7_75t_R _12661_ (.A1(_05715_),
    .A2(_05725_),
    .B1(_05741_),
    .B2(_05753_),
    .Y(_05754_));
 BUFx4f_ASAP7_75t_R _12662_ (.A(_05754_),
    .Y(_10027_));
 INVx4_ASAP7_75t_R _12663_ (.A(_10027_),
    .Y(_10029_));
 AND2x2_ASAP7_75t_R _12664_ (.A(_03378_),
    .B(_03483_),
    .Y(_05755_));
 AO32x1_ASAP7_75t_R _12665_ (.A1(_04171_),
    .A2(_04172_),
    .A3(_05640_),
    .B1(_05755_),
    .B2(_04848_),
    .Y(_05756_));
 OA21x2_ASAP7_75t_R _12666_ (.A1(_05347_),
    .A2(_05756_),
    .B(_04168_),
    .Y(_05757_));
 OA211x2_ASAP7_75t_R _12667_ (.A1(_05347_),
    .A2(_05641_),
    .B(_04174_),
    .C(_04168_),
    .Y(_05758_));
 AO21x2_ASAP7_75t_R _12668_ (.A1(_05346_),
    .A2(_05757_),
    .B(_05758_),
    .Y(_10138_));
 AND2x2_ASAP7_75t_R _12669_ (.A(_03933_),
    .B(_00569_),
    .Y(_05759_));
 AO21x1_ASAP7_75t_R _12670_ (.A1(_03930_),
    .A2(_00568_),
    .B(_05759_),
    .Y(_05760_));
 AO21x1_ASAP7_75t_R _12671_ (.A1(_03927_),
    .A2(_05760_),
    .B(_04032_),
    .Y(_05761_));
 AO22x1_ASAP7_75t_R _12672_ (.A1(_03950_),
    .A2(_00566_),
    .B1(_00567_),
    .B2(_04101_),
    .Y(_05762_));
 AO22x1_ASAP7_75t_R _12673_ (.A1(_04071_),
    .A2(_00566_),
    .B1(_05762_),
    .B2(_04114_),
    .Y(_05763_));
 AO21x1_ASAP7_75t_R _12674_ (.A1(_03381_),
    .A2(_05761_),
    .B(_05763_),
    .Y(_05764_));
 AND2x2_ASAP7_75t_R _12675_ (.A(_04015_),
    .B(_00573_),
    .Y(_05765_));
 AO21x1_ASAP7_75t_R _12676_ (.A1(_04556_),
    .A2(_00572_),
    .B(_05765_),
    .Y(_05766_));
 AND3x1_ASAP7_75t_R _12677_ (.A(_04532_),
    .B(_04559_),
    .C(_00571_),
    .Y(_05767_));
 AO21x1_ASAP7_75t_R _12678_ (.A1(_00570_),
    .A2(_04535_),
    .B(_05767_),
    .Y(_05768_));
 AO221x1_ASAP7_75t_R _12679_ (.A1(_04530_),
    .A2(_05766_),
    .B1(_05768_),
    .B2(_04540_),
    .C(_04542_),
    .Y(_05769_));
 AND2x2_ASAP7_75t_R _12680_ (.A(_04015_),
    .B(_00581_),
    .Y(_05770_));
 AO21x1_ASAP7_75t_R _12681_ (.A1(_04556_),
    .A2(_00580_),
    .B(_05770_),
    .Y(_05771_));
 AND3x1_ASAP7_75t_R _12682_ (.A(_04532_),
    .B(_04559_),
    .C(_00579_),
    .Y(_05772_));
 AO21x1_ASAP7_75t_R _12683_ (.A1(_00578_),
    .A2(_04535_),
    .B(_05772_),
    .Y(_05773_));
 AO221x1_ASAP7_75t_R _12684_ (.A1(_04502_),
    .A2(_05771_),
    .B1(_05773_),
    .B2(_04540_),
    .C(_04094_),
    .Y(_05774_));
 AND2x2_ASAP7_75t_R _12685_ (.A(_04105_),
    .B(_00576_),
    .Y(_05775_));
 AO21x1_ASAP7_75t_R _12686_ (.A1(_04103_),
    .A2(_00574_),
    .B(_05775_),
    .Y(_05776_));
 AO22x1_ASAP7_75t_R _12687_ (.A1(_00577_),
    .A2(_04090_),
    .B1(_05776_),
    .B2(_04079_),
    .Y(_05777_));
 AO21x1_ASAP7_75t_R _12688_ (.A1(_00575_),
    .A2(_04983_),
    .B(_04130_),
    .Y(_05778_));
 OA21x2_ASAP7_75t_R _12689_ (.A1(_05777_),
    .A2(_05778_),
    .B(_04280_),
    .Y(_05779_));
 AO32x1_ASAP7_75t_R _12690_ (.A1(_04099_),
    .A2(_05764_),
    .A3(_05769_),
    .B1(_05774_),
    .B2(_05779_),
    .Y(_05780_));
 AND2x2_ASAP7_75t_R _12691_ (.A(_04992_),
    .B(_00589_),
    .Y(_05781_));
 AO21x1_ASAP7_75t_R _12692_ (.A1(_04079_),
    .A2(_00588_),
    .B(_05781_),
    .Y(_05782_));
 AND3x1_ASAP7_75t_R _12693_ (.A(_04992_),
    .B(_04315_),
    .C(_00587_),
    .Y(_05783_));
 AO21x1_ASAP7_75t_R _12694_ (.A1(_00586_),
    .A2(_04991_),
    .B(_05783_),
    .Y(_05784_));
 AO221x1_ASAP7_75t_R _12695_ (.A1(_04988_),
    .A2(_05782_),
    .B1(_05784_),
    .B2(_04996_),
    .C(_04298_),
    .Y(_05785_));
 AND2x2_ASAP7_75t_R _12696_ (.A(_04992_),
    .B(_00597_),
    .Y(_05786_));
 AO21x1_ASAP7_75t_R _12697_ (.A1(_04079_),
    .A2(_00596_),
    .B(_05786_),
    .Y(_05787_));
 AND3x1_ASAP7_75t_R _12698_ (.A(_04992_),
    .B(_04315_),
    .C(_00595_),
    .Y(_05788_));
 AO21x1_ASAP7_75t_R _12699_ (.A1(_00594_),
    .A2(_04991_),
    .B(_05788_),
    .Y(_05789_));
 AO221x1_ASAP7_75t_R _12700_ (.A1(_04988_),
    .A2(_05787_),
    .B1(_05789_),
    .B2(_04996_),
    .C(_04304_),
    .Y(_05790_));
 AND3x1_ASAP7_75t_R _12701_ (.A(_04763_),
    .B(_05785_),
    .C(_05790_),
    .Y(_05791_));
 AO221x1_ASAP7_75t_R _12702_ (.A1(_04643_),
    .A2(_00593_),
    .B1(_04069_),
    .B2(_00591_),
    .C(_04414_),
    .Y(_05792_));
 AO221x1_ASAP7_75t_R _12703_ (.A1(_04643_),
    .A2(_00585_),
    .B1(_04632_),
    .B2(_00583_),
    .C(_04156_),
    .Y(_05793_));
 AO21x1_ASAP7_75t_R _12704_ (.A1(_05792_),
    .A2(_05793_),
    .B(_04089_),
    .Y(_05794_));
 INVx1_ASAP7_75t_R _12705_ (.A(_00584_),
    .Y(_05795_));
 NAND2x1_ASAP7_75t_R _12706_ (.A(_04084_),
    .B(_00582_),
    .Y(_05796_));
 OA211x2_ASAP7_75t_R _12707_ (.A1(_04074_),
    .A2(_05795_),
    .B(_03997_),
    .C(_05796_),
    .Y(_05797_));
 INVx1_ASAP7_75t_R _12708_ (.A(_00590_),
    .Y(_05798_));
 NAND2x1_ASAP7_75t_R _12709_ (.A(_03975_),
    .B(_00592_),
    .Y(_05799_));
 OA211x2_ASAP7_75t_R _12710_ (.A1(_04530_),
    .A2(_05798_),
    .B(_04156_),
    .C(_05799_),
    .Y(_05800_));
 OAI21x1_ASAP7_75t_R _12711_ (.A1(_05797_),
    .A2(_05800_),
    .B(_04089_),
    .Y(_05801_));
 AO21x1_ASAP7_75t_R _12712_ (.A1(_05794_),
    .A2(_05801_),
    .B(_04120_),
    .Y(_05802_));
 AO221x2_ASAP7_75t_R _12713_ (.A1(_04122_),
    .A2(_05780_),
    .B1(_05791_),
    .B2(_05802_),
    .C(_04565_),
    .Y(_05803_));
 NAND2x1_ASAP7_75t_R _12714_ (.A(_05547_),
    .B(_05803_),
    .Y(_05804_));
 OA21x2_ASAP7_75t_R _12715_ (.A1(_05547_),
    .A2(_10138_),
    .B(_05804_),
    .Y(_05805_));
 XNOR2x1_ASAP7_75t_R _12716_ (.B(_05805_),
    .Y(_10033_),
    .A(_03914_));
 INVx1_ASAP7_75t_R _12717_ (.A(_10033_),
    .Y(_10035_));
 OR4x1_ASAP7_75t_R _12718_ (.A(_00570_),
    .B(_03820_),
    .C(_04591_),
    .D(_03783_),
    .Y(_05806_));
 AO221x1_ASAP7_75t_R _12719_ (.A1(_03815_),
    .A2(_04624_),
    .B1(_03804_),
    .B2(_03803_),
    .C(_00572_),
    .Y(_05807_));
 AND4x1_ASAP7_75t_R _12720_ (.A(_03822_),
    .B(_04920_),
    .C(_05806_),
    .D(_05807_),
    .Y(_05808_));
 OR3x1_ASAP7_75t_R _12721_ (.A(_00571_),
    .B(_03820_),
    .C(_03783_),
    .Y(_05809_));
 AO21x1_ASAP7_75t_R _12722_ (.A1(_03862_),
    .A2(_03889_),
    .B(_00573_),
    .Y(_05810_));
 AO21x1_ASAP7_75t_R _12723_ (.A1(_05809_),
    .A2(_05810_),
    .B(_03587_),
    .Y(_05811_));
 OR3x1_ASAP7_75t_R _12724_ (.A(_00576_),
    .B(_05640_),
    .C(_04948_),
    .Y(_05812_));
 OR3x1_ASAP7_75t_R _12725_ (.A(_00580_),
    .B(_03837_),
    .C(_03887_),
    .Y(_05813_));
 OR3x1_ASAP7_75t_R _12726_ (.A(_00577_),
    .B(_03796_),
    .C(_04948_),
    .Y(_05814_));
 AND3x1_ASAP7_75t_R _12727_ (.A(_04916_),
    .B(_03853_),
    .C(_00581_),
    .Y(_05815_));
 AO21x1_ASAP7_75t_R _12728_ (.A1(_00580_),
    .A2(_03891_),
    .B(_05815_),
    .Y(_05816_));
 OA21x2_ASAP7_75t_R _12729_ (.A1(_03707_),
    .A2(_05816_),
    .B(_03868_),
    .Y(_05817_));
 AND4x2_ASAP7_75t_R _12730_ (.A(_05812_),
    .B(_05813_),
    .C(_05814_),
    .D(_05817_),
    .Y(_05818_));
 INVx1_ASAP7_75t_R _12731_ (.A(_00574_),
    .Y(_05819_));
 AND2x2_ASAP7_75t_R _12732_ (.A(_05332_),
    .B(_00579_),
    .Y(_05820_));
 AO21x1_ASAP7_75t_R _12733_ (.A1(_05331_),
    .A2(_00575_),
    .B(_05820_),
    .Y(_05821_));
 AOI22x1_ASAP7_75t_R _12734_ (.A1(_00578_),
    .A2(_04936_),
    .B1(_05821_),
    .B2(_04624_),
    .Y(_05822_));
 OA211x2_ASAP7_75t_R _12735_ (.A1(_03482_),
    .A2(_05822_),
    .B(_03889_),
    .C(_03862_),
    .Y(_05823_));
 OAI22x1_ASAP7_75t_R _12736_ (.A1(_05819_),
    .A2(_04934_),
    .B1(_05823_),
    .B2(_04165_),
    .Y(_05824_));
 AO221x2_ASAP7_75t_R _12737_ (.A1(_05808_),
    .A2(_05811_),
    .B1(_05818_),
    .B2(_05824_),
    .C(_04452_),
    .Y(_05825_));
 AND2x2_ASAP7_75t_R _12738_ (.A(_00587_),
    .B(_04591_),
    .Y(_05826_));
 AO21x1_ASAP7_75t_R _12739_ (.A1(_00586_),
    .A2(_03879_),
    .B(_05826_),
    .Y(_05827_));
 AND2x2_ASAP7_75t_R _12740_ (.A(_00588_),
    .B(_03711_),
    .Y(_05828_));
 AO221x1_ASAP7_75t_R _12741_ (.A1(_00589_),
    .A2(_03887_),
    .B1(_03889_),
    .B2(_03862_),
    .C(_05828_),
    .Y(_05829_));
 OA211x2_ASAP7_75t_R _12742_ (.A1(_03852_),
    .A2(_05827_),
    .B(_05829_),
    .C(_05403_),
    .Y(_05830_));
 AND3x1_ASAP7_75t_R _12743_ (.A(_03376_),
    .B(_04436_),
    .C(_00585_),
    .Y(_05831_));
 AO21x1_ASAP7_75t_R _12744_ (.A1(_00584_),
    .A2(_04595_),
    .B(_05831_),
    .Y(_05832_));
 AO32x1_ASAP7_75t_R _12745_ (.A1(_03655_),
    .A2(_04587_),
    .A3(_05832_),
    .B1(_03703_),
    .B2(_00582_),
    .Y(_05833_));
 AND2x2_ASAP7_75t_R _12746_ (.A(_04915_),
    .B(_05833_),
    .Y(_05834_));
 AO21x1_ASAP7_75t_R _12747_ (.A1(_00583_),
    .A2(_05409_),
    .B(_03809_),
    .Y(_05835_));
 AND3x1_ASAP7_75t_R _12748_ (.A(_00592_),
    .B(_03873_),
    .C(_03830_),
    .Y(_05836_));
 AO221x1_ASAP7_75t_R _12749_ (.A1(_00597_),
    .A2(_04198_),
    .B1(_04476_),
    .B2(_00596_),
    .C(_05836_),
    .Y(_05837_));
 AO21x1_ASAP7_75t_R _12750_ (.A1(_00593_),
    .A2(_05233_),
    .B(_05218_),
    .Y(_05838_));
 AND2x2_ASAP7_75t_R _12751_ (.A(_04938_),
    .B(_00595_),
    .Y(_05839_));
 AO21x1_ASAP7_75t_R _12752_ (.A1(_04937_),
    .A2(_00591_),
    .B(_05839_),
    .Y(_05840_));
 AOI22x1_ASAP7_75t_R _12753_ (.A1(_00594_),
    .A2(_05221_),
    .B1(_05840_),
    .B2(_05224_),
    .Y(_05841_));
 OA211x2_ASAP7_75t_R _12754_ (.A1(_05417_),
    .A2(_05841_),
    .B(_04592_),
    .C(_03873_),
    .Y(_05842_));
 OAI22x1_ASAP7_75t_R _12755_ (.A1(_05798_),
    .A2(_04934_),
    .B1(_05842_),
    .B2(_03786_),
    .Y(_05843_));
 OA211x2_ASAP7_75t_R _12756_ (.A1(_05837_),
    .A2(_05838_),
    .B(_03850_),
    .C(_05843_),
    .Y(_05844_));
 OR4x2_ASAP7_75t_R _12757_ (.A(_05830_),
    .B(_05834_),
    .C(_05835_),
    .D(_05844_),
    .Y(_05845_));
 AND3x4_ASAP7_75t_R _12758_ (.A(_03646_),
    .B(_03607_),
    .C(_04192_),
    .Y(_05846_));
 AND3x1_ASAP7_75t_R _12759_ (.A(_04053_),
    .B(_04624_),
    .C(_00569_),
    .Y(_05847_));
 AO21x1_ASAP7_75t_R _12760_ (.A1(_00568_),
    .A2(_04623_),
    .B(_05847_),
    .Y(_05848_));
 AO32x1_ASAP7_75t_R _12761_ (.A1(_00567_),
    .A2(_03814_),
    .A3(_05846_),
    .B1(_03901_),
    .B2(_05848_),
    .Y(_05849_));
 AO21x2_ASAP7_75t_R _12762_ (.A1(_00566_),
    .A2(_04622_),
    .B(_05849_),
    .Y(_05850_));
 AO21x2_ASAP7_75t_R _12763_ (.A1(_05825_),
    .A2(_05845_),
    .B(_05850_),
    .Y(_05851_));
 BUFx10_ASAP7_75t_R _12764_ (.A(_05851_),
    .Y(_10034_));
 NAND2x2_ASAP7_75t_R _12765_ (.A(_03843_),
    .B(_03528_),
    .Y(_05852_));
 INVx3_ASAP7_75t_R _12766_ (.A(_05852_),
    .Y(_05853_));
 AO32x1_ASAP7_75t_R _12767_ (.A1(_04171_),
    .A2(_04172_),
    .A3(_05755_),
    .B1(_05853_),
    .B2(_04848_),
    .Y(_05854_));
 OA21x2_ASAP7_75t_R _12768_ (.A1(_05347_),
    .A2(_05854_),
    .B(_05346_),
    .Y(_05855_));
 AO21x2_ASAP7_75t_R _12769_ (.A1(_04174_),
    .A2(_05757_),
    .B(_05855_),
    .Y(_10136_));
 AND2x2_ASAP7_75t_R _12770_ (.A(_03942_),
    .B(_00603_),
    .Y(_05856_));
 AO21x1_ASAP7_75t_R _12771_ (.A1(_04671_),
    .A2(_00602_),
    .B(_05856_),
    .Y(_05857_));
 AO21x1_ASAP7_75t_R _12772_ (.A1(_04502_),
    .A2(_05857_),
    .B(_04032_),
    .Y(_05858_));
 AO22x1_ASAP7_75t_R _12773_ (.A1(_04281_),
    .A2(_00600_),
    .B1(_00601_),
    .B2(_05073_),
    .Y(_05859_));
 AO22x1_ASAP7_75t_R _12774_ (.A1(_04504_),
    .A2(_00600_),
    .B1(_05859_),
    .B2(_04104_),
    .Y(_05860_));
 AO21x1_ASAP7_75t_R _12775_ (.A1(_04060_),
    .A2(_05858_),
    .B(_05860_),
    .Y(_05861_));
 AND2x2_ASAP7_75t_R _12776_ (.A(_04537_),
    .B(_00607_),
    .Y(_05862_));
 AO21x1_ASAP7_75t_R _12777_ (.A1(_04647_),
    .A2(_00606_),
    .B(_05862_),
    .Y(_05863_));
 AND3x1_ASAP7_75t_R _12778_ (.A(_04992_),
    .B(_03971_),
    .C(_00605_),
    .Y(_05864_));
 AO21x1_ASAP7_75t_R _12779_ (.A1(_00604_),
    .A2(_04991_),
    .B(_05864_),
    .Y(_05865_));
 AO221x1_ASAP7_75t_R _12780_ (.A1(_04988_),
    .A2(_05863_),
    .B1(_05865_),
    .B2(_04996_),
    .C(_04542_),
    .Y(_05866_));
 AND2x2_ASAP7_75t_R _12781_ (.A(_04532_),
    .B(_00615_),
    .Y(_05867_));
 AO21x1_ASAP7_75t_R _12782_ (.A1(_04531_),
    .A2(_00614_),
    .B(_05867_),
    .Y(_05868_));
 AND3x1_ASAP7_75t_R _12783_ (.A(_04537_),
    .B(_03971_),
    .C(_00613_),
    .Y(_05869_));
 AO21x1_ASAP7_75t_R _12784_ (.A1(_00612_),
    .A2(_04991_),
    .B(_05869_),
    .Y(_05870_));
 AO221x1_ASAP7_75t_R _12785_ (.A1(_04530_),
    .A2(_05868_),
    .B1(_05870_),
    .B2(_04540_),
    .C(_04542_),
    .Y(_05871_));
 AND2x2_ASAP7_75t_R _12786_ (.A(_04075_),
    .B(_00610_),
    .Y(_05872_));
 AO21x1_ASAP7_75t_R _12787_ (.A1(_04073_),
    .A2(_00608_),
    .B(_05872_),
    .Y(_05873_));
 AO22x1_ASAP7_75t_R _12788_ (.A1(_00611_),
    .A2(_04262_),
    .B1(_05873_),
    .B2(_04088_),
    .Y(_05874_));
 AO21x1_ASAP7_75t_R _12789_ (.A1(_00609_),
    .A2(_04983_),
    .B(_04130_),
    .Y(_05875_));
 OA21x2_ASAP7_75t_R _12790_ (.A1(_05874_),
    .A2(_05875_),
    .B(_03921_),
    .Y(_05876_));
 AO32x1_ASAP7_75t_R _12791_ (.A1(_04099_),
    .A2(_05861_),
    .A3(_05866_),
    .B1(_05871_),
    .B2(_05876_),
    .Y(_05877_));
 AND2x2_ASAP7_75t_R _12792_ (.A(_04307_),
    .B(_00623_),
    .Y(_05878_));
 AO21x1_ASAP7_75t_R _12793_ (.A1(_04088_),
    .A2(_00622_),
    .B(_05878_),
    .Y(_05879_));
 AND3x1_ASAP7_75t_R _12794_ (.A(_04307_),
    .B(_04315_),
    .C(_00621_),
    .Y(_05880_));
 AO21x1_ASAP7_75t_R _12795_ (.A1(_00620_),
    .A2(_04991_),
    .B(_05880_),
    .Y(_05881_));
 AO221x1_ASAP7_75t_R _12796_ (.A1(_04656_),
    .A2(_05879_),
    .B1(_05881_),
    .B2(_04996_),
    .C(_04298_),
    .Y(_05882_));
 AND2x2_ASAP7_75t_R _12797_ (.A(_04992_),
    .B(_00631_),
    .Y(_05883_));
 AO21x1_ASAP7_75t_R _12798_ (.A1(_04088_),
    .A2(_00630_),
    .B(_05883_),
    .Y(_05884_));
 AND3x1_ASAP7_75t_R _12799_ (.A(_04307_),
    .B(_04315_),
    .C(_00629_),
    .Y(_05885_));
 AO21x1_ASAP7_75t_R _12800_ (.A1(_00628_),
    .A2(_04991_),
    .B(_05885_),
    .Y(_05886_));
 AO221x1_ASAP7_75t_R _12801_ (.A1(_04988_),
    .A2(_05884_),
    .B1(_05886_),
    .B2(_04996_),
    .C(_04304_),
    .Y(_05887_));
 AND3x1_ASAP7_75t_R _12802_ (.A(_04763_),
    .B(_05882_),
    .C(_05887_),
    .Y(_05888_));
 AO221x1_ASAP7_75t_R _12803_ (.A1(_04255_),
    .A2(_00627_),
    .B1(_04069_),
    .B2(_00625_),
    .C(_03997_),
    .Y(_05889_));
 AO221x1_ASAP7_75t_R _12804_ (.A1(_04255_),
    .A2(_00619_),
    .B1(_04069_),
    .B2(_00617_),
    .C(_04156_),
    .Y(_05890_));
 AO21x1_ASAP7_75t_R _12805_ (.A1(_05889_),
    .A2(_05890_),
    .B(_04089_),
    .Y(_05891_));
 INVx1_ASAP7_75t_R _12806_ (.A(_00616_),
    .Y(_05892_));
 NAND2x1_ASAP7_75t_R _12807_ (.A(_03975_),
    .B(_00618_),
    .Y(_05893_));
 OA211x2_ASAP7_75t_R _12808_ (.A1(_04988_),
    .A2(_05892_),
    .B(_03997_),
    .C(_05893_),
    .Y(_05894_));
 INVx1_ASAP7_75t_R _12809_ (.A(_00624_),
    .Y(_05895_));
 NAND2x1_ASAP7_75t_R _12810_ (.A(_04643_),
    .B(_00626_),
    .Y(_05896_));
 OA211x2_ASAP7_75t_R _12811_ (.A1(_04988_),
    .A2(_05895_),
    .B(_04280_),
    .C(_05896_),
    .Y(_05897_));
 OAI21x1_ASAP7_75t_R _12812_ (.A1(_05894_),
    .A2(_05897_),
    .B(_04089_),
    .Y(_05898_));
 AO21x1_ASAP7_75t_R _12813_ (.A1(_05891_),
    .A2(_05898_),
    .B(_04120_),
    .Y(_05899_));
 AO221x2_ASAP7_75t_R _12814_ (.A1(_04122_),
    .A2(_05877_),
    .B1(_05888_),
    .B2(_05899_),
    .C(_04565_),
    .Y(_05900_));
 NAND2x1_ASAP7_75t_R _12815_ (.A(_05547_),
    .B(_05900_),
    .Y(_05901_));
 OA21x2_ASAP7_75t_R _12816_ (.A1(_05547_),
    .A2(_10136_),
    .B(_05901_),
    .Y(_05902_));
 XNOR2x1_ASAP7_75t_R _12817_ (.B(_05902_),
    .Y(_10038_),
    .A(_03913_));
 INVx1_ASAP7_75t_R _12818_ (.A(_10038_),
    .Y(_10040_));
 AND3x1_ASAP7_75t_R _12819_ (.A(_03376_),
    .B(_05224_),
    .C(_00623_),
    .Y(_05903_));
 AO21x1_ASAP7_75t_R _12820_ (.A1(_00622_),
    .A2(_04434_),
    .B(_05903_),
    .Y(_05904_));
 OA22x2_ASAP7_75t_R _12821_ (.A1(_00620_),
    .A2(_04492_),
    .B1(_05904_),
    .B2(_03826_),
    .Y(_05905_));
 OA211x2_ASAP7_75t_R _12822_ (.A1(_00621_),
    .A2(_04952_),
    .B(_04920_),
    .C(_03655_),
    .Y(_05906_));
 NAND2x1_ASAP7_75t_R _12823_ (.A(_05905_),
    .B(_05906_),
    .Y(_05907_));
 AND3x1_ASAP7_75t_R _12824_ (.A(_04596_),
    .B(_04436_),
    .C(_00627_),
    .Y(_05908_));
 AO21x1_ASAP7_75t_R _12825_ (.A1(_00626_),
    .A2(_04595_),
    .B(_05908_),
    .Y(_05909_));
 AND3x1_ASAP7_75t_R _12826_ (.A(_03663_),
    .B(_03853_),
    .C(_00631_),
    .Y(_05910_));
 AO221x1_ASAP7_75t_R _12827_ (.A1(_00630_),
    .A2(_03711_),
    .B1(_03874_),
    .B2(_03705_),
    .C(_05910_),
    .Y(_05911_));
 OAI21x1_ASAP7_75t_R _12828_ (.A1(_04602_),
    .A2(_05909_),
    .B(_05911_),
    .Y(_05912_));
 AND2x2_ASAP7_75t_R _12829_ (.A(_03610_),
    .B(_00629_),
    .Y(_05913_));
 AO21x1_ASAP7_75t_R _12830_ (.A1(_04831_),
    .A2(_00625_),
    .B(_05913_),
    .Y(_05914_));
 AO22x1_ASAP7_75t_R _12831_ (.A1(_00628_),
    .A2(_04800_),
    .B1(_05914_),
    .B2(_04597_),
    .Y(_05915_));
 NAND2x1_ASAP7_75t_R _12832_ (.A(_03815_),
    .B(_05915_),
    .Y(_05916_));
 AO21x1_ASAP7_75t_R _12833_ (.A1(_03825_),
    .A2(_05916_),
    .B(_04164_),
    .Y(_05917_));
 NAND2x1_ASAP7_75t_R _12834_ (.A(_00624_),
    .B(_03750_),
    .Y(_05918_));
 AO221x1_ASAP7_75t_R _12835_ (.A1(_03795_),
    .A2(_05912_),
    .B1(_05917_),
    .B2(_05918_),
    .C(_04468_),
    .Y(_05919_));
 AND3x1_ASAP7_75t_R _12836_ (.A(_04596_),
    .B(_04436_),
    .C(_00619_),
    .Y(_05920_));
 AO21x1_ASAP7_75t_R _12837_ (.A1(_00618_),
    .A2(_04595_),
    .B(_05920_),
    .Y(_05921_));
 AO222x2_ASAP7_75t_R _12838_ (.A1(_00616_),
    .A2(_03703_),
    .B1(_04628_),
    .B2(_00617_),
    .C1(_05921_),
    .C2(_03733_),
    .Y(_05922_));
 AOI21x1_ASAP7_75t_R _12839_ (.A1(_04915_),
    .A2(_05922_),
    .B(_03809_),
    .Y(_05923_));
 AND3x1_ASAP7_75t_R _12840_ (.A(_03815_),
    .B(_04930_),
    .C(_00607_),
    .Y(_05924_));
 AO21x1_ASAP7_75t_R _12841_ (.A1(_00606_),
    .A2(_04929_),
    .B(_05924_),
    .Y(_05925_));
 AND2x2_ASAP7_75t_R _12842_ (.A(_00602_),
    .B(_03890_),
    .Y(_05926_));
 AO221x1_ASAP7_75t_R _12843_ (.A1(_00603_),
    .A2(_04921_),
    .B1(_04804_),
    .B2(_03861_),
    .C(_05926_),
    .Y(_05927_));
 OA211x2_ASAP7_75t_R _12844_ (.A1(_00601_),
    .A2(_04952_),
    .B(_04627_),
    .C(_05927_),
    .Y(_05928_));
 AND3x1_ASAP7_75t_R _12845_ (.A(_03844_),
    .B(_05224_),
    .C(_00605_),
    .Y(_05929_));
 AO21x1_ASAP7_75t_R _12846_ (.A1(_00604_),
    .A2(_04434_),
    .B(_05929_),
    .Y(_05930_));
 AO21x1_ASAP7_75t_R _12847_ (.A1(_04727_),
    .A2(_05930_),
    .B(_04959_),
    .Y(_05931_));
 AOI211x1_ASAP7_75t_R _12848_ (.A1(_04440_),
    .A2(_05925_),
    .B(_05928_),
    .C(_05931_),
    .Y(_05932_));
 INVx1_ASAP7_75t_R _12849_ (.A(_00608_),
    .Y(_05933_));
 AND2x2_ASAP7_75t_R _12850_ (.A(_04610_),
    .B(_00613_),
    .Y(_05934_));
 AO21x1_ASAP7_75t_R _12851_ (.A1(_04457_),
    .A2(_00609_),
    .B(_05934_),
    .Y(_05935_));
 AOI22x1_ASAP7_75t_R _12852_ (.A1(_00612_),
    .A2(_04576_),
    .B1(_05935_),
    .B2(_03665_),
    .Y(_05936_));
 OA211x2_ASAP7_75t_R _12853_ (.A1(_03839_),
    .A2(_05936_),
    .B(_03775_),
    .C(_03737_),
    .Y(_05937_));
 OA22x2_ASAP7_75t_R _12854_ (.A1(_05933_),
    .A2(_04575_),
    .B1(_05937_),
    .B2(_03785_),
    .Y(_05938_));
 AND3x1_ASAP7_75t_R _12855_ (.A(_00611_),
    .B(_03705_),
    .C(_03874_),
    .Y(_05939_));
 AOI211x1_ASAP7_75t_R _12856_ (.A1(_00615_),
    .A2(_04602_),
    .B(_03869_),
    .C(_05939_),
    .Y(_05940_));
 AND3x1_ASAP7_75t_R _12857_ (.A(_00610_),
    .B(_03705_),
    .C(_03874_),
    .Y(_05941_));
 AOI211x1_ASAP7_75t_R _12858_ (.A1(_00614_),
    .A2(_04602_),
    .B(_03866_),
    .C(_05941_),
    .Y(_05942_));
 OR4x1_ASAP7_75t_R _12859_ (.A(_04468_),
    .B(_05938_),
    .C(_05940_),
    .D(_05942_),
    .Y(_05943_));
 AO32x2_ASAP7_75t_R _12860_ (.A1(_05907_),
    .A2(_05919_),
    .A3(_05923_),
    .B1(_05932_),
    .B2(_05943_),
    .Y(_05944_));
 BUFx16f_ASAP7_75t_R _12861_ (.A(_05944_),
    .Y(_10037_));
 INVx1_ASAP7_75t_R _12862_ (.A(_10037_),
    .Y(_10039_));
 NAND2x2_ASAP7_75t_R _12863_ (.A(_03382_),
    .B(_03534_),
    .Y(_05945_));
 INVx2_ASAP7_75t_R _12864_ (.A(_05945_),
    .Y(_05946_));
 AO32x1_ASAP7_75t_R _12865_ (.A1(_04171_),
    .A2(_04172_),
    .A3(_05853_),
    .B1(_05946_),
    .B2(_04848_),
    .Y(_05947_));
 OAI21x1_ASAP7_75t_R _12866_ (.A1(_05347_),
    .A2(_05947_),
    .B(_04168_),
    .Y(_05948_));
 INVx1_ASAP7_75t_R _12867_ (.A(_05948_),
    .Y(_05949_));
 OA211x2_ASAP7_75t_R _12868_ (.A1(_05347_),
    .A2(_05854_),
    .B(_04174_),
    .C(_04168_),
    .Y(_05950_));
 AO21x2_ASAP7_75t_R _12869_ (.A1(_05346_),
    .A2(_05949_),
    .B(_05950_),
    .Y(_10134_));
 AO22x1_ASAP7_75t_R _12870_ (.A1(_04502_),
    .A2(_00656_),
    .B1(_04069_),
    .B2(_00654_),
    .Y(_05951_));
 AND2x2_ASAP7_75t_R _12871_ (.A(_03957_),
    .B(_00655_),
    .Y(_05952_));
 AO21x1_ASAP7_75t_R _12872_ (.A1(_03955_),
    .A2(_00653_),
    .B(_05952_),
    .Y(_05953_));
 AO221x1_ASAP7_75t_R _12873_ (.A1(_04071_),
    .A2(_00653_),
    .B1(_05953_),
    .B2(_04265_),
    .C(_04156_),
    .Y(_05954_));
 AO21x1_ASAP7_75t_R _12874_ (.A1(_04066_),
    .A2(_05951_),
    .B(_05954_),
    .Y(_05955_));
 AND2x2_ASAP7_75t_R _12875_ (.A(_03926_),
    .B(_00663_),
    .Y(_05956_));
 AO21x1_ASAP7_75t_R _12876_ (.A1(_04104_),
    .A2(_00661_),
    .B(_05956_),
    .Y(_05957_));
 AO21x1_ASAP7_75t_R _12877_ (.A1(_00664_),
    .A2(_03962_),
    .B(_04009_),
    .Y(_05958_));
 AO221x1_ASAP7_75t_R _12878_ (.A1(_00662_),
    .A2(_04083_),
    .B1(_05957_),
    .B2(_04080_),
    .C(_05958_),
    .Y(_05959_));
 AO21x1_ASAP7_75t_R _12879_ (.A1(_05955_),
    .A2(_05959_),
    .B(_04095_),
    .Y(_05960_));
 AND3x1_ASAP7_75t_R _12880_ (.A(_04016_),
    .B(_04289_),
    .C(_00660_),
    .Y(_05961_));
 AND2x2_ASAP7_75t_R _12881_ (.A(_03957_),
    .B(_00659_),
    .Y(_05962_));
 AO21x1_ASAP7_75t_R _12882_ (.A1(_03955_),
    .A2(_00657_),
    .B(_05962_),
    .Y(_05963_));
 AO32x1_ASAP7_75t_R _12883_ (.A1(_04104_),
    .A2(_00658_),
    .A3(_04102_),
    .B1(_05963_),
    .B2(_03951_),
    .Y(_05964_));
 OR3x1_ASAP7_75t_R _12884_ (.A(_04514_),
    .B(_05961_),
    .C(_05964_),
    .Y(_05965_));
 AND2x2_ASAP7_75t_R _12885_ (.A(_04075_),
    .B(_00651_),
    .Y(_05966_));
 AO21x1_ASAP7_75t_R _12886_ (.A1(_04073_),
    .A2(_00649_),
    .B(_05966_),
    .Y(_05967_));
 AO32x1_ASAP7_75t_R _12887_ (.A1(_04521_),
    .A2(_00650_),
    .A3(_04522_),
    .B1(_05967_),
    .B2(_04088_),
    .Y(_05968_));
 AO221x1_ASAP7_75t_R _12888_ (.A1(_04112_),
    .A2(_03381_),
    .B1(_00652_),
    .B2(_04091_),
    .C(_05968_),
    .Y(_05969_));
 AO21x1_ASAP7_75t_R _12889_ (.A1(_05965_),
    .A2(_05969_),
    .B(_04120_),
    .Y(_05970_));
 AOI21x1_ASAP7_75t_R _12890_ (.A1(_05960_),
    .A2(_05970_),
    .B(_04122_),
    .Y(_05971_));
 AND2x2_ASAP7_75t_R _12891_ (.A(_04137_),
    .B(_00636_),
    .Y(_05972_));
 AO21x1_ASAP7_75t_R _12892_ (.A1(_04663_),
    .A2(_00635_),
    .B(_05972_),
    .Y(_05973_));
 AO21x1_ASAP7_75t_R _12893_ (.A1(_04502_),
    .A2(_05973_),
    .B(_04032_),
    .Y(_05974_));
 AO22x1_ASAP7_75t_R _12894_ (.A1(_04281_),
    .A2(_00633_),
    .B1(_00634_),
    .B2(_05073_),
    .Y(_05975_));
 AO22x2_ASAP7_75t_R _12895_ (.A1(_04504_),
    .A2(_00633_),
    .B1(_05975_),
    .B2(_04114_),
    .Y(_05976_));
 AO21x1_ASAP7_75t_R _12896_ (.A1(_04060_),
    .A2(_05974_),
    .B(_05976_),
    .Y(_05977_));
 AND2x2_ASAP7_75t_R _12897_ (.A(_04532_),
    .B(_00640_),
    .Y(_05978_));
 AO21x1_ASAP7_75t_R _12898_ (.A1(_04531_),
    .A2(_00639_),
    .B(_05978_),
    .Y(_05979_));
 AND3x1_ASAP7_75t_R _12899_ (.A(_04537_),
    .B(_03971_),
    .C(_00638_),
    .Y(_05980_));
 AO21x1_ASAP7_75t_R _12900_ (.A1(_00637_),
    .A2(_04535_),
    .B(_05980_),
    .Y(_05981_));
 AO221x1_ASAP7_75t_R _12901_ (.A1(_04530_),
    .A2(_05979_),
    .B1(_05981_),
    .B2(_04540_),
    .C(_04542_),
    .Y(_05982_));
 AND2x2_ASAP7_75t_R _12902_ (.A(_04532_),
    .B(_00648_),
    .Y(_05983_));
 AO21x1_ASAP7_75t_R _12903_ (.A1(_04531_),
    .A2(_00647_),
    .B(_05983_),
    .Y(_05984_));
 AND3x1_ASAP7_75t_R _12904_ (.A(_04537_),
    .B(_03971_),
    .C(_00646_),
    .Y(_05985_));
 AO21x1_ASAP7_75t_R _12905_ (.A1(_00645_),
    .A2(_04535_),
    .B(_05985_),
    .Y(_05986_));
 AO221x1_ASAP7_75t_R _12906_ (.A1(_04530_),
    .A2(_05984_),
    .B1(_05986_),
    .B2(_04540_),
    .C(_04542_),
    .Y(_05987_));
 AND2x2_ASAP7_75t_R _12907_ (.A(_04075_),
    .B(_00643_),
    .Y(_05988_));
 AO21x1_ASAP7_75t_R _12908_ (.A1(_04073_),
    .A2(_00641_),
    .B(_05988_),
    .Y(_05989_));
 AO22x1_ASAP7_75t_R _12909_ (.A1(_00644_),
    .A2(_04262_),
    .B1(_05989_),
    .B2(_04079_),
    .Y(_05990_));
 AO21x1_ASAP7_75t_R _12910_ (.A1(_00642_),
    .A2(_04983_),
    .B(_04130_),
    .Y(_05991_));
 OA21x2_ASAP7_75t_R _12911_ (.A1(_05990_),
    .A2(_05991_),
    .B(_03921_),
    .Y(_05992_));
 AO32x2_ASAP7_75t_R _12912_ (.A1(_04099_),
    .A2(_05977_),
    .A3(_05982_),
    .B1(_05987_),
    .B2(_05992_),
    .Y(_05993_));
 NOR2x1_ASAP7_75t_R _12913_ (.A(_04124_),
    .B(_05993_),
    .Y(_05994_));
 OAI21x1_ASAP7_75t_R _12914_ (.A1(_05971_),
    .A2(_05994_),
    .B(_03447_),
    .Y(_05995_));
 NAND2x1_ASAP7_75t_R _12915_ (.A(_05547_),
    .B(_05995_),
    .Y(_05996_));
 OA21x2_ASAP7_75t_R _12916_ (.A1(_05547_),
    .A2(_10134_),
    .B(_05996_),
    .Y(_05997_));
 XNOR2x1_ASAP7_75t_R _12917_ (.B(_05997_),
    .Y(_10043_),
    .A(_03913_));
 INVx1_ASAP7_75t_R _12918_ (.A(_10043_),
    .Y(_10045_));
 OR2x2_ASAP7_75t_R _12919_ (.A(_03816_),
    .B(_00654_),
    .Y(_05998_));
 OA211x2_ASAP7_75t_R _12920_ (.A1(_00656_),
    .A2(_04792_),
    .B(_05998_),
    .C(_05640_),
    .Y(_05999_));
 OA21x2_ASAP7_75t_R _12921_ (.A1(_00655_),
    .A2(_04792_),
    .B(_04623_),
    .Y(_06000_));
 OA211x2_ASAP7_75t_R _12922_ (.A1(_00653_),
    .A2(_04492_),
    .B(_04920_),
    .C(_03822_),
    .Y(_06001_));
 OAI21x1_ASAP7_75t_R _12923_ (.A1(_05999_),
    .A2(_06000_),
    .B(_06001_),
    .Y(_06002_));
 AND2x2_ASAP7_75t_R _12924_ (.A(_05332_),
    .B(_00662_),
    .Y(_06003_));
 AO21x1_ASAP7_75t_R _12925_ (.A1(_05331_),
    .A2(_00658_),
    .B(_06003_),
    .Y(_06004_));
 AO22x1_ASAP7_75t_R _12926_ (.A1(_00661_),
    .A2(_04936_),
    .B1(_06004_),
    .B2(_03798_),
    .Y(_06005_));
 NAND2x1_ASAP7_75t_R _12927_ (.A(_04053_),
    .B(_06005_),
    .Y(_06006_));
 AO21x1_ASAP7_75t_R _12928_ (.A1(_03826_),
    .A2(_06006_),
    .B(_03786_),
    .Y(_06007_));
 NAND2x1_ASAP7_75t_R _12929_ (.A(_00657_),
    .B(_03811_),
    .Y(_06008_));
 AND2x2_ASAP7_75t_R _12930_ (.A(_00663_),
    .B(_04434_),
    .Y(_06009_));
 AND2x2_ASAP7_75t_R _12931_ (.A(_00659_),
    .B(_03805_),
    .Y(_06010_));
 AO32x1_ASAP7_75t_R _12932_ (.A1(_03837_),
    .A2(_03838_),
    .A3(_06010_),
    .B1(_03834_),
    .B2(_00660_),
    .Y(_06011_));
 AOI221x1_ASAP7_75t_R _12933_ (.A1(_00664_),
    .A2(_05230_),
    .B1(_06009_),
    .B2(_03872_),
    .C(_06011_),
    .Y(_06012_));
 AO221x2_ASAP7_75t_R _12934_ (.A1(_06007_),
    .A2(_06008_),
    .B1(_06012_),
    .B2(_03852_),
    .C(_05235_),
    .Y(_06013_));
 AND3x1_ASAP7_75t_R _12935_ (.A(_03797_),
    .B(_03798_),
    .C(_00652_),
    .Y(_06014_));
 AO21x1_ASAP7_75t_R _12936_ (.A1(_00651_),
    .A2(_03796_),
    .B(_06014_),
    .Y(_06015_));
 AO222x2_ASAP7_75t_R _12937_ (.A1(_00649_),
    .A2(_03703_),
    .B1(_04628_),
    .B2(_00650_),
    .C1(_06015_),
    .C2(_03733_),
    .Y(_06016_));
 AOI21x1_ASAP7_75t_R _12938_ (.A1(_04915_),
    .A2(_06016_),
    .B(_03809_),
    .Y(_06017_));
 AND3x1_ASAP7_75t_R _12939_ (.A(_03969_),
    .B(_04624_),
    .C(_00640_),
    .Y(_06018_));
 AO21x1_ASAP7_75t_R _12940_ (.A1(_00639_),
    .A2(_04623_),
    .B(_06018_),
    .Y(_06019_));
 AND2x2_ASAP7_75t_R _12941_ (.A(_00635_),
    .B(_03714_),
    .Y(_06020_));
 AO221x1_ASAP7_75t_R _12942_ (.A1(_00636_),
    .A2(_03887_),
    .B1(_03803_),
    .B2(_03837_),
    .C(_06020_),
    .Y(_06021_));
 OA211x2_ASAP7_75t_R _12943_ (.A1(_00634_),
    .A2(_04952_),
    .B(_04627_),
    .C(_06021_),
    .Y(_06022_));
 AND3x1_ASAP7_75t_R _12944_ (.A(_03377_),
    .B(_04624_),
    .C(_00638_),
    .Y(_06023_));
 AO21x1_ASAP7_75t_R _12945_ (.A1(_00637_),
    .A2(_04623_),
    .B(_06023_),
    .Y(_06024_));
 AO21x1_ASAP7_75t_R _12946_ (.A1(_04727_),
    .A2(_06024_),
    .B(_04959_),
    .Y(_06025_));
 AOI211x1_ASAP7_75t_R _12947_ (.A1(_04440_),
    .A2(_06019_),
    .B(_06022_),
    .C(_06025_),
    .Y(_06026_));
 AND3x1_ASAP7_75t_R _12948_ (.A(_00643_),
    .B(_03837_),
    .C(_03838_),
    .Y(_06027_));
 AOI211x1_ASAP7_75t_R _12949_ (.A1(_00647_),
    .A2(_03872_),
    .B(_03866_),
    .C(_06027_),
    .Y(_06028_));
 AND3x1_ASAP7_75t_R _12950_ (.A(_00644_),
    .B(_03837_),
    .C(_03838_),
    .Y(_06029_));
 AOI211x1_ASAP7_75t_R _12951_ (.A1(_00648_),
    .A2(_03872_),
    .B(_03869_),
    .C(_06029_),
    .Y(_06030_));
 INVx1_ASAP7_75t_R _12952_ (.A(_00641_),
    .Y(_06031_));
 AND2x2_ASAP7_75t_R _12953_ (.A(_04938_),
    .B(_00646_),
    .Y(_06032_));
 AO21x1_ASAP7_75t_R _12954_ (.A1(_04831_),
    .A2(_00642_),
    .B(_06032_),
    .Y(_06033_));
 AOI22x1_ASAP7_75t_R _12955_ (.A1(_00645_),
    .A2(_05221_),
    .B1(_06033_),
    .B2(_05224_),
    .Y(_06034_));
 OA211x2_ASAP7_75t_R _12956_ (.A1(_05417_),
    .A2(_06034_),
    .B(_04592_),
    .C(_03873_),
    .Y(_06035_));
 OA22x2_ASAP7_75t_R _12957_ (.A1(_06031_),
    .A2(_04799_),
    .B1(_06035_),
    .B2(_05227_),
    .Y(_06036_));
 OR4x2_ASAP7_75t_R _12958_ (.A(_05235_),
    .B(_06028_),
    .C(_06030_),
    .D(_06036_),
    .Y(_06037_));
 AO32x2_ASAP7_75t_R _12959_ (.A1(_06002_),
    .A2(_06013_),
    .A3(_06017_),
    .B1(_06026_),
    .B2(_06037_),
    .Y(_06038_));
 BUFx10_ASAP7_75t_R _12960_ (.A(_06038_),
    .Y(_10042_));
 INVx3_ASAP7_75t_R _12961_ (.A(_10042_),
    .Y(_10044_));
 AND2x2_ASAP7_75t_R _12962_ (.A(_03932_),
    .B(_00669_),
    .Y(_06039_));
 AO21x1_ASAP7_75t_R _12963_ (.A1(_04037_),
    .A2(_00668_),
    .B(_06039_),
    .Y(_06040_));
 AO21x1_ASAP7_75t_R _12964_ (.A1(_04018_),
    .A2(_06040_),
    .B(_03966_),
    .Y(_06041_));
 AO22x1_ASAP7_75t_R _12965_ (.A1(_03949_),
    .A2(_00666_),
    .B1(_00667_),
    .B2(_03988_),
    .Y(_06042_));
 AO22x1_ASAP7_75t_R _12966_ (.A1(_04023_),
    .A2(_00666_),
    .B1(_06042_),
    .B2(_04113_),
    .Y(_06043_));
 AO21x1_ASAP7_75t_R _12967_ (.A1(_04142_),
    .A2(_06041_),
    .B(_06043_),
    .Y(_06044_));
 AND2x2_ASAP7_75t_R _12968_ (.A(_04014_),
    .B(_00673_),
    .Y(_06045_));
 AO21x1_ASAP7_75t_R _12969_ (.A1(_04274_),
    .A2(_00672_),
    .B(_06045_),
    .Y(_06046_));
 AND3x1_ASAP7_75t_R _12970_ (.A(_04403_),
    .B(_03970_),
    .C(_00671_),
    .Y(_06047_));
 AO21x1_ASAP7_75t_R _12971_ (.A1(_00670_),
    .A2(_04001_),
    .B(_06047_),
    .Y(_06048_));
 AO221x1_ASAP7_75t_R _12972_ (.A1(_04076_),
    .A2(_06046_),
    .B1(_06048_),
    .B2(_04004_),
    .C(_04541_),
    .Y(_06049_));
 AND2x2_ASAP7_75t_R _12973_ (.A(_04014_),
    .B(_00681_),
    .Y(_06050_));
 AO21x1_ASAP7_75t_R _12974_ (.A1(_03998_),
    .A2(_00680_),
    .B(_06050_),
    .Y(_06051_));
 AND3x1_ASAP7_75t_R _12975_ (.A(_04014_),
    .B(_03970_),
    .C(_00679_),
    .Y(_06052_));
 AO21x1_ASAP7_75t_R _12976_ (.A1(_00678_),
    .A2(_04001_),
    .B(_06052_),
    .Y(_06053_));
 AO221x1_ASAP7_75t_R _12977_ (.A1(_04076_),
    .A2(_06051_),
    .B1(_06053_),
    .B2(_04004_),
    .C(_03946_),
    .Y(_06054_));
 AND2x2_ASAP7_75t_R _12978_ (.A(_04025_),
    .B(_00676_),
    .Y(_06055_));
 AO21x1_ASAP7_75t_R _12979_ (.A1(_04024_),
    .A2(_00674_),
    .B(_06055_),
    .Y(_06056_));
 AO22x1_ASAP7_75t_R _12980_ (.A1(_00677_),
    .A2(_03960_),
    .B1(_06056_),
    .B2(_03986_),
    .Y(_06057_));
 AO21x1_ASAP7_75t_R _12981_ (.A1(_00675_),
    .A2(_04266_),
    .B(_03965_),
    .Y(_06058_));
 OA21x2_ASAP7_75t_R _12982_ (.A1(_06057_),
    .A2(_06058_),
    .B(_03920_),
    .Y(_06059_));
 AO32x1_ASAP7_75t_R _12983_ (.A1(_03997_),
    .A2(_06044_),
    .A3(_06049_),
    .B1(_06054_),
    .B2(_06059_),
    .Y(_06060_));
 AND2x2_ASAP7_75t_R _12984_ (.A(_04403_),
    .B(_00689_),
    .Y(_06061_));
 AO21x1_ASAP7_75t_R _12985_ (.A1(_03986_),
    .A2(_00688_),
    .B(_06061_),
    .Y(_06062_));
 AND3x1_ASAP7_75t_R _12986_ (.A(_04536_),
    .B(_04314_),
    .C(_00687_),
    .Y(_06063_));
 AO21x1_ASAP7_75t_R _12987_ (.A1(_00686_),
    .A2(_05590_),
    .B(_06063_),
    .Y(_06064_));
 AO221x1_ASAP7_75t_R _12988_ (.A1(_04529_),
    .A2(_06062_),
    .B1(_06064_),
    .B2(_04995_),
    .C(_04298_),
    .Y(_06065_));
 AND2x2_ASAP7_75t_R _12989_ (.A(_04403_),
    .B(_00697_),
    .Y(_06066_));
 AO21x1_ASAP7_75t_R _12990_ (.A1(_03986_),
    .A2(_00696_),
    .B(_06066_),
    .Y(_06067_));
 AND3x1_ASAP7_75t_R _12991_ (.A(_04536_),
    .B(_03970_),
    .C(_00695_),
    .Y(_06068_));
 AO21x1_ASAP7_75t_R _12992_ (.A1(_00694_),
    .A2(_05590_),
    .B(_06068_),
    .Y(_06069_));
 AO221x1_ASAP7_75t_R _12993_ (.A1(_04529_),
    .A2(_06067_),
    .B1(_06069_),
    .B2(_04004_),
    .C(_04304_),
    .Y(_06070_));
 AND3x1_ASAP7_75t_R _12994_ (.A(_04051_),
    .B(_06065_),
    .C(_06070_),
    .Y(_06071_));
 AO22x1_ASAP7_75t_R _12995_ (.A1(_03974_),
    .A2(_00685_),
    .B1(_04021_),
    .B2(_00683_),
    .Y(_06072_));
 AO221x1_ASAP7_75t_R _12996_ (.A1(_04075_),
    .A2(_00693_),
    .B1(_04021_),
    .B2(_00691_),
    .C(_03996_),
    .Y(_06073_));
 OA211x2_ASAP7_75t_R _12997_ (.A1(_04279_),
    .A2(_06072_),
    .B(_06073_),
    .C(_04127_),
    .Y(_06074_));
 AND2x2_ASAP7_75t_R _12998_ (.A(_04043_),
    .B(_00692_),
    .Y(_06075_));
 AO21x1_ASAP7_75t_R _12999_ (.A1(_04520_),
    .A2(_00690_),
    .B(_06075_),
    .Y(_06076_));
 AND2x2_ASAP7_75t_R _13000_ (.A(_03956_),
    .B(_00684_),
    .Y(_06077_));
 AO221x1_ASAP7_75t_R _13001_ (.A1(_04111_),
    .A2(_03379_),
    .B1(_00682_),
    .B2(_03954_),
    .C(_06077_),
    .Y(_06078_));
 OA211x2_ASAP7_75t_R _13002_ (.A1(_04097_),
    .A2(_06076_),
    .B(_06078_),
    .C(_04663_),
    .Y(_06079_));
 OR3x1_ASAP7_75t_R _13003_ (.A(_04119_),
    .B(_06074_),
    .C(_06079_),
    .Y(_06080_));
 AO221x2_ASAP7_75t_R _13004_ (.A1(_03916_),
    .A2(_06060_),
    .B1(_06071_),
    .B2(_06080_),
    .C(_04055_),
    .Y(_06081_));
 AO21x1_ASAP7_75t_R _13005_ (.A1(_04173_),
    .A2(_05946_),
    .B(_05347_),
    .Y(_06082_));
 NOR2x1_ASAP7_75t_R _13006_ (.A(_05346_),
    .B(_05948_),
    .Y(_06083_));
 AO21x2_ASAP7_75t_R _13007_ (.A1(_05346_),
    .A2(_06082_),
    .B(_06083_),
    .Y(_10132_));
 NAND2x1_ASAP7_75t_R _13008_ (.A(_04254_),
    .B(_10132_),
    .Y(_06084_));
 OA21x2_ASAP7_75t_R _13009_ (.A1(_04250_),
    .A2(_06081_),
    .B(_06084_),
    .Y(_06085_));
 XNOR2x1_ASAP7_75t_R _13010_ (.B(_06085_),
    .Y(_10048_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _13011_ (.A(_10048_),
    .Y(_10050_));
 AND3x1_ASAP7_75t_R _13012_ (.A(_00693_),
    .B(_04350_),
    .C(_03734_),
    .Y(_06086_));
 AOI211x1_ASAP7_75t_R _13013_ (.A1(_00697_),
    .A2(_03871_),
    .B(_06086_),
    .C(_03761_),
    .Y(_06087_));
 AND3x1_ASAP7_75t_R _13014_ (.A(_00692_),
    .B(_04350_),
    .C(_03734_),
    .Y(_06088_));
 AOI211x1_ASAP7_75t_R _13015_ (.A1(_00696_),
    .A2(_03871_),
    .B(_06088_),
    .C(_03886_),
    .Y(_06089_));
 OR4x1_ASAP7_75t_R _13016_ (.A(_03740_),
    .B(_03659_),
    .C(_06087_),
    .D(_06089_),
    .Y(_06090_));
 AND3x1_ASAP7_75t_R _13017_ (.A(_03443_),
    .B(_03716_),
    .C(_00689_),
    .Y(_06091_));
 AO21x1_ASAP7_75t_R _13018_ (.A1(_00688_),
    .A2(_03710_),
    .B(_06091_),
    .Y(_06092_));
 OA222x2_ASAP7_75t_R _13019_ (.A1(_00687_),
    .A2(_04952_),
    .B1(_06092_),
    .B2(_03824_),
    .C1(_04491_),
    .C2(_00686_),
    .Y(_06093_));
 AO221x2_ASAP7_75t_R _13020_ (.A1(_03554_),
    .A2(_03657_),
    .B1(_03570_),
    .B2(_03661_),
    .C(_03600_),
    .Y(_06094_));
 OA211x2_ASAP7_75t_R _13021_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03885_),
    .C(_00691_),
    .Y(_06095_));
 AOI21x1_ASAP7_75t_R _13022_ (.A1(_00690_),
    .A2(_03878_),
    .B(_06095_),
    .Y(_06096_));
 AO32x2_ASAP7_75t_R _13023_ (.A1(_03486_),
    .A2(_03489_),
    .A3(_03495_),
    .B1(_04610_),
    .B2(_03395_),
    .Y(_06097_));
 NAND2x1_ASAP7_75t_R _13024_ (.A(_00695_),
    .B(_03885_),
    .Y(_06098_));
 NAND2x1_ASAP7_75t_R _13025_ (.A(_00694_),
    .B(_03612_),
    .Y(_06099_));
 AND5x1_ASAP7_75t_R _13026_ (.A(_03509_),
    .B(_03516_),
    .C(_06097_),
    .D(_06098_),
    .E(_06099_),
    .Y(_06100_));
 NAND2x2_ASAP7_75t_R _13027_ (.A(_03775_),
    .B(_03697_),
    .Y(_06101_));
 AOI211x1_ASAP7_75t_R _13028_ (.A1(_06094_),
    .A2(_06096_),
    .B(_06100_),
    .C(_06101_),
    .Y(_06102_));
 INVx1_ASAP7_75t_R _13029_ (.A(_00684_),
    .Y(_06103_));
 INVx1_ASAP7_75t_R _13030_ (.A(_00683_),
    .Y(_06104_));
 NAND2x1_ASAP7_75t_R _13031_ (.A(_03619_),
    .B(_00685_),
    .Y(_06105_));
 OA211x2_ASAP7_75t_R _13032_ (.A1(_03636_),
    .A2(_06104_),
    .B(_06105_),
    .C(_03672_),
    .Y(_06106_));
 AOI21x1_ASAP7_75t_R _13033_ (.A1(_06103_),
    .A2(_04442_),
    .B(_06106_),
    .Y(_06107_));
 OA22x2_ASAP7_75t_R _13034_ (.A1(_00682_),
    .A2(_04344_),
    .B1(_06107_),
    .B2(_04811_),
    .Y(_06108_));
 AO21x1_ASAP7_75t_R _13035_ (.A1(_03772_),
    .A2(_06108_),
    .B(_03722_),
    .Y(_06109_));
 AOI211x1_ASAP7_75t_R _13036_ (.A1(_03791_),
    .A2(_06093_),
    .B(_06102_),
    .C(_06109_),
    .Y(_06110_));
 AND2x2_ASAP7_75t_R _13037_ (.A(_03608_),
    .B(_00679_),
    .Y(_06111_));
 AO21x1_ASAP7_75t_R _13038_ (.A1(_03683_),
    .A2(_00675_),
    .B(_06111_),
    .Y(_06112_));
 AO22x1_ASAP7_75t_R _13039_ (.A1(_00678_),
    .A2(_04210_),
    .B1(_06112_),
    .B2(_03716_),
    .Y(_06113_));
 NAND2x1_ASAP7_75t_R _13040_ (.A(_03639_),
    .B(_06113_),
    .Y(_06114_));
 AO21x1_ASAP7_75t_R _13041_ (.A1(_03824_),
    .A2(_06114_),
    .B(_04214_),
    .Y(_06115_));
 NAND2x1_ASAP7_75t_R _13042_ (.A(_00674_),
    .B(_03750_),
    .Y(_06116_));
 AND2x2_ASAP7_75t_R _13043_ (.A(_03614_),
    .B(_00681_),
    .Y(_06117_));
 AO21x1_ASAP7_75t_R _13044_ (.A1(_03629_),
    .A2(_00680_),
    .B(_06117_),
    .Y(_06118_));
 OA222x2_ASAP7_75t_R _13045_ (.A1(_03415_),
    .A2(_04457_),
    .B1(_00677_),
    .B2(_03709_),
    .C1(_04832_),
    .C2(_00676_),
    .Y(_06119_));
 AO21x1_ASAP7_75t_R _13046_ (.A1(_03670_),
    .A2(_06118_),
    .B(_06119_),
    .Y(_06120_));
 OR3x1_ASAP7_75t_R _13047_ (.A(_00676_),
    .B(_03657_),
    .C(_04204_),
    .Y(_06121_));
 OR4x1_ASAP7_75t_R _13048_ (.A(_00680_),
    .B(_04836_),
    .C(_03642_),
    .D(_03727_),
    .Y(_06122_));
 NAND3x1_ASAP7_75t_R _13049_ (.A(_06120_),
    .B(_06121_),
    .C(_06122_),
    .Y(_06123_));
 AO221x1_ASAP7_75t_R _13050_ (.A1(_06115_),
    .A2(_06116_),
    .B1(_06123_),
    .B2(_03733_),
    .C(_03740_),
    .Y(_06124_));
 OAI22x1_ASAP7_75t_R _13051_ (.A1(_00672_),
    .A2(_03881_),
    .B1(_03585_),
    .B2(_00673_),
    .Y(_06125_));
 AND2x2_ASAP7_75t_R _13052_ (.A(_03733_),
    .B(_06125_),
    .Y(_06126_));
 INVx1_ASAP7_75t_R _13053_ (.A(_00671_),
    .Y(_06127_));
 NAND2x1_ASAP7_75t_R _13054_ (.A(_00670_),
    .B(_03584_),
    .Y(_06128_));
 OA211x2_ASAP7_75t_R _13055_ (.A1(_06127_),
    .A2(_03585_),
    .B(_03658_),
    .C(_06128_),
    .Y(_06129_));
 AO221x1_ASAP7_75t_R _13056_ (.A1(_03510_),
    .A2(_03490_),
    .B1(_03402_),
    .B2(_03619_),
    .C(_00667_),
    .Y(_06130_));
 OA21x2_ASAP7_75t_R _13057_ (.A1(_00669_),
    .A2(_03593_),
    .B(_06130_),
    .Y(_06131_));
 OR3x1_ASAP7_75t_R _13058_ (.A(_03614_),
    .B(_03632_),
    .C(_00668_),
    .Y(_06132_));
 OR3x1_ASAP7_75t_R _13059_ (.A(_03618_),
    .B(_03636_),
    .C(_00667_),
    .Y(_06133_));
 AO21x1_ASAP7_75t_R _13060_ (.A1(_06132_),
    .A2(_06133_),
    .B(_03628_),
    .Y(_06134_));
 OA21x2_ASAP7_75t_R _13061_ (.A1(_03710_),
    .A2(_06131_),
    .B(_06134_),
    .Y(_06135_));
 AOI21x1_ASAP7_75t_R _13062_ (.A1(_03772_),
    .A2(_06135_),
    .B(_04194_),
    .Y(_06136_));
 OA31x2_ASAP7_75t_R _13063_ (.A1(_05698_),
    .A2(_06126_),
    .A3(_06129_),
    .B1(_06136_),
    .Y(_06137_));
 AO22x2_ASAP7_75t_R _13064_ (.A1(_06090_),
    .A2(_06110_),
    .B1(_06124_),
    .B2(_06137_),
    .Y(_06138_));
 BUFx6f_ASAP7_75t_R _13065_ (.A(_06138_),
    .Y(_10047_));
 INVx4_ASAP7_75t_R _13066_ (.A(_10047_),
    .Y(_10049_));
 INVx1_ASAP7_75t_R _13067_ (.A(_03504_),
    .Y(_06139_));
 AO21x2_ASAP7_75t_R _13068_ (.A1(_03382_),
    .A2(net28),
    .B(_03820_),
    .Y(_06140_));
 AND3x1_ASAP7_75t_R _13069_ (.A(_04174_),
    .B(_04168_),
    .C(_05347_),
    .Y(_06141_));
 AO221x2_ASAP7_75t_R _13070_ (.A1(_06139_),
    .A2(_06140_),
    .B1(_04102_),
    .B2(_04173_),
    .C(_06141_),
    .Y(_10130_));
 AO22x1_ASAP7_75t_R _13071_ (.A1(_04987_),
    .A2(_00722_),
    .B1(_04068_),
    .B2(_00720_),
    .Y(_06142_));
 AND2x2_ASAP7_75t_R _13072_ (.A(_03973_),
    .B(_00721_),
    .Y(_06143_));
 AO21x1_ASAP7_75t_R _13073_ (.A1(_03991_),
    .A2(_00719_),
    .B(_06143_),
    .Y(_06144_));
 AO221x1_ASAP7_75t_R _13074_ (.A1(_04023_),
    .A2(_00719_),
    .B1(_06144_),
    .B2(_03930_),
    .C(_04279_),
    .Y(_06145_));
 AO21x1_ASAP7_75t_R _13075_ (.A1(_04308_),
    .A2(_06142_),
    .B(_06145_),
    .Y(_06146_));
 AND2x2_ASAP7_75t_R _13076_ (.A(_03957_),
    .B(_00729_),
    .Y(_06147_));
 AO21x1_ASAP7_75t_R _13077_ (.A1(_03955_),
    .A2(_00727_),
    .B(_06147_),
    .Y(_06148_));
 AO21x1_ASAP7_75t_R _13078_ (.A1(_00730_),
    .A2(_03961_),
    .B(_04009_),
    .Y(_06149_));
 AO221x1_ASAP7_75t_R _13079_ (.A1(_00728_),
    .A2(_04983_),
    .B1(_06148_),
    .B2(_03951_),
    .C(_06149_),
    .Y(_06150_));
 AO21x1_ASAP7_75t_R _13080_ (.A1(_06146_),
    .A2(_06150_),
    .B(_04008_),
    .Y(_06151_));
 AND3x1_ASAP7_75t_R _13081_ (.A(_04034_),
    .B(_04076_),
    .C(_00726_),
    .Y(_06152_));
 AND2x2_ASAP7_75t_R _13082_ (.A(_03956_),
    .B(_00725_),
    .Y(_06153_));
 AO21x1_ASAP7_75t_R _13083_ (.A1(_04040_),
    .A2(_00723_),
    .B(_06153_),
    .Y(_06154_));
 AO32x1_ASAP7_75t_R _13084_ (.A1(_03955_),
    .A2(_00724_),
    .A3(_05073_),
    .B1(_06154_),
    .B2(_04281_),
    .Y(_06155_));
 OR3x1_ASAP7_75t_R _13085_ (.A(_03997_),
    .B(_06152_),
    .C(_06155_),
    .Y(_06156_));
 AND2x2_ASAP7_75t_R _13086_ (.A(_03956_),
    .B(_00717_),
    .Y(_06157_));
 AO21x1_ASAP7_75t_R _13087_ (.A1(_04040_),
    .A2(_00715_),
    .B(_06157_),
    .Y(_06158_));
 AO32x1_ASAP7_75t_R _13088_ (.A1(_04073_),
    .A2(_00716_),
    .A3(_05073_),
    .B1(_06158_),
    .B2(_04281_),
    .Y(_06159_));
 AO221x1_ASAP7_75t_R _13089_ (.A1(_04112_),
    .A2(_03972_),
    .B1(_00718_),
    .B2(_04262_),
    .C(_06159_),
    .Y(_06160_));
 AO21x1_ASAP7_75t_R _13090_ (.A1(_06156_),
    .A2(_06160_),
    .B(_04131_),
    .Y(_06161_));
 AO21x2_ASAP7_75t_R _13091_ (.A1(_06151_),
    .A2(_06161_),
    .B(_03917_),
    .Y(_06162_));
 AND2x2_ASAP7_75t_R _13092_ (.A(_03978_),
    .B(_00714_),
    .Y(_06163_));
 AO21x1_ASAP7_75t_R _13093_ (.A1(_03976_),
    .A2(_00713_),
    .B(_06163_),
    .Y(_06164_));
 AND3x1_ASAP7_75t_R _13094_ (.A(_04033_),
    .B(_04314_),
    .C(_00712_),
    .Y(_06165_));
 AO21x1_ASAP7_75t_R _13095_ (.A1(_00711_),
    .A2(_05590_),
    .B(_06165_),
    .Y(_06166_));
 AO221x1_ASAP7_75t_R _13096_ (.A1(_04270_),
    .A2(_06164_),
    .B1(_06166_),
    .B2(_04995_),
    .C(_04541_),
    .Y(_06167_));
 AND2x2_ASAP7_75t_R _13097_ (.A(_03925_),
    .B(_00709_),
    .Y(_06168_));
 AO21x1_ASAP7_75t_R _13098_ (.A1(_04113_),
    .A2(_00707_),
    .B(_06168_),
    .Y(_06169_));
 AO21x1_ASAP7_75t_R _13099_ (.A1(_00708_),
    .A2(_04266_),
    .B(_03966_),
    .Y(_06170_));
 AO221x1_ASAP7_75t_R _13100_ (.A1(_00710_),
    .A2(_04090_),
    .B1(_06169_),
    .B2(_04647_),
    .C(_06170_),
    .Y(_06171_));
 AND3x1_ASAP7_75t_R _13101_ (.A(_03921_),
    .B(_06167_),
    .C(_06171_),
    .Y(_06172_));
 AND2x2_ASAP7_75t_R _13102_ (.A(_03932_),
    .B(_00702_),
    .Y(_06173_));
 AO21x1_ASAP7_75t_R _13103_ (.A1(_03929_),
    .A2(_00701_),
    .B(_06173_),
    .Y(_06174_));
 AO21x1_ASAP7_75t_R _13104_ (.A1(_03926_),
    .A2(_06174_),
    .B(_03966_),
    .Y(_06175_));
 AND2x2_ASAP7_75t_R _13105_ (.A(_04142_),
    .B(_06175_),
    .Y(_06176_));
 AO22x1_ASAP7_75t_R _13106_ (.A1(_03976_),
    .A2(_00699_),
    .B1(_00700_),
    .B2(_04101_),
    .Y(_06177_));
 AO22x1_ASAP7_75t_R _13107_ (.A1(_04071_),
    .A2(_00699_),
    .B1(_06177_),
    .B2(_04521_),
    .Y(_06178_));
 AND2x2_ASAP7_75t_R _13108_ (.A(_04403_),
    .B(_00706_),
    .Y(_06179_));
 AO21x1_ASAP7_75t_R _13109_ (.A1(_03986_),
    .A2(_00705_),
    .B(_06179_),
    .Y(_06180_));
 AND3x1_ASAP7_75t_R _13110_ (.A(_04536_),
    .B(_03970_),
    .C(_00704_),
    .Y(_06181_));
 AO21x1_ASAP7_75t_R _13111_ (.A1(_00703_),
    .A2(_05590_),
    .B(_06181_),
    .Y(_06182_));
 AO221x1_ASAP7_75t_R _13112_ (.A1(_04529_),
    .A2(_06180_),
    .B1(_06182_),
    .B2(_04004_),
    .C(_04541_),
    .Y(_06183_));
 OA211x2_ASAP7_75t_R _13113_ (.A1(_06176_),
    .A2(_06178_),
    .B(_06183_),
    .C(_04098_),
    .Y(_06184_));
 OR3x1_ASAP7_75t_R _13114_ (.A(_04763_),
    .B(_06172_),
    .C(_06184_),
    .Y(_06185_));
 AOI21x1_ASAP7_75t_R _13115_ (.A1(_06162_),
    .A2(_06185_),
    .B(_04565_),
    .Y(_06186_));
 OR2x2_ASAP7_75t_R _13116_ (.A(_03915_),
    .B(_06186_),
    .Y(_06187_));
 OA21x2_ASAP7_75t_R _13117_ (.A1(_05547_),
    .A2(_10130_),
    .B(_06187_),
    .Y(_06188_));
 XNOR2x2_ASAP7_75t_R _13118_ (.A(_03913_),
    .B(_06188_),
    .Y(_10053_));
 INVx1_ASAP7_75t_R _13119_ (.A(_10053_),
    .Y(_10055_));
 AND2x2_ASAP7_75t_R _13120_ (.A(_03717_),
    .B(_00714_),
    .Y(_06189_));
 AO21x1_ASAP7_75t_R _13121_ (.A1(_03840_),
    .A2(_00713_),
    .B(_06189_),
    .Y(_06190_));
 OA222x2_ASAP7_75t_R _13122_ (.A1(_03839_),
    .A2(_05331_),
    .B1(_00710_),
    .B2(_04242_),
    .C1(_04832_),
    .C2(_00709_),
    .Y(_06191_));
 AO21x1_ASAP7_75t_R _13123_ (.A1(_03817_),
    .A2(_06190_),
    .B(_06191_),
    .Y(_06192_));
 OR3x1_ASAP7_75t_R _13124_ (.A(_00709_),
    .B(_03657_),
    .C(_04204_),
    .Y(_06193_));
 OR4x1_ASAP7_75t_R _13125_ (.A(_00713_),
    .B(_04836_),
    .C(_03642_),
    .D(_04921_),
    .Y(_06194_));
 AND3x1_ASAP7_75t_R _13126_ (.A(_06192_),
    .B(_06193_),
    .C(_06194_),
    .Y(_06195_));
 INVx1_ASAP7_75t_R _13127_ (.A(_00707_),
    .Y(_06196_));
 AND2x2_ASAP7_75t_R _13128_ (.A(_05332_),
    .B(_00712_),
    .Y(_06197_));
 AO21x1_ASAP7_75t_R _13129_ (.A1(_05331_),
    .A2(_00708_),
    .B(_06197_),
    .Y(_06198_));
 AOI22x1_ASAP7_75t_R _13130_ (.A1(_00711_),
    .A2(_04936_),
    .B1(_06198_),
    .B2(_04930_),
    .Y(_06199_));
 OA211x2_ASAP7_75t_R _13131_ (.A1(_04935_),
    .A2(_06199_),
    .B(_03803_),
    .C(_03804_),
    .Y(_06200_));
 OAI22x1_ASAP7_75t_R _13132_ (.A1(_06196_),
    .A2(_04934_),
    .B1(_06200_),
    .B2(_04165_),
    .Y(_06201_));
 OA21x2_ASAP7_75t_R _13133_ (.A1(_04583_),
    .A2(_06195_),
    .B(_06201_),
    .Y(_06202_));
 AND2x2_ASAP7_75t_R _13134_ (.A(_00700_),
    .B(_04583_),
    .Y(_06203_));
 AND2x2_ASAP7_75t_R _13135_ (.A(_00702_),
    .B(_03733_),
    .Y(_06204_));
 OA21x2_ASAP7_75t_R _13136_ (.A1(_00701_),
    .A2(_03866_),
    .B(_04627_),
    .Y(_06205_));
 OA33x2_ASAP7_75t_R _13137_ (.A1(_03587_),
    .A2(_06203_),
    .A3(_06204_),
    .B1(_06205_),
    .B2(_03600_),
    .B3(_04061_),
    .Y(_06206_));
 AO21x2_ASAP7_75t_R _13138_ (.A1(_04839_),
    .A2(_06202_),
    .B(_06206_),
    .Y(_06207_));
 AND3x1_ASAP7_75t_R _13139_ (.A(_04455_),
    .B(_04584_),
    .C(_00726_),
    .Y(_06208_));
 AO21x1_ASAP7_75t_R _13140_ (.A1(_00725_),
    .A2(_03891_),
    .B(_06208_),
    .Y(_06209_));
 AND3x1_ASAP7_75t_R _13141_ (.A(_03663_),
    .B(_03665_),
    .C(_00730_),
    .Y(_06210_));
 AO221x1_ASAP7_75t_R _13142_ (.A1(_00729_),
    .A2(_03714_),
    .B1(_03874_),
    .B2(_03861_),
    .C(_06210_),
    .Y(_06211_));
 OA21x2_ASAP7_75t_R _13143_ (.A1(_04602_),
    .A2(_06209_),
    .B(_06211_),
    .Y(_06212_));
 INVx1_ASAP7_75t_R _13144_ (.A(_00723_),
    .Y(_06213_));
 AND2x2_ASAP7_75t_R _13145_ (.A(_03610_),
    .B(_00728_),
    .Y(_06214_));
 AO21x1_ASAP7_75t_R _13146_ (.A1(_04831_),
    .A2(_00724_),
    .B(_06214_),
    .Y(_06215_));
 AOI22x1_ASAP7_75t_R _13147_ (.A1(_00727_),
    .A2(_05221_),
    .B1(_06215_),
    .B2(_05215_),
    .Y(_06216_));
 OA211x2_ASAP7_75t_R _13148_ (.A1(_05417_),
    .A2(_06216_),
    .B(_03888_),
    .C(_03873_),
    .Y(_06217_));
 OAI22x1_ASAP7_75t_R _13149_ (.A1(_06213_),
    .A2(_04799_),
    .B1(_06217_),
    .B2(_05227_),
    .Y(_06218_));
 OA211x2_ASAP7_75t_R _13150_ (.A1(_04792_),
    .A2(_06212_),
    .B(_06218_),
    .C(_03850_),
    .Y(_06219_));
 INVx1_ASAP7_75t_R _13151_ (.A(_00717_),
    .Y(_06220_));
 INVx1_ASAP7_75t_R _13152_ (.A(_00716_),
    .Y(_06221_));
 NAND2x1_ASAP7_75t_R _13153_ (.A(_03897_),
    .B(_00718_),
    .Y(_06222_));
 OA211x2_ASAP7_75t_R _13154_ (.A1(_03816_),
    .A2(_06221_),
    .B(_06222_),
    .C(_03762_),
    .Y(_06223_));
 AO21x1_ASAP7_75t_R _13155_ (.A1(_06220_),
    .A2(_04442_),
    .B(_06223_),
    .Y(_06224_));
 NAND2x1_ASAP7_75t_R _13156_ (.A(_03377_),
    .B(_06224_),
    .Y(_06225_));
 AO21x1_ASAP7_75t_R _13157_ (.A1(_03773_),
    .A2(_06225_),
    .B(_04806_),
    .Y(_06226_));
 OR2x2_ASAP7_75t_R _13158_ (.A(_00715_),
    .B(_03759_),
    .Y(_06227_));
 AO32x1_ASAP7_75t_R _13159_ (.A1(_00720_),
    .A2(_05640_),
    .A3(_03721_),
    .B1(_06226_),
    .B2(_06227_),
    .Y(_06228_));
 AND3x1_ASAP7_75t_R _13160_ (.A(_04596_),
    .B(_04436_),
    .C(_00722_),
    .Y(_06229_));
 AO21x1_ASAP7_75t_R _13161_ (.A1(_00721_),
    .A2(_04595_),
    .B(_06229_),
    .Y(_06230_));
 AO32x1_ASAP7_75t_R _13162_ (.A1(_00719_),
    .A2(_03862_),
    .A3(_03648_),
    .B1(_06230_),
    .B2(_03795_),
    .Y(_06231_));
 AO21x1_ASAP7_75t_R _13163_ (.A1(_03792_),
    .A2(_06231_),
    .B(_04499_),
    .Y(_06232_));
 OA211x2_ASAP7_75t_R _13164_ (.A1(_03524_),
    .A2(_03880_),
    .B(_03886_),
    .C(_00704_),
    .Y(_06233_));
 AO21x1_ASAP7_75t_R _13165_ (.A1(_00703_),
    .A2(_03586_),
    .B(_06233_),
    .Y(_06234_));
 OA222x2_ASAP7_75t_R _13166_ (.A1(_00705_),
    .A2(_03882_),
    .B1(_03586_),
    .B2(_00706_),
    .C1(_03783_),
    .C2(_03780_),
    .Y(_06235_));
 AO21x1_ASAP7_75t_R _13167_ (.A1(_03826_),
    .A2(_06234_),
    .B(_06235_),
    .Y(_06236_));
 AO21x1_ASAP7_75t_R _13168_ (.A1(_05403_),
    .A2(_06236_),
    .B(_03907_),
    .Y(_06237_));
 OA31x2_ASAP7_75t_R _13169_ (.A1(_06219_),
    .A2(_06228_),
    .A3(_06232_),
    .B1(_06237_),
    .Y(_06238_));
 OR2x2_ASAP7_75t_R _13170_ (.A(_06207_),
    .B(_06238_),
    .Y(_06239_));
 BUFx3_ASAP7_75t_R _13171_ (.A(_06239_),
    .Y(_10054_));
 AO22x1_ASAP7_75t_R _13172_ (.A1(_04076_),
    .A2(_00755_),
    .B1(_04068_),
    .B2(_00753_),
    .Y(_06240_));
 AND2x2_ASAP7_75t_R _13173_ (.A(_03956_),
    .B(_00754_),
    .Y(_06241_));
 AO21x1_ASAP7_75t_R _13174_ (.A1(_04040_),
    .A2(_00752_),
    .B(_06241_),
    .Y(_06242_));
 AO221x1_ASAP7_75t_R _13175_ (.A1(_04023_),
    .A2(_00752_),
    .B1(_06242_),
    .B2(_04281_),
    .C(_04279_),
    .Y(_06243_));
 AO21x1_ASAP7_75t_R _13176_ (.A1(_04308_),
    .A2(_06240_),
    .B(_06243_),
    .Y(_06244_));
 AND2x2_ASAP7_75t_R _13177_ (.A(_04105_),
    .B(_00762_),
    .Y(_06245_));
 AO21x1_ASAP7_75t_R _13178_ (.A1(_04103_),
    .A2(_00760_),
    .B(_06245_),
    .Y(_06246_));
 AO21x1_ASAP7_75t_R _13179_ (.A1(_00763_),
    .A2(_03961_),
    .B(_03413_),
    .Y(_06247_));
 AO221x1_ASAP7_75t_R _13180_ (.A1(_00761_),
    .A2(_03964_),
    .B1(_06246_),
    .B2(_04079_),
    .C(_06247_),
    .Y(_06248_));
 AO21x1_ASAP7_75t_R _13181_ (.A1(_06244_),
    .A2(_06248_),
    .B(_04008_),
    .Y(_06249_));
 AND3x1_ASAP7_75t_R _13182_ (.A(_04034_),
    .B(_03926_),
    .C(_00759_),
    .Y(_06250_));
 AND2x2_ASAP7_75t_R _13183_ (.A(_04025_),
    .B(_00758_),
    .Y(_06251_));
 AO21x1_ASAP7_75t_R _13184_ (.A1(_03954_),
    .A2(_00756_),
    .B(_06251_),
    .Y(_06252_));
 AO32x1_ASAP7_75t_R _13185_ (.A1(_04103_),
    .A2(_00757_),
    .A3(_04101_),
    .B1(_06252_),
    .B2(_03950_),
    .Y(_06253_));
 OR3x1_ASAP7_75t_R _13186_ (.A(_04414_),
    .B(_06250_),
    .C(_06253_),
    .Y(_06254_));
 AND2x2_ASAP7_75t_R _13187_ (.A(_04025_),
    .B(_00750_),
    .Y(_06255_));
 AO21x1_ASAP7_75t_R _13188_ (.A1(_03954_),
    .A2(_00748_),
    .B(_06255_),
    .Y(_06256_));
 AO32x1_ASAP7_75t_R _13189_ (.A1(_04113_),
    .A2(_00749_),
    .A3(_04101_),
    .B1(_06256_),
    .B2(_03976_),
    .Y(_06257_));
 AO221x1_ASAP7_75t_R _13190_ (.A1(_04111_),
    .A2(_04142_),
    .B1(_00751_),
    .B2(_04262_),
    .C(_06257_),
    .Y(_06258_));
 AO21x1_ASAP7_75t_R _13191_ (.A1(_06254_),
    .A2(_06258_),
    .B(_04131_),
    .Y(_06259_));
 AO21x1_ASAP7_75t_R _13192_ (.A1(_06249_),
    .A2(_06259_),
    .B(_03917_),
    .Y(_06260_));
 AND2x2_ASAP7_75t_R _13193_ (.A(_04403_),
    .B(_00747_),
    .Y(_06261_));
 AO21x1_ASAP7_75t_R _13194_ (.A1(_04028_),
    .A2(_00746_),
    .B(_06261_),
    .Y(_06262_));
 AND3x1_ASAP7_75t_R _13195_ (.A(_04536_),
    .B(_04314_),
    .C(_00745_),
    .Y(_06263_));
 AO21x1_ASAP7_75t_R _13196_ (.A1(_00744_),
    .A2(_05590_),
    .B(_06263_),
    .Y(_06264_));
 AO221x1_ASAP7_75t_R _13197_ (.A1(_04987_),
    .A2(_06262_),
    .B1(_06264_),
    .B2(_04995_),
    .C(_04541_),
    .Y(_06265_));
 AND2x2_ASAP7_75t_R _13198_ (.A(_04043_),
    .B(_00742_),
    .Y(_06266_));
 AO21x1_ASAP7_75t_R _13199_ (.A1(_04520_),
    .A2(_00740_),
    .B(_06266_),
    .Y(_06267_));
 AO21x1_ASAP7_75t_R _13200_ (.A1(_00741_),
    .A2(_03963_),
    .B(_03965_),
    .Y(_06268_));
 AO221x1_ASAP7_75t_R _13201_ (.A1(_00743_),
    .A2(_04090_),
    .B1(_06267_),
    .B2(_04671_),
    .C(_06268_),
    .Y(_06269_));
 AND3x1_ASAP7_75t_R _13202_ (.A(_04280_),
    .B(_06265_),
    .C(_06269_),
    .Y(_06270_));
 AO22x1_ASAP7_75t_R _13203_ (.A1(_04274_),
    .A2(_00732_),
    .B1(_00733_),
    .B2(_03989_),
    .Y(_06271_));
 AND2x2_ASAP7_75t_R _13204_ (.A(_03977_),
    .B(_00735_),
    .Y(_06272_));
 AO21x1_ASAP7_75t_R _13205_ (.A1(_03949_),
    .A2(_00734_),
    .B(_06272_),
    .Y(_06273_));
 AO21x1_ASAP7_75t_R _13206_ (.A1(_04544_),
    .A2(_06273_),
    .B(_03965_),
    .Y(_06274_));
 AND2x2_ASAP7_75t_R _13207_ (.A(_04023_),
    .B(_00732_),
    .Y(_06275_));
 AO221x1_ASAP7_75t_R _13208_ (.A1(_04276_),
    .A2(_06271_),
    .B1(_06274_),
    .B2(_03380_),
    .C(_06275_),
    .Y(_06276_));
 AND2x2_ASAP7_75t_R _13209_ (.A(_04403_),
    .B(_00739_),
    .Y(_06277_));
 AO21x1_ASAP7_75t_R _13210_ (.A1(_03986_),
    .A2(_00738_),
    .B(_06277_),
    .Y(_06278_));
 AND3x1_ASAP7_75t_R _13211_ (.A(_04536_),
    .B(_04314_),
    .C(_00737_),
    .Y(_06279_));
 AO21x1_ASAP7_75t_R _13212_ (.A1(_00736_),
    .A2(_05590_),
    .B(_06279_),
    .Y(_06280_));
 AO221x1_ASAP7_75t_R _13213_ (.A1(_04529_),
    .A2(_06278_),
    .B1(_06280_),
    .B2(_04995_),
    .C(_04541_),
    .Y(_06281_));
 AND3x1_ASAP7_75t_R _13214_ (.A(_04098_),
    .B(_06276_),
    .C(_06281_),
    .Y(_06282_));
 OR3x1_ASAP7_75t_R _13215_ (.A(_04763_),
    .B(_06270_),
    .C(_06282_),
    .Y(_06283_));
 AOI21x1_ASAP7_75t_R _13216_ (.A1(_06260_),
    .A2(_06283_),
    .B(_04055_),
    .Y(_06284_));
 BUFx10_ASAP7_75t_R _13217_ (.A(_03742_),
    .Y(_06285_));
 AND2x2_ASAP7_75t_R _13218_ (.A(_06285_),
    .B(_04169_),
    .Y(_10128_));
 AND2x2_ASAP7_75t_R _13219_ (.A(_04254_),
    .B(_10128_),
    .Y(_06286_));
 AOI21x1_ASAP7_75t_R _13220_ (.A1(_04065_),
    .A2(_06284_),
    .B(_06286_),
    .Y(_06287_));
 XNOR2x1_ASAP7_75t_R _13221_ (.B(_06287_),
    .Y(_10101_),
    .A(_03538_));
 INVx1_ASAP7_75t_R _13222_ (.A(_10101_),
    .Y(_10103_));
 AND3x1_ASAP7_75t_R _13223_ (.A(_04596_),
    .B(_04597_),
    .C(_00735_),
    .Y(_06288_));
 AO21x1_ASAP7_75t_R _13224_ (.A1(_00734_),
    .A2(_04595_),
    .B(_06288_),
    .Y(_06289_));
 AO222x2_ASAP7_75t_R _13225_ (.A1(_00732_),
    .A2(_04622_),
    .B1(_03901_),
    .B2(_06289_),
    .C1(_04629_),
    .C2(_00733_),
    .Y(_06290_));
 AO221x1_ASAP7_75t_R _13226_ (.A1(_00763_),
    .A2(_04198_),
    .B1(_03834_),
    .B2(_00759_),
    .C(_03825_),
    .Y(_06291_));
 AND3x1_ASAP7_75t_R _13227_ (.A(_00758_),
    .B(_03861_),
    .C(_03874_),
    .Y(_06292_));
 OA21x2_ASAP7_75t_R _13228_ (.A1(_03780_),
    .A2(_03817_),
    .B(_00762_),
    .Y(_06293_));
 OA21x2_ASAP7_75t_R _13229_ (.A1(_06292_),
    .A2(_06293_),
    .B(_03796_),
    .Y(_06294_));
 INVx1_ASAP7_75t_R _13230_ (.A(_00756_),
    .Y(_06295_));
 AND2x2_ASAP7_75t_R _13231_ (.A(_03610_),
    .B(_00761_),
    .Y(_06296_));
 AO21x1_ASAP7_75t_R _13232_ (.A1(_04831_),
    .A2(_00757_),
    .B(_06296_),
    .Y(_06297_));
 AOI22x1_ASAP7_75t_R _13233_ (.A1(_00760_),
    .A2(_04800_),
    .B1(_06297_),
    .B2(_04597_),
    .Y(_06298_));
 OA211x2_ASAP7_75t_R _13234_ (.A1(_03481_),
    .A2(_06298_),
    .B(_04804_),
    .C(_03861_),
    .Y(_06299_));
 OAI22x1_ASAP7_75t_R _13235_ (.A1(_06295_),
    .A2(_04799_),
    .B1(_06299_),
    .B2(_04806_),
    .Y(_06300_));
 OA211x2_ASAP7_75t_R _13236_ (.A1(_06291_),
    .A2(_06294_),
    .B(_03850_),
    .C(_06300_),
    .Y(_06301_));
 OA211x2_ASAP7_75t_R _13237_ (.A1(_03523_),
    .A2(_03696_),
    .B(_03881_),
    .C(_00753_),
    .Y(_06302_));
 AO21x1_ASAP7_75t_R _13238_ (.A1(_00752_),
    .A2(_03586_),
    .B(_06302_),
    .Y(_06303_));
 AND2x2_ASAP7_75t_R _13239_ (.A(_00754_),
    .B(_03890_),
    .Y(_06304_));
 AO221x1_ASAP7_75t_R _13240_ (.A1(_00755_),
    .A2(_04921_),
    .B1(_03888_),
    .B2(_03705_),
    .C(_06304_),
    .Y(_06305_));
 OA21x2_ASAP7_75t_R _13241_ (.A1(_03795_),
    .A2(_06303_),
    .B(_06305_),
    .Y(_06306_));
 AO21x2_ASAP7_75t_R _13242_ (.A1(_05403_),
    .A2(_06306_),
    .B(_04499_),
    .Y(_06307_));
 AND3x1_ASAP7_75t_R _13243_ (.A(_04916_),
    .B(_03853_),
    .C(_00751_),
    .Y(_06308_));
 AO21x1_ASAP7_75t_R _13244_ (.A1(_00750_),
    .A2(_03891_),
    .B(_06308_),
    .Y(_06309_));
 AO32x1_ASAP7_75t_R _13245_ (.A1(_03655_),
    .A2(_04587_),
    .A3(_06309_),
    .B1(_03702_),
    .B2(_00748_),
    .Y(_06310_));
 AND3x1_ASAP7_75t_R _13246_ (.A(_00749_),
    .B(_03814_),
    .C(_03889_),
    .Y(_06311_));
 OA21x2_ASAP7_75t_R _13247_ (.A1(_06310_),
    .A2(_06311_),
    .B(_04915_),
    .Y(_06312_));
 OA22x2_ASAP7_75t_R _13248_ (.A1(_00747_),
    .A2(_04478_),
    .B1(_04948_),
    .B2(_00743_),
    .Y(_06313_));
 OR2x2_ASAP7_75t_R _13249_ (.A(_00742_),
    .B(_04948_),
    .Y(_06314_));
 OA211x2_ASAP7_75t_R _13250_ (.A1(_00746_),
    .A2(_03836_),
    .B(_03761_),
    .C(_06314_),
    .Y(_06315_));
 AO21x1_ASAP7_75t_R _13251_ (.A1(_03887_),
    .A2(_06313_),
    .B(_06315_),
    .Y(_06316_));
 AND3x1_ASAP7_75t_R _13252_ (.A(_03715_),
    .B(_03717_),
    .C(_00747_),
    .Y(_06317_));
 AO21x1_ASAP7_75t_R _13253_ (.A1(_00746_),
    .A2(_03714_),
    .B(_06317_),
    .Y(_06318_));
 OA21x2_ASAP7_75t_R _13254_ (.A1(_03707_),
    .A2(_06318_),
    .B(_03698_),
    .Y(_06319_));
 INVx1_ASAP7_75t_R _13255_ (.A(_00740_),
    .Y(_06320_));
 AND2x2_ASAP7_75t_R _13256_ (.A(_04610_),
    .B(_00745_),
    .Y(_06321_));
 AO21x1_ASAP7_75t_R _13257_ (.A1(_04609_),
    .A2(_00741_),
    .B(_06321_),
    .Y(_06322_));
 AOI22x1_ASAP7_75t_R _13258_ (.A1(_00744_),
    .A2(_04800_),
    .B1(_06322_),
    .B2(_04584_),
    .Y(_06323_));
 OA211x2_ASAP7_75t_R _13259_ (.A1(_03481_),
    .A2(_06323_),
    .B(_04804_),
    .C(_04478_),
    .Y(_06324_));
 OAI22x1_ASAP7_75t_R _13260_ (.A1(_06320_),
    .A2(_04799_),
    .B1(_06324_),
    .B2(_04806_),
    .Y(_06325_));
 AND3x2_ASAP7_75t_R _13261_ (.A(_06316_),
    .B(_06319_),
    .C(_06325_),
    .Y(_06326_));
 AND4x1_ASAP7_75t_R _13262_ (.A(_00739_),
    .B(_03677_),
    .C(_03516_),
    .D(_03731_),
    .Y(_06327_));
 AO21x1_ASAP7_75t_R _13263_ (.A1(_00737_),
    .A2(_03659_),
    .B(_06327_),
    .Y(_06328_));
 OA22x2_ASAP7_75t_R _13264_ (.A1(_00736_),
    .A2(_04492_),
    .B1(_03866_),
    .B2(_00738_),
    .Y(_06329_));
 OA211x2_ASAP7_75t_R _13265_ (.A1(_03879_),
    .A2(_06328_),
    .B(_06329_),
    .C(_03791_),
    .Y(_06330_));
 OA33x2_ASAP7_75t_R _13266_ (.A1(_06301_),
    .A2(_06307_),
    .A3(_06312_),
    .B1(_06326_),
    .B2(_06330_),
    .B3(_04452_),
    .Y(_06331_));
 OR2x2_ASAP7_75t_R _13267_ (.A(_06290_),
    .B(_06331_),
    .Y(_06332_));
 BUFx6f_ASAP7_75t_R _13268_ (.A(_06332_),
    .Y(_10102_));
 AO22x1_ASAP7_75t_R _13269_ (.A1(_04529_),
    .A2(_00787_),
    .B1(_04068_),
    .B2(_00785_),
    .Y(_06333_));
 AND2x2_ASAP7_75t_R _13270_ (.A(_03973_),
    .B(_00786_),
    .Y(_06334_));
 AO21x1_ASAP7_75t_R _13271_ (.A1(_04040_),
    .A2(_00784_),
    .B(_06334_),
    .Y(_06335_));
 AO221x1_ASAP7_75t_R _13272_ (.A1(_04023_),
    .A2(_00784_),
    .B1(_06335_),
    .B2(_04281_),
    .C(_04279_),
    .Y(_06336_));
 AO21x1_ASAP7_75t_R _13273_ (.A1(_04308_),
    .A2(_06333_),
    .B(_06336_),
    .Y(_06337_));
 AND2x2_ASAP7_75t_R _13274_ (.A(_04075_),
    .B(_00794_),
    .Y(_06338_));
 AO21x1_ASAP7_75t_R _13275_ (.A1(_03955_),
    .A2(_00792_),
    .B(_06338_),
    .Y(_06339_));
 AO21x1_ASAP7_75t_R _13276_ (.A1(_00795_),
    .A2(_03961_),
    .B(_03413_),
    .Y(_06340_));
 AO221x1_ASAP7_75t_R _13277_ (.A1(_00793_),
    .A2(_04983_),
    .B1(_06339_),
    .B2(_03951_),
    .C(_06340_),
    .Y(_06341_));
 AO21x1_ASAP7_75t_R _13278_ (.A1(_06337_),
    .A2(_06341_),
    .B(_04008_),
    .Y(_06342_));
 AND3x1_ASAP7_75t_R _13279_ (.A(_04034_),
    .B(_04106_),
    .C(_00791_),
    .Y(_06343_));
 AND2x2_ASAP7_75t_R _13280_ (.A(_03956_),
    .B(_00790_),
    .Y(_06344_));
 AO21x1_ASAP7_75t_R _13281_ (.A1(_03954_),
    .A2(_00788_),
    .B(_06344_),
    .Y(_06345_));
 AO32x1_ASAP7_75t_R _13282_ (.A1(_04073_),
    .A2(_00789_),
    .A3(_05073_),
    .B1(_06345_),
    .B2(_03950_),
    .Y(_06346_));
 OR3x1_ASAP7_75t_R _13283_ (.A(_04414_),
    .B(_06343_),
    .C(_06346_),
    .Y(_06347_));
 AND2x2_ASAP7_75t_R _13284_ (.A(_04025_),
    .B(_00782_),
    .Y(_06348_));
 AO21x1_ASAP7_75t_R _13285_ (.A1(_03954_),
    .A2(_00780_),
    .B(_06348_),
    .Y(_06349_));
 AO32x1_ASAP7_75t_R _13286_ (.A1(_04103_),
    .A2(_00781_),
    .A3(_04101_),
    .B1(_06349_),
    .B2(_03950_),
    .Y(_06350_));
 AO221x1_ASAP7_75t_R _13287_ (.A1(_04112_),
    .A2(_03972_),
    .B1(_00783_),
    .B2(_04262_),
    .C(_06350_),
    .Y(_06351_));
 AO21x1_ASAP7_75t_R _13288_ (.A1(_06347_),
    .A2(_06351_),
    .B(_04131_),
    .Y(_06352_));
 AO21x2_ASAP7_75t_R _13289_ (.A1(_06342_),
    .A2(_06352_),
    .B(_03917_),
    .Y(_06353_));
 AND2x2_ASAP7_75t_R _13290_ (.A(_03978_),
    .B(_00779_),
    .Y(_06354_));
 AO21x1_ASAP7_75t_R _13291_ (.A1(_04028_),
    .A2(_00778_),
    .B(_06354_),
    .Y(_06355_));
 AND3x1_ASAP7_75t_R _13292_ (.A(_03978_),
    .B(_04314_),
    .C(_00777_),
    .Y(_06356_));
 AO21x1_ASAP7_75t_R _13293_ (.A1(_00776_),
    .A2(_05590_),
    .B(_06356_),
    .Y(_06357_));
 AO221x1_ASAP7_75t_R _13294_ (.A1(_04987_),
    .A2(_06355_),
    .B1(_06357_),
    .B2(_04995_),
    .C(_04541_),
    .Y(_06358_));
 AND2x2_ASAP7_75t_R _13295_ (.A(_04017_),
    .B(_00774_),
    .Y(_06359_));
 AO21x1_ASAP7_75t_R _13296_ (.A1(_04520_),
    .A2(_00772_),
    .B(_06359_),
    .Y(_06360_));
 AO21x1_ASAP7_75t_R _13297_ (.A1(_00773_),
    .A2(_04266_),
    .B(_03965_),
    .Y(_06361_));
 AO221x1_ASAP7_75t_R _13298_ (.A1(_00775_),
    .A2(_04090_),
    .B1(_06360_),
    .B2(_04556_),
    .C(_06361_),
    .Y(_06362_));
 AND3x1_ASAP7_75t_R _13299_ (.A(_04280_),
    .B(_06358_),
    .C(_06362_),
    .Y(_06363_));
 AO22x1_ASAP7_75t_R _13300_ (.A1(_04274_),
    .A2(_00764_),
    .B1(_00765_),
    .B2(_03989_),
    .Y(_06364_));
 AND2x2_ASAP7_75t_R _13301_ (.A(_03932_),
    .B(_00767_),
    .Y(_06365_));
 AO21x1_ASAP7_75t_R _13302_ (.A1(_04037_),
    .A2(_00766_),
    .B(_06365_),
    .Y(_06366_));
 AO21x1_ASAP7_75t_R _13303_ (.A1(_04544_),
    .A2(_06366_),
    .B(_03965_),
    .Y(_06367_));
 AND2x2_ASAP7_75t_R _13304_ (.A(_04023_),
    .B(_00764_),
    .Y(_06368_));
 AO221x1_ASAP7_75t_R _13305_ (.A1(_03992_),
    .A2(_06364_),
    .B1(_06367_),
    .B2(_04142_),
    .C(_06368_),
    .Y(_06369_));
 AND2x2_ASAP7_75t_R _13306_ (.A(_04536_),
    .B(_00771_),
    .Y(_06370_));
 AO21x1_ASAP7_75t_R _13307_ (.A1(_04028_),
    .A2(_00770_),
    .B(_06370_),
    .Y(_06371_));
 AND3x1_ASAP7_75t_R _13308_ (.A(_03978_),
    .B(_04314_),
    .C(_00769_),
    .Y(_06372_));
 AO21x1_ASAP7_75t_R _13309_ (.A1(_00768_),
    .A2(_05590_),
    .B(_06372_),
    .Y(_06373_));
 AO221x1_ASAP7_75t_R _13310_ (.A1(_04987_),
    .A2(_06371_),
    .B1(_06373_),
    .B2(_04995_),
    .C(_04541_),
    .Y(_06374_));
 AND3x1_ASAP7_75t_R _13311_ (.A(_04098_),
    .B(_06369_),
    .C(_06374_),
    .Y(_06375_));
 OR3x1_ASAP7_75t_R _13312_ (.A(_04763_),
    .B(_06363_),
    .C(_06375_),
    .Y(_06376_));
 AOI21x1_ASAP7_75t_R _13313_ (.A1(_06353_),
    .A2(_06376_),
    .B(_04565_),
    .Y(_06377_));
 AND3x2_ASAP7_75t_R _13314_ (.A(net89),
    .B(net20),
    .C(_06285_),
    .Y(_10126_));
 AND2x2_ASAP7_75t_R _13315_ (.A(_04254_),
    .B(_10126_),
    .Y(_06378_));
 AOI21x1_ASAP7_75t_R _13316_ (.A1(_04065_),
    .A2(_06377_),
    .B(_06378_),
    .Y(_06379_));
 XNOR2x2_ASAP7_75t_R _13317_ (.A(_03537_),
    .B(_06379_),
    .Y(_10058_));
 INVx1_ASAP7_75t_R _13318_ (.A(_10058_),
    .Y(_10060_));
 AND3x1_ASAP7_75t_R _13319_ (.A(_03715_),
    .B(_03717_),
    .C(_00769_),
    .Y(_06380_));
 AO22x1_ASAP7_75t_R _13320_ (.A1(_00768_),
    .A2(_03878_),
    .B1(_06380_),
    .B2(_03677_),
    .Y(_06381_));
 OA222x2_ASAP7_75t_R _13321_ (.A1(_00770_),
    .A2(_03886_),
    .B1(_03878_),
    .B2(_00771_),
    .C1(_03765_),
    .C2(_03667_),
    .Y(_06382_));
 AO21x1_ASAP7_75t_R _13322_ (.A1(_03825_),
    .A2(_06381_),
    .B(_06382_),
    .Y(_06383_));
 AO21x1_ASAP7_75t_R _13323_ (.A1(_05403_),
    .A2(_06383_),
    .B(_03907_),
    .Y(_06384_));
 AND3x1_ASAP7_75t_R _13324_ (.A(_00785_),
    .B(_04591_),
    .C(_04727_),
    .Y(_06385_));
 INVx1_ASAP7_75t_R _13325_ (.A(_00782_),
    .Y(_06386_));
 INVx1_ASAP7_75t_R _13326_ (.A(_00781_),
    .Y(_06387_));
 NAND2x1_ASAP7_75t_R _13327_ (.A(_03636_),
    .B(_00783_),
    .Y(_06388_));
 OA211x2_ASAP7_75t_R _13328_ (.A1(_03897_),
    .A2(_06387_),
    .B(_06388_),
    .C(_03672_),
    .Y(_06389_));
 AOI21x1_ASAP7_75t_R _13329_ (.A1(_06386_),
    .A2(_04442_),
    .B(_06389_),
    .Y(_06390_));
 OA211x2_ASAP7_75t_R _13330_ (.A1(_04811_),
    .A2(_06390_),
    .B(_03771_),
    .C(_03828_),
    .Y(_06391_));
 OA22x2_ASAP7_75t_R _13331_ (.A1(_00780_),
    .A2(_03759_),
    .B1(_06391_),
    .B2(_03785_),
    .Y(_06392_));
 AND3x1_ASAP7_75t_R _13332_ (.A(_03443_),
    .B(_03716_),
    .C(_00787_),
    .Y(_06393_));
 AO21x1_ASAP7_75t_R _13333_ (.A1(_00786_),
    .A2(_03671_),
    .B(_06393_),
    .Y(_06394_));
 OA21x2_ASAP7_75t_R _13334_ (.A1(_03667_),
    .A2(_03765_),
    .B(_06394_),
    .Y(_06395_));
 AND3x1_ASAP7_75t_R _13335_ (.A(_00784_),
    .B(_03828_),
    .C(_03648_),
    .Y(_06396_));
 OA211x2_ASAP7_75t_R _13336_ (.A1(_06395_),
    .A2(_06396_),
    .B(_03518_),
    .C(_03653_),
    .Y(_06397_));
 OR4x1_ASAP7_75t_R _13337_ (.A(_04499_),
    .B(_06385_),
    .C(_06392_),
    .D(_06397_),
    .Y(_06398_));
 AND3x1_ASAP7_75t_R _13338_ (.A(_04916_),
    .B(_03853_),
    .C(_00791_),
    .Y(_06399_));
 AO21x1_ASAP7_75t_R _13339_ (.A1(_00790_),
    .A2(_03891_),
    .B(_06399_),
    .Y(_06400_));
 AND3x1_ASAP7_75t_R _13340_ (.A(_03715_),
    .B(_03717_),
    .C(_00795_),
    .Y(_06401_));
 AO221x1_ASAP7_75t_R _13341_ (.A1(_00794_),
    .A2(_03805_),
    .B1(_03735_),
    .B2(_04478_),
    .C(_06401_),
    .Y(_06402_));
 OA21x2_ASAP7_75t_R _13342_ (.A1(_04602_),
    .A2(_06400_),
    .B(_06402_),
    .Y(_06403_));
 OA21x2_ASAP7_75t_R _13343_ (.A1(_04792_),
    .A2(_06403_),
    .B(_03850_),
    .Y(_06404_));
 INVx1_ASAP7_75t_R _13344_ (.A(_00788_),
    .Y(_06405_));
 AND2x2_ASAP7_75t_R _13345_ (.A(_04610_),
    .B(_00793_),
    .Y(_06406_));
 AO21x1_ASAP7_75t_R _13346_ (.A1(_04609_),
    .A2(_00789_),
    .B(_06406_),
    .Y(_06407_));
 AOI22x1_ASAP7_75t_R _13347_ (.A1(_00792_),
    .A2(_04800_),
    .B1(_06407_),
    .B2(_04584_),
    .Y(_06408_));
 OA211x2_ASAP7_75t_R _13348_ (.A1(_03481_),
    .A2(_06408_),
    .B(_03802_),
    .C(_04478_),
    .Y(_06409_));
 OAI22x1_ASAP7_75t_R _13349_ (.A1(_06405_),
    .A2(_04799_),
    .B1(_06409_),
    .B2(_04806_),
    .Y(_06410_));
 AO21x1_ASAP7_75t_R _13350_ (.A1(_03518_),
    .A2(_04920_),
    .B(_03906_),
    .Y(_06411_));
 OA211x2_ASAP7_75t_R _13351_ (.A1(_03907_),
    .A2(_06383_),
    .B(_06410_),
    .C(_06411_),
    .Y(_06412_));
 INVx1_ASAP7_75t_R _13352_ (.A(_00772_),
    .Y(_06413_));
 AND2x2_ASAP7_75t_R _13353_ (.A(_03610_),
    .B(_00777_),
    .Y(_06414_));
 AO21x1_ASAP7_75t_R _13354_ (.A1(_04831_),
    .A2(_00773_),
    .B(_06414_),
    .Y(_06415_));
 AOI22x1_ASAP7_75t_R _13355_ (.A1(_00776_),
    .A2(_04800_),
    .B1(_06415_),
    .B2(_04436_),
    .Y(_06416_));
 OA211x2_ASAP7_75t_R _13356_ (.A1(_03481_),
    .A2(_06416_),
    .B(_03888_),
    .C(_03705_),
    .Y(_06417_));
 OAI22x1_ASAP7_75t_R _13357_ (.A1(_06413_),
    .A2(_04799_),
    .B1(_06417_),
    .B2(_05227_),
    .Y(_06418_));
 AND2x2_ASAP7_75t_R _13358_ (.A(_04435_),
    .B(_00779_),
    .Y(_06419_));
 AO21x1_ASAP7_75t_R _13359_ (.A1(_03629_),
    .A2(_00778_),
    .B(_06419_),
    .Y(_06420_));
 OA222x2_ASAP7_75t_R _13360_ (.A1(_04811_),
    .A2(_04937_),
    .B1(_00775_),
    .B2(_03710_),
    .C1(_04832_),
    .C2(_00774_),
    .Y(_06421_));
 AO21x1_ASAP7_75t_R _13361_ (.A1(_03817_),
    .A2(_06420_),
    .B(_06421_),
    .Y(_06422_));
 OR3x1_ASAP7_75t_R _13362_ (.A(_00774_),
    .B(_03657_),
    .C(_04204_),
    .Y(_06423_));
 OR4x1_ASAP7_75t_R _13363_ (.A(_00778_),
    .B(_04836_),
    .C(_03642_),
    .D(_03886_),
    .Y(_06424_));
 AO31x2_ASAP7_75t_R _13364_ (.A1(_06422_),
    .A2(_06423_),
    .A3(_06424_),
    .B(_03659_),
    .Y(_06425_));
 AND4x1_ASAP7_75t_R _13365_ (.A(_00767_),
    .B(_03677_),
    .C(_03678_),
    .D(_03731_),
    .Y(_06426_));
 AO211x2_ASAP7_75t_R _13366_ (.A1(_00765_),
    .A2(_03659_),
    .B(_06426_),
    .C(_03879_),
    .Y(_06427_));
 AO221x1_ASAP7_75t_R _13367_ (.A1(_03376_),
    .A2(_05224_),
    .B1(_04478_),
    .B2(_04804_),
    .C(_00766_),
    .Y(_06428_));
 AO21x1_ASAP7_75t_R _13368_ (.A1(_04627_),
    .A2(_06428_),
    .B(_04806_),
    .Y(_06429_));
 AO32x1_ASAP7_75t_R _13369_ (.A1(_04839_),
    .A2(_06418_),
    .A3(_06425_),
    .B1(_06427_),
    .B2(_06429_),
    .Y(_06430_));
 AO221x2_ASAP7_75t_R _13370_ (.A1(_06384_),
    .A2(_06398_),
    .B1(_06404_),
    .B2(_06412_),
    .C(_06430_),
    .Y(_06431_));
 BUFx10_ASAP7_75t_R _13371_ (.A(_06431_),
    .Y(_10059_));
 AND2x2_ASAP7_75t_R _13372_ (.A(_04043_),
    .B(_00816_),
    .Y(_06432_));
 AO21x1_ASAP7_75t_R _13373_ (.A1(_03991_),
    .A2(_00814_),
    .B(_06432_),
    .Y(_06433_));
 AO222x2_ASAP7_75t_R _13374_ (.A1(_00817_),
    .A2(_03961_),
    .B1(_04266_),
    .B2(_00815_),
    .C1(_04663_),
    .C2(_06433_),
    .Y(_06434_));
 OR3x1_ASAP7_75t_R _13375_ (.A(_04119_),
    .B(_04280_),
    .C(_06434_),
    .Y(_06435_));
 AO22x1_ASAP7_75t_R _13376_ (.A1(_04643_),
    .A2(_00821_),
    .B1(_04632_),
    .B2(_00819_),
    .Y(_06436_));
 AND2x2_ASAP7_75t_R _13377_ (.A(_03957_),
    .B(_00820_),
    .Y(_06437_));
 AO21x1_ASAP7_75t_R _13378_ (.A1(_03955_),
    .A2(_00818_),
    .B(_06437_),
    .Y(_06438_));
 AO21x1_ASAP7_75t_R _13379_ (.A1(_03951_),
    .A2(_06438_),
    .B(_04298_),
    .Y(_06439_));
 AO21x1_ASAP7_75t_R _13380_ (.A1(_04308_),
    .A2(_06436_),
    .B(_06439_),
    .Y(_06440_));
 AND2x2_ASAP7_75t_R _13381_ (.A(_03926_),
    .B(_00828_),
    .Y(_06441_));
 AO21x1_ASAP7_75t_R _13382_ (.A1(_04114_),
    .A2(_00826_),
    .B(_06441_),
    .Y(_06442_));
 AO221x1_ASAP7_75t_R _13383_ (.A1(_00829_),
    .A2(_04090_),
    .B1(_03964_),
    .B2(_00827_),
    .C(_04304_),
    .Y(_06443_));
 AO21x1_ASAP7_75t_R _13384_ (.A1(_04080_),
    .A2(_06442_),
    .B(_06443_),
    .Y(_06444_));
 AND2x2_ASAP7_75t_R _13385_ (.A(_03973_),
    .B(_00824_),
    .Y(_06445_));
 AO21x1_ASAP7_75t_R _13386_ (.A1(_03991_),
    .A2(_00822_),
    .B(_06445_),
    .Y(_06446_));
 AO222x2_ASAP7_75t_R _13387_ (.A1(_00825_),
    .A2(_03961_),
    .B1(_04266_),
    .B2(_00823_),
    .C1(_03930_),
    .C2(_06446_),
    .Y(_06447_));
 OR3x1_ASAP7_75t_R _13388_ (.A(_04119_),
    .B(_03997_),
    .C(_06447_),
    .Y(_06448_));
 AND4x2_ASAP7_75t_R _13389_ (.A(_06435_),
    .B(_06440_),
    .C(_06444_),
    .D(_06448_),
    .Y(_06449_));
 AND2x2_ASAP7_75t_R _13390_ (.A(_03942_),
    .B(_00801_),
    .Y(_06450_));
 AO21x1_ASAP7_75t_R _13391_ (.A1(_04663_),
    .A2(_00800_),
    .B(_06450_),
    .Y(_06451_));
 AO21x1_ASAP7_75t_R _13392_ (.A1(_04502_),
    .A2(_06451_),
    .B(_04032_),
    .Y(_06452_));
 AO22x1_ASAP7_75t_R _13393_ (.A1(_04281_),
    .A2(_00798_),
    .B1(_00799_),
    .B2(_05073_),
    .Y(_06453_));
 AO22x1_ASAP7_75t_R _13394_ (.A1(_04504_),
    .A2(_00798_),
    .B1(_06453_),
    .B2(_04104_),
    .Y(_06454_));
 AO21x1_ASAP7_75t_R _13395_ (.A1(_04060_),
    .A2(_06452_),
    .B(_06454_),
    .Y(_06455_));
 AND2x2_ASAP7_75t_R _13396_ (.A(_04537_),
    .B(_00805_),
    .Y(_06456_));
 AO21x1_ASAP7_75t_R _13397_ (.A1(_04647_),
    .A2(_00804_),
    .B(_06456_),
    .Y(_06457_));
 AND3x1_ASAP7_75t_R _13398_ (.A(_04992_),
    .B(_03971_),
    .C(_00803_),
    .Y(_06458_));
 AO21x1_ASAP7_75t_R _13399_ (.A1(_00802_),
    .A2(_04991_),
    .B(_06458_),
    .Y(_06459_));
 AO221x1_ASAP7_75t_R _13400_ (.A1(_04988_),
    .A2(_06457_),
    .B1(_06459_),
    .B2(_04996_),
    .C(_04542_),
    .Y(_06460_));
 AND2x2_ASAP7_75t_R _13401_ (.A(_04532_),
    .B(_00813_),
    .Y(_06461_));
 AO21x1_ASAP7_75t_R _13402_ (.A1(_04531_),
    .A2(_00812_),
    .B(_06461_),
    .Y(_06462_));
 AND3x1_ASAP7_75t_R _13403_ (.A(_04537_),
    .B(_03971_),
    .C(_00811_),
    .Y(_06463_));
 AO21x1_ASAP7_75t_R _13404_ (.A1(_00810_),
    .A2(_04535_),
    .B(_06463_),
    .Y(_06464_));
 AO221x1_ASAP7_75t_R _13405_ (.A1(_04530_),
    .A2(_06462_),
    .B1(_06464_),
    .B2(_04540_),
    .C(_04542_),
    .Y(_06465_));
 AND2x2_ASAP7_75t_R _13406_ (.A(_04075_),
    .B(_00808_),
    .Y(_06466_));
 AO21x1_ASAP7_75t_R _13407_ (.A1(_04073_),
    .A2(_00806_),
    .B(_06466_),
    .Y(_06467_));
 AO22x1_ASAP7_75t_R _13408_ (.A1(_00809_),
    .A2(_04262_),
    .B1(_06467_),
    .B2(_04088_),
    .Y(_06468_));
 AO21x1_ASAP7_75t_R _13409_ (.A1(_00807_),
    .A2(_04983_),
    .B(_04130_),
    .Y(_06469_));
 OA21x2_ASAP7_75t_R _13410_ (.A1(_06468_),
    .A2(_06469_),
    .B(_03921_),
    .Y(_06470_));
 AO32x2_ASAP7_75t_R _13411_ (.A1(_04099_),
    .A2(_06455_),
    .A3(_06460_),
    .B1(_06465_),
    .B2(_06470_),
    .Y(_06471_));
 OAI22x1_ASAP7_75t_R _13412_ (.A1(_04122_),
    .A2(_06449_),
    .B1(_06471_),
    .B2(_04429_),
    .Y(_06472_));
 AND3x2_ASAP7_75t_R _13413_ (.A(net89),
    .B(net19),
    .C(_06285_),
    .Y(_10124_));
 AND2x2_ASAP7_75t_R _13414_ (.A(_04162_),
    .B(_10124_),
    .Y(_06473_));
 AOI21x1_ASAP7_75t_R _13415_ (.A1(_04065_),
    .A2(_06472_),
    .B(_06473_),
    .Y(_06474_));
 XNOR2x2_ASAP7_75t_R _13416_ (.A(_03537_),
    .B(_06474_),
    .Y(_10063_));
 INVx1_ASAP7_75t_R _13417_ (.A(_10063_),
    .Y(_10065_));
 AND2x2_ASAP7_75t_R _13418_ (.A(_00802_),
    .B(_03878_),
    .Y(_06475_));
 AND2x2_ASAP7_75t_R _13419_ (.A(_00803_),
    .B(_03813_),
    .Y(_06476_));
 OR4x2_ASAP7_75t_R _13420_ (.A(_03794_),
    .B(_03906_),
    .C(_06475_),
    .D(_06476_),
    .Y(_06477_));
 AND2x2_ASAP7_75t_R _13421_ (.A(_00804_),
    .B(_03710_),
    .Y(_06478_));
 AO221x1_ASAP7_75t_R _13422_ (.A1(_00805_),
    .A2(_03886_),
    .B1(_03802_),
    .B2(_03836_),
    .C(_06478_),
    .Y(_06479_));
 AO32x2_ASAP7_75t_R _13423_ (.A1(_03655_),
    .A2(_04920_),
    .A3(_06479_),
    .B1(_03905_),
    .B2(_03742_),
    .Y(_06480_));
 AND2x2_ASAP7_75t_R _13424_ (.A(_06477_),
    .B(_06480_),
    .Y(_06481_));
 OR2x2_ASAP7_75t_R _13425_ (.A(_00814_),
    .B(_03759_),
    .Y(_06482_));
 INVx1_ASAP7_75t_R _13426_ (.A(_00816_),
    .Y(_06483_));
 INVx1_ASAP7_75t_R _13427_ (.A(_00815_),
    .Y(_06484_));
 NAND2x1_ASAP7_75t_R _13428_ (.A(_03897_),
    .B(_00817_),
    .Y(_06485_));
 OA211x2_ASAP7_75t_R _13429_ (.A1(_03897_),
    .A2(_06484_),
    .B(_06485_),
    .C(_04435_),
    .Y(_06486_));
 AO21x1_ASAP7_75t_R _13430_ (.A1(_06483_),
    .A2(_04442_),
    .B(_06486_),
    .Y(_06487_));
 NAND2x1_ASAP7_75t_R _13431_ (.A(_03815_),
    .B(_06487_),
    .Y(_06488_));
 AO221x1_ASAP7_75t_R _13432_ (.A1(_00819_),
    .A2(_05497_),
    .B1(_06488_),
    .B2(_03773_),
    .C(_04164_),
    .Y(_06489_));
 AND3x1_ASAP7_75t_R _13433_ (.A(_04455_),
    .B(_04597_),
    .C(_00821_),
    .Y(_06490_));
 AO21x1_ASAP7_75t_R _13434_ (.A1(_00820_),
    .A2(_03782_),
    .B(_06490_),
    .Y(_06491_));
 AO32x1_ASAP7_75t_R _13435_ (.A1(_00818_),
    .A2(_03862_),
    .A3(_03648_),
    .B1(_06491_),
    .B2(_03795_),
    .Y(_06492_));
 AO221x1_ASAP7_75t_R _13436_ (.A1(_06482_),
    .A2(_06489_),
    .B1(_06492_),
    .B2(_05403_),
    .C(_04499_),
    .Y(_06493_));
 AND2x2_ASAP7_75t_R _13437_ (.A(_00828_),
    .B(_03890_),
    .Y(_06494_));
 AO221x1_ASAP7_75t_R _13438_ (.A1(_00829_),
    .A2(_04921_),
    .B1(_03874_),
    .B2(_03861_),
    .C(_06494_),
    .Y(_06495_));
 AND3x1_ASAP7_75t_R _13439_ (.A(_03375_),
    .B(_04460_),
    .C(_00825_),
    .Y(_06496_));
 AO21x1_ASAP7_75t_R _13440_ (.A1(_00824_),
    .A2(_04242_),
    .B(_06496_),
    .Y(_06497_));
 OR3x1_ASAP7_75t_R _13441_ (.A(_03780_),
    .B(_03817_),
    .C(_06497_),
    .Y(_06498_));
 AO21x1_ASAP7_75t_R _13442_ (.A1(_06495_),
    .A2(_06498_),
    .B(_05218_),
    .Y(_06499_));
 INVx1_ASAP7_75t_R _13443_ (.A(_00822_),
    .Y(_06500_));
 AND2x2_ASAP7_75t_R _13444_ (.A(_04938_),
    .B(_00827_),
    .Y(_06501_));
 AO21x1_ASAP7_75t_R _13445_ (.A1(_04831_),
    .A2(_00823_),
    .B(_06501_),
    .Y(_06502_));
 AOI22x1_ASAP7_75t_R _13446_ (.A1(_00826_),
    .A2(_05221_),
    .B1(_06502_),
    .B2(_05224_),
    .Y(_06503_));
 OA211x2_ASAP7_75t_R _13447_ (.A1(_05417_),
    .A2(_06503_),
    .B(_04592_),
    .C(_03873_),
    .Y(_06504_));
 OAI22x1_ASAP7_75t_R _13448_ (.A1(_06500_),
    .A2(_04934_),
    .B1(_06504_),
    .B2(_05227_),
    .Y(_06505_));
 AND5x1_ASAP7_75t_R _13449_ (.A(_03850_),
    .B(_06477_),
    .C(_06480_),
    .D(_06499_),
    .E(_06505_),
    .Y(_06506_));
 INVx1_ASAP7_75t_R _13450_ (.A(_00806_),
    .Y(_06507_));
 AND2x2_ASAP7_75t_R _13451_ (.A(_05332_),
    .B(_00811_),
    .Y(_06508_));
 AO21x1_ASAP7_75t_R _13452_ (.A1(_05331_),
    .A2(_00807_),
    .B(_06508_),
    .Y(_06509_));
 AOI22x1_ASAP7_75t_R _13453_ (.A1(_00810_),
    .A2(_04936_),
    .B1(_06509_),
    .B2(_04930_),
    .Y(_06510_));
 OA211x2_ASAP7_75t_R _13454_ (.A1(_04935_),
    .A2(_06510_),
    .B(_03803_),
    .C(_03804_),
    .Y(_06511_));
 OAI22x1_ASAP7_75t_R _13455_ (.A1(_06507_),
    .A2(_04934_),
    .B1(_06511_),
    .B2(_04165_),
    .Y(_06512_));
 NAND2x1_ASAP7_75t_R _13456_ (.A(_00813_),
    .B(_03774_),
    .Y(_06513_));
 NAND2x1_ASAP7_75t_R _13457_ (.A(_00812_),
    .B(_03891_),
    .Y(_06514_));
 AOI22x1_ASAP7_75t_R _13458_ (.A1(_03837_),
    .A2(_03838_),
    .B1(_06513_),
    .B2(_06514_),
    .Y(_06515_));
 AND2x2_ASAP7_75t_R _13459_ (.A(_00808_),
    .B(_04242_),
    .Y(_06516_));
 AO32x1_ASAP7_75t_R _13460_ (.A1(_03829_),
    .A2(_03874_),
    .A3(_06516_),
    .B1(_03834_),
    .B2(_00809_),
    .Y(_06517_));
 OR3x1_ASAP7_75t_R _13461_ (.A(_04583_),
    .B(_06515_),
    .C(_06517_),
    .Y(_06518_));
 AO221x1_ASAP7_75t_R _13462_ (.A1(_03815_),
    .A2(_04930_),
    .B1(_03829_),
    .B2(_03776_),
    .C(_00800_),
    .Y(_06519_));
 AO21x1_ASAP7_75t_R _13463_ (.A1(_04627_),
    .A2(_06519_),
    .B(_03786_),
    .Y(_06520_));
 AND4x2_ASAP7_75t_R _13464_ (.A(_00801_),
    .B(_03742_),
    .C(_03678_),
    .D(_04587_),
    .Y(_06521_));
 AO211x2_ASAP7_75t_R _13465_ (.A1(_00799_),
    .A2(_04583_),
    .B(_06521_),
    .C(_03879_),
    .Y(_06522_));
 AO32x2_ASAP7_75t_R _13466_ (.A1(_04839_),
    .A2(_06512_),
    .A3(_06518_),
    .B1(_06520_),
    .B2(_06522_),
    .Y(_06523_));
 AO211x2_ASAP7_75t_R _13467_ (.A1(_06481_),
    .A2(_06493_),
    .B(_06506_),
    .C(_06523_),
    .Y(_06524_));
 BUFx10_ASAP7_75t_R _13468_ (.A(_06524_),
    .Y(_10064_));
 INVx1_ASAP7_75t_R _13469_ (.A(_00855_),
    .Y(_06525_));
 NAND2x1_ASAP7_75t_R _13470_ (.A(_04017_),
    .B(_00857_),
    .Y(_06526_));
 OA211x2_ASAP7_75t_R _13471_ (.A1(_04269_),
    .A2(_06525_),
    .B(_06526_),
    .C(_03929_),
    .Y(_06527_));
 INVx1_ASAP7_75t_R _13472_ (.A(_00856_),
    .Y(_06528_));
 NAND2x1_ASAP7_75t_R _13473_ (.A(_04043_),
    .B(_00858_),
    .Y(_06529_));
 OA211x2_ASAP7_75t_R _13474_ (.A1(_04269_),
    .A2(_06528_),
    .B(_06529_),
    .C(_04256_),
    .Y(_06530_));
 OR3x1_ASAP7_75t_R _13475_ (.A(_04097_),
    .B(_06527_),
    .C(_06530_),
    .Y(_06531_));
 AND2x2_ASAP7_75t_R _13476_ (.A(_03956_),
    .B(_00849_),
    .Y(_06532_));
 AO21x1_ASAP7_75t_R _13477_ (.A1(_04040_),
    .A2(_00847_),
    .B(_06532_),
    .Y(_06533_));
 AO221x1_ASAP7_75t_R _13478_ (.A1(_04043_),
    .A2(_00850_),
    .B1(_04021_),
    .B2(_00848_),
    .C(_03949_),
    .Y(_06534_));
 OA211x2_ASAP7_75t_R _13479_ (.A1(_04307_),
    .A2(_06533_),
    .B(_06534_),
    .C(_03996_),
    .Y(_06535_));
 INVx1_ASAP7_75t_R _13480_ (.A(_06535_),
    .Y(_06536_));
 AND4x2_ASAP7_75t_R _13481_ (.A(_04296_),
    .B(_04051_),
    .C(_06531_),
    .D(_06536_),
    .Y(_06537_));
 AND2x2_ASAP7_75t_R _13482_ (.A(_04025_),
    .B(_00861_),
    .Y(_06538_));
 AO21x1_ASAP7_75t_R _13483_ (.A1(_03954_),
    .A2(_00859_),
    .B(_06538_),
    .Y(_06539_));
 AO222x2_ASAP7_75t_R _13484_ (.A1(_00862_),
    .A2(_03960_),
    .B1(_04266_),
    .B2(_00860_),
    .C1(_03976_),
    .C2(_06539_),
    .Y(_06540_));
 INVx1_ASAP7_75t_R _13485_ (.A(_00853_),
    .Y(_06541_));
 NAND2x1_ASAP7_75t_R _13486_ (.A(_03977_),
    .B(_00854_),
    .Y(_06542_));
 OA211x2_ASAP7_75t_R _13487_ (.A1(_04014_),
    .A2(_06541_),
    .B(_06542_),
    .C(_03973_),
    .Y(_06543_));
 INVx1_ASAP7_75t_R _13488_ (.A(_06543_),
    .Y(_06544_));
 AO221x1_ASAP7_75t_R _13489_ (.A1(_03949_),
    .A2(_00851_),
    .B1(_00852_),
    .B2(_03988_),
    .C(_03925_),
    .Y(_06545_));
 AO221x1_ASAP7_75t_R _13490_ (.A1(_04023_),
    .A2(_00851_),
    .B1(_06544_),
    .B2(_06545_),
    .C(_04279_),
    .Y(_06546_));
 OA21x2_ASAP7_75t_R _13491_ (.A1(_04414_),
    .A2(_06540_),
    .B(_06546_),
    .Y(_06547_));
 OR3x4_ASAP7_75t_R _13492_ (.A(_03418_),
    .B(_03429_),
    .C(_03419_),
    .Y(_06548_));
 NOR2x2_ASAP7_75t_R _13493_ (.A(_06547_),
    .B(_06548_),
    .Y(_06549_));
 AND2x2_ASAP7_75t_R _13494_ (.A(_03932_),
    .B(_00842_),
    .Y(_06550_));
 AO21x1_ASAP7_75t_R _13495_ (.A1(_04037_),
    .A2(_00841_),
    .B(_06550_),
    .Y(_06551_));
 AO221x1_ASAP7_75t_R _13496_ (.A1(_03985_),
    .A2(_00839_),
    .B1(_00840_),
    .B2(_03988_),
    .C(_04017_),
    .Y(_06552_));
 OA21x2_ASAP7_75t_R _13497_ (.A1(_04113_),
    .A2(_06551_),
    .B(_06552_),
    .Y(_06553_));
 AND2x2_ASAP7_75t_R _13498_ (.A(_03977_),
    .B(_00846_),
    .Y(_06554_));
 AO21x1_ASAP7_75t_R _13499_ (.A1(_03985_),
    .A2(_00845_),
    .B(_06554_),
    .Y(_06555_));
 AND3x1_ASAP7_75t_R _13500_ (.A(_03977_),
    .B(_03969_),
    .C(_00844_),
    .Y(_06556_));
 AO21x1_ASAP7_75t_R _13501_ (.A1(_00843_),
    .A2(_03548_),
    .B(_06556_),
    .Y(_06557_));
 AO221x1_ASAP7_75t_R _13502_ (.A1(_04269_),
    .A2(_06555_),
    .B1(_06557_),
    .B2(_03937_),
    .C(_03946_),
    .Y(_06558_));
 OA211x2_ASAP7_75t_R _13503_ (.A1(_04130_),
    .A2(_06553_),
    .B(_06558_),
    .C(_03920_),
    .Y(_06559_));
 AO22x1_ASAP7_75t_R _13504_ (.A1(_04037_),
    .A2(_00831_),
    .B1(_00832_),
    .B2(_03988_),
    .Y(_06560_));
 AND2x2_ASAP7_75t_R _13505_ (.A(_03931_),
    .B(_00834_),
    .Y(_06561_));
 AO21x1_ASAP7_75t_R _13506_ (.A1(_03928_),
    .A2(_00833_),
    .B(_06561_),
    .Y(_06562_));
 AO221x1_ASAP7_75t_R _13507_ (.A1(_03983_),
    .A2(_00831_),
    .B1(_04412_),
    .B2(_06562_),
    .C(_04406_),
    .Y(_06563_));
 AO21x1_ASAP7_75t_R _13508_ (.A1(_04073_),
    .A2(_06560_),
    .B(_06563_),
    .Y(_06564_));
 AND2x2_ASAP7_75t_R _13509_ (.A(_03977_),
    .B(_00838_),
    .Y(_06565_));
 AO21x1_ASAP7_75t_R _13510_ (.A1(_03949_),
    .A2(_00837_),
    .B(_06565_),
    .Y(_06566_));
 AND3x1_ASAP7_75t_R _13511_ (.A(_03977_),
    .B(_03378_),
    .C(_00836_),
    .Y(_06567_));
 AO21x1_ASAP7_75t_R _13512_ (.A1(_00835_),
    .A2(_03548_),
    .B(_06567_),
    .Y(_06568_));
 AO221x1_ASAP7_75t_R _13513_ (.A1(_03974_),
    .A2(_06566_),
    .B1(_06568_),
    .B2(_03937_),
    .C(_03946_),
    .Y(_06569_));
 AND3x4_ASAP7_75t_R _13514_ (.A(_04414_),
    .B(_06564_),
    .C(_06569_),
    .Y(_06570_));
 NOR3x2_ASAP7_75t_R _13515_ (.B(_06559_),
    .C(_06570_),
    .Y(_06571_),
    .A(_04429_));
 NOR3x2_ASAP7_75t_R _13516_ (.B(_06549_),
    .C(_06571_),
    .Y(_06572_),
    .A(_06537_));
 CKINVDCx12_ASAP7_75t_R _13517_ (.A(_06572_),
    .Y(net128));
 AND3x2_ASAP7_75t_R _13518_ (.A(net89),
    .B(net18),
    .C(_06285_),
    .Y(_10122_));
 AND2x2_ASAP7_75t_R _13519_ (.A(_04162_),
    .B(_10122_),
    .Y(_06573_));
 AOI21x1_ASAP7_75t_R _13520_ (.A1(_04065_),
    .A2(net128),
    .B(_06573_),
    .Y(_06574_));
 XNOR2x2_ASAP7_75t_R _13521_ (.A(_03537_),
    .B(_06574_),
    .Y(_10068_));
 INVx1_ASAP7_75t_R _13522_ (.A(_10068_),
    .Y(_10070_));
 AND3x1_ASAP7_75t_R _13523_ (.A(_06285_),
    .B(_03889_),
    .C(_03817_),
    .Y(_06575_));
 OR3x1_ASAP7_75t_R _13524_ (.A(_03482_),
    .B(_03840_),
    .C(_00844_),
    .Y(_06576_));
 OAI21x1_ASAP7_75t_R _13525_ (.A1(_00843_),
    .A2(_05640_),
    .B(_06576_),
    .Y(_06577_));
 AO21x1_ASAP7_75t_R _13526_ (.A1(_03662_),
    .A2(_03648_),
    .B(_03786_),
    .Y(_06578_));
 INVx1_ASAP7_75t_R _13527_ (.A(_00839_),
    .Y(_06579_));
 AND2x2_ASAP7_75t_R _13528_ (.A(_03853_),
    .B(_00842_),
    .Y(_06580_));
 AO21x1_ASAP7_75t_R _13529_ (.A1(_03840_),
    .A2(_00841_),
    .B(_06580_),
    .Y(_06581_));
 AND2x2_ASAP7_75t_R _13530_ (.A(_03853_),
    .B(_00846_),
    .Y(_06582_));
 AO21x1_ASAP7_75t_R _13531_ (.A1(_03840_),
    .A2(_00845_),
    .B(_06582_),
    .Y(_06583_));
 OAI22x1_ASAP7_75t_R _13532_ (.A1(_04948_),
    .A2(_06581_),
    .B1(_06583_),
    .B2(_03707_),
    .Y(_06584_));
 INVx1_ASAP7_75t_R _13533_ (.A(_00840_),
    .Y(_06585_));
 AND4x1_ASAP7_75t_R _13534_ (.A(_05331_),
    .B(_06585_),
    .C(_04591_),
    .D(_03776_),
    .Y(_06586_));
 OR3x1_ASAP7_75t_R _13535_ (.A(_04468_),
    .B(_06584_),
    .C(_06586_),
    .Y(_06587_));
 AOI221x1_ASAP7_75t_R _13536_ (.A1(_06575_),
    .A2(_06577_),
    .B1(_06578_),
    .B2(_06579_),
    .C(_06587_),
    .Y(_06588_));
 OA211x2_ASAP7_75t_R _13537_ (.A1(_03523_),
    .A2(_03880_),
    .B(_03728_),
    .C(_00836_),
    .Y(_06589_));
 AO21x1_ASAP7_75t_R _13538_ (.A1(_00835_),
    .A2(_03586_),
    .B(_06589_),
    .Y(_06590_));
 AO21x1_ASAP7_75t_R _13539_ (.A1(_03506_),
    .A2(_03508_),
    .B(_00838_),
    .Y(_06591_));
 AND2x2_ASAP7_75t_R _13540_ (.A(_00837_),
    .B(_03781_),
    .Y(_06592_));
 AO221x1_ASAP7_75t_R _13541_ (.A1(_03861_),
    .A2(_03888_),
    .B1(_06591_),
    .B2(_03882_),
    .C(_06592_),
    .Y(_06593_));
 OA21x2_ASAP7_75t_R _13542_ (.A1(_03795_),
    .A2(_06590_),
    .B(_06593_),
    .Y(_06594_));
 OA211x2_ASAP7_75t_R _13543_ (.A1(_03524_),
    .A2(_03880_),
    .B(_03728_),
    .C(_00832_),
    .Y(_06595_));
 AO21x1_ASAP7_75t_R _13544_ (.A1(_00831_),
    .A2(_03586_),
    .B(_06595_),
    .Y(_06596_));
 AND3x1_ASAP7_75t_R _13545_ (.A(_03843_),
    .B(_04460_),
    .C(_00834_),
    .Y(_06597_));
 AO21x1_ASAP7_75t_R _13546_ (.A1(_00833_),
    .A2(_04242_),
    .B(_06597_),
    .Y(_06598_));
 AND4x1_ASAP7_75t_R _13547_ (.A(_03742_),
    .B(_03557_),
    .C(_03783_),
    .D(_06598_),
    .Y(_06599_));
 AO21x1_ASAP7_75t_R _13548_ (.A1(_03889_),
    .A2(_06596_),
    .B(_06599_),
    .Y(_06600_));
 AO221x2_ASAP7_75t_R _13549_ (.A1(_05403_),
    .A2(_06594_),
    .B1(_06600_),
    .B2(_03773_),
    .C(_04452_),
    .Y(_06601_));
 AO32x1_ASAP7_75t_R _13550_ (.A1(_00857_),
    .A2(_03862_),
    .A3(_03831_),
    .B1(_04476_),
    .B2(_00861_),
    .Y(_06602_));
 AND3x1_ASAP7_75t_R _13551_ (.A(_03377_),
    .B(_04624_),
    .C(_00862_),
    .Y(_06603_));
 AND4x1_ASAP7_75t_R _13552_ (.A(_00858_),
    .B(_03777_),
    .C(_03774_),
    .D(_03838_),
    .Y(_06604_));
 AO21x1_ASAP7_75t_R _13553_ (.A1(_03872_),
    .A2(_06603_),
    .B(_06604_),
    .Y(_06605_));
 AND4x2_ASAP7_75t_R _13554_ (.A(_06285_),
    .B(_03678_),
    .C(_03868_),
    .D(_04587_),
    .Y(_06606_));
 OA21x2_ASAP7_75t_R _13555_ (.A1(_06602_),
    .A2(_06605_),
    .B(_06606_),
    .Y(_06607_));
 OA211x2_ASAP7_75t_R _13556_ (.A1(_03524_),
    .A2(_03880_),
    .B(_03728_),
    .C(_00856_),
    .Y(_06608_));
 AO21x1_ASAP7_75t_R _13557_ (.A1(_00855_),
    .A2(_03586_),
    .B(_06608_),
    .Y(_06609_));
 AND3x1_ASAP7_75t_R _13558_ (.A(_03375_),
    .B(_04435_),
    .C(_00860_),
    .Y(_06610_));
 AO21x1_ASAP7_75t_R _13559_ (.A1(_00859_),
    .A2(_04242_),
    .B(_06610_),
    .Y(_06611_));
 AND4x1_ASAP7_75t_R _13560_ (.A(_03742_),
    .B(_03678_),
    .C(_06097_),
    .D(_06611_),
    .Y(_06612_));
 AO21x1_ASAP7_75t_R _13561_ (.A1(_06094_),
    .A2(_06609_),
    .B(_06612_),
    .Y(_06613_));
 AND3x1_ASAP7_75t_R _13562_ (.A(_04596_),
    .B(_04436_),
    .C(_00852_),
    .Y(_06614_));
 AO21x1_ASAP7_75t_R _13563_ (.A1(_00851_),
    .A2(_04595_),
    .B(_06614_),
    .Y(_06615_));
 AND2x2_ASAP7_75t_R _13564_ (.A(_00853_),
    .B(_03781_),
    .Y(_06616_));
 AO221x1_ASAP7_75t_R _13565_ (.A1(_00854_),
    .A2(_03882_),
    .B1(_03888_),
    .B2(_03873_),
    .C(_06616_),
    .Y(_06617_));
 OA21x2_ASAP7_75t_R _13566_ (.A1(_03795_),
    .A2(_06615_),
    .B(_06617_),
    .Y(_06618_));
 OA22x2_ASAP7_75t_R _13567_ (.A1(_04436_),
    .A2(_00847_),
    .B1(_00848_),
    .B2(_04236_),
    .Y(_06619_));
 OA22x2_ASAP7_75t_R _13568_ (.A1(_03815_),
    .A2(_00847_),
    .B1(_06619_),
    .B2(_03816_),
    .Y(_06620_));
 AND2x2_ASAP7_75t_R _13569_ (.A(_00849_),
    .B(_04242_),
    .Y(_06621_));
 AO221x1_ASAP7_75t_R _13570_ (.A1(_00850_),
    .A2(_03882_),
    .B1(_04592_),
    .B2(_03873_),
    .C(_06621_),
    .Y(_06622_));
 AO31x2_ASAP7_75t_R _13571_ (.A1(_03773_),
    .A2(_06620_),
    .A3(_06622_),
    .B(_04499_),
    .Y(_06623_));
 AO221x2_ASAP7_75t_R _13572_ (.A1(_05510_),
    .A2(_06613_),
    .B1(_06618_),
    .B2(_05403_),
    .C(_06623_),
    .Y(_06624_));
 OAI22x1_ASAP7_75t_R _13573_ (.A1(_06588_),
    .A2(_06601_),
    .B1(_06607_),
    .B2(_06624_),
    .Y(_10067_));
 INVx6_ASAP7_75t_R _13574_ (.A(_10067_),
    .Y(_10069_));
 AO22x1_ASAP7_75t_R _13575_ (.A1(_04544_),
    .A2(_00888_),
    .B1(_04021_),
    .B2(_00886_),
    .Y(_06625_));
 AND2x2_ASAP7_75t_R _13576_ (.A(_03924_),
    .B(_00887_),
    .Y(_06626_));
 AO21x1_ASAP7_75t_R _13577_ (.A1(_04024_),
    .A2(_00885_),
    .B(_06626_),
    .Y(_06627_));
 AO221x1_ASAP7_75t_R _13578_ (.A1(_03983_),
    .A2(_00885_),
    .B1(_06627_),
    .B2(_04274_),
    .C(_03919_),
    .Y(_06628_));
 AO21x1_ASAP7_75t_R _13579_ (.A1(_04138_),
    .A2(_06625_),
    .B(_06628_),
    .Y(_06629_));
 AND2x2_ASAP7_75t_R _13580_ (.A(_03973_),
    .B(_00895_),
    .Y(_06630_));
 AO21x1_ASAP7_75t_R _13581_ (.A1(_04040_),
    .A2(_00893_),
    .B(_06630_),
    .Y(_06631_));
 AO21x1_ASAP7_75t_R _13582_ (.A1(_00896_),
    .A2(_03960_),
    .B(_03413_),
    .Y(_06632_));
 AO221x1_ASAP7_75t_R _13583_ (.A1(_00894_),
    .A2(_04266_),
    .B1(_06631_),
    .B2(_04125_),
    .C(_06632_),
    .Y(_06633_));
 AO21x1_ASAP7_75t_R _13584_ (.A1(_06629_),
    .A2(_06633_),
    .B(_04094_),
    .Y(_06634_));
 AND3x1_ASAP7_75t_R _13585_ (.A(_04666_),
    .B(_04269_),
    .C(_00892_),
    .Y(_06635_));
 AND2x2_ASAP7_75t_R _13586_ (.A(_03924_),
    .B(_00891_),
    .Y(_06636_));
 AO21x1_ASAP7_75t_R _13587_ (.A1(_04024_),
    .A2(_00889_),
    .B(_06636_),
    .Y(_06637_));
 AO32x1_ASAP7_75t_R _13588_ (.A1(_04040_),
    .A2(_00890_),
    .A3(_03989_),
    .B1(_06637_),
    .B2(_03998_),
    .Y(_06638_));
 OR3x1_ASAP7_75t_R _13589_ (.A(_04097_),
    .B(_06635_),
    .C(_06638_),
    .Y(_06639_));
 AND2x2_ASAP7_75t_R _13590_ (.A(_03924_),
    .B(_00883_),
    .Y(_06640_));
 AO21x1_ASAP7_75t_R _13591_ (.A1(_04024_),
    .A2(_00881_),
    .B(_06640_),
    .Y(_06641_));
 AO32x1_ASAP7_75t_R _13592_ (.A1(_04040_),
    .A2(_00882_),
    .A3(_03989_),
    .B1(_06641_),
    .B2(_03929_),
    .Y(_06642_));
 AO221x1_ASAP7_75t_R _13593_ (.A1(_04111_),
    .A2(_04315_),
    .B1(_00884_),
    .B2(_03961_),
    .C(_06642_),
    .Y(_06643_));
 AO21x1_ASAP7_75t_R _13594_ (.A1(_06639_),
    .A2(_06643_),
    .B(_04032_),
    .Y(_06644_));
 AOI21x1_ASAP7_75t_R _13595_ (.A1(_06634_),
    .A2(_06644_),
    .B(_03916_),
    .Y(_06645_));
 AND2x2_ASAP7_75t_R _13596_ (.A(_04536_),
    .B(_00868_),
    .Y(_06646_));
 AO21x1_ASAP7_75t_R _13597_ (.A1(_04028_),
    .A2(_00867_),
    .B(_06646_),
    .Y(_06647_));
 AO21x1_ASAP7_75t_R _13598_ (.A1(_04987_),
    .A2(_06647_),
    .B(_03981_),
    .Y(_06648_));
 AO22x1_ASAP7_75t_R _13599_ (.A1(_03998_),
    .A2(_00865_),
    .B1(_00866_),
    .B2(_03989_),
    .Y(_06649_));
 AO22x1_ASAP7_75t_R _13600_ (.A1(_03984_),
    .A2(_00865_),
    .B1(_06649_),
    .B2(_04276_),
    .Y(_06650_));
 AO21x1_ASAP7_75t_R _13601_ (.A1(_03972_),
    .A2(_06648_),
    .B(_06650_),
    .Y(_06651_));
 AND2x2_ASAP7_75t_R _13602_ (.A(_03932_),
    .B(_00872_),
    .Y(_06652_));
 AO21x1_ASAP7_75t_R _13603_ (.A1(_04037_),
    .A2(_00871_),
    .B(_06652_),
    .Y(_06653_));
 AND3x1_ASAP7_75t_R _13604_ (.A(_03932_),
    .B(_03378_),
    .C(_00870_),
    .Y(_06654_));
 AO21x1_ASAP7_75t_R _13605_ (.A1(_00869_),
    .A2(_03548_),
    .B(_06654_),
    .Y(_06655_));
 AO221x1_ASAP7_75t_R _13606_ (.A1(_04018_),
    .A2(_06653_),
    .B1(_06655_),
    .B2(_03937_),
    .C(_03946_),
    .Y(_06656_));
 AND2x2_ASAP7_75t_R _13607_ (.A(_04414_),
    .B(_06656_),
    .Y(_06657_));
 AND2x2_ASAP7_75t_R _13608_ (.A(_03932_),
    .B(_00880_),
    .Y(_06658_));
 AO21x1_ASAP7_75t_R _13609_ (.A1(_03929_),
    .A2(_00879_),
    .B(_06658_),
    .Y(_06659_));
 AND3x1_ASAP7_75t_R _13610_ (.A(_03941_),
    .B(_03378_),
    .C(_00878_),
    .Y(_06660_));
 AO21x1_ASAP7_75t_R _13611_ (.A1(_00877_),
    .A2(_04001_),
    .B(_06660_),
    .Y(_06661_));
 AO221x1_ASAP7_75t_R _13612_ (.A1(_04018_),
    .A2(_06659_),
    .B1(_06661_),
    .B2(_03937_),
    .C(_03946_),
    .Y(_06662_));
 AND2x2_ASAP7_75t_R _13613_ (.A(_03956_),
    .B(_00875_),
    .Y(_06663_));
 AO21x1_ASAP7_75t_R _13614_ (.A1(_04040_),
    .A2(_00873_),
    .B(_06663_),
    .Y(_06664_));
 AO21x1_ASAP7_75t_R _13615_ (.A1(_00874_),
    .A2(_03963_),
    .B(_03965_),
    .Y(_06665_));
 AO221x1_ASAP7_75t_R _13616_ (.A1(_00876_),
    .A2(_03961_),
    .B1(_06664_),
    .B2(_04281_),
    .C(_06665_),
    .Y(_06666_));
 AND3x1_ASAP7_75t_R _13617_ (.A(_04156_),
    .B(_06662_),
    .C(_06666_),
    .Y(_06667_));
 AOI211x1_ASAP7_75t_R _13618_ (.A1(_06651_),
    .A2(_06657_),
    .B(_04051_),
    .C(_06667_),
    .Y(_06668_));
 OAI21x1_ASAP7_75t_R _13619_ (.A1(_06645_),
    .A2(_06668_),
    .B(_03447_),
    .Y(_06669_));
 CKINVDCx11_ASAP7_75t_R _13620_ (.A(_06669_),
    .Y(net127));
 AND3x2_ASAP7_75t_R _13621_ (.A(net89),
    .B(net17),
    .C(_06285_),
    .Y(_10120_));
 AND2x2_ASAP7_75t_R _13622_ (.A(_04162_),
    .B(_10120_),
    .Y(_06670_));
 AOI21x1_ASAP7_75t_R _13623_ (.A1(_04065_),
    .A2(net127),
    .B(_06670_),
    .Y(_06671_));
 XNOR2x1_ASAP7_75t_R _13624_ (.B(_06671_),
    .Y(_10073_),
    .A(_03537_));
 INVx1_ASAP7_75t_R _13625_ (.A(_10073_),
    .Y(_10075_));
 AND3x1_ASAP7_75t_R _13626_ (.A(_04455_),
    .B(_04584_),
    .C(_00872_),
    .Y(_06672_));
 AO21x1_ASAP7_75t_R _13627_ (.A1(_00871_),
    .A2(_03891_),
    .B(_06672_),
    .Y(_06673_));
 OR2x2_ASAP7_75t_R _13628_ (.A(_04583_),
    .B(_06673_),
    .Y(_06674_));
 OA33x2_ASAP7_75t_R _13629_ (.A1(_00870_),
    .A2(_03586_),
    .A3(_03765_),
    .B1(_04344_),
    .B2(_03780_),
    .B3(_00869_),
    .Y(_06675_));
 AND3x1_ASAP7_75t_R _13630_ (.A(_03822_),
    .B(_04920_),
    .C(_06675_),
    .Y(_06676_));
 OR3x1_ASAP7_75t_R _13631_ (.A(_03482_),
    .B(_03840_),
    .C(_00866_),
    .Y(_06677_));
 AND3x1_ASAP7_75t_R _13632_ (.A(_03844_),
    .B(_03845_),
    .C(_00868_),
    .Y(_06678_));
 AO21x1_ASAP7_75t_R _13633_ (.A1(_00867_),
    .A2(_03796_),
    .B(_06678_),
    .Y(_06679_));
 AO21x1_ASAP7_75t_R _13634_ (.A1(_03901_),
    .A2(_06679_),
    .B(_04959_),
    .Y(_06680_));
 AO221x2_ASAP7_75t_R _13635_ (.A1(_06674_),
    .A2(_06676_),
    .B1(_06677_),
    .B2(_05846_),
    .C(_06680_),
    .Y(_06681_));
 AND3x1_ASAP7_75t_R _13636_ (.A(_00875_),
    .B(_03829_),
    .C(_03831_),
    .Y(_06682_));
 AO221x1_ASAP7_75t_R _13637_ (.A1(_00880_),
    .A2(_05230_),
    .B1(_04476_),
    .B2(_00879_),
    .C(_06682_),
    .Y(_06683_));
 AO21x1_ASAP7_75t_R _13638_ (.A1(_00876_),
    .A2(_05233_),
    .B(_03826_),
    .Y(_06684_));
 INVx1_ASAP7_75t_R _13639_ (.A(_00873_),
    .Y(_06685_));
 AND2x2_ASAP7_75t_R _13640_ (.A(_05332_),
    .B(_00878_),
    .Y(_06686_));
 AO21x1_ASAP7_75t_R _13641_ (.A1(_05331_),
    .A2(_00874_),
    .B(_06686_),
    .Y(_06687_));
 AOI22x1_ASAP7_75t_R _13642_ (.A1(_00877_),
    .A2(_04936_),
    .B1(_06687_),
    .B2(_03798_),
    .Y(_06688_));
 OA211x2_ASAP7_75t_R _13643_ (.A1(_04935_),
    .A2(_06688_),
    .B(_03776_),
    .C(_03777_),
    .Y(_06689_));
 OAI22x1_ASAP7_75t_R _13644_ (.A1(_06685_),
    .A2(_04934_),
    .B1(_06689_),
    .B2(_04165_),
    .Y(_06690_));
 OA211x2_ASAP7_75t_R _13645_ (.A1(_06683_),
    .A2(_06684_),
    .B(_03850_),
    .C(_06690_),
    .Y(_06691_));
 AO221x1_ASAP7_75t_R _13646_ (.A1(_00896_),
    .A2(_05230_),
    .B1(_05233_),
    .B2(_00892_),
    .C(_05218_),
    .Y(_06692_));
 AND3x1_ASAP7_75t_R _13647_ (.A(_00891_),
    .B(_03804_),
    .C(_03838_),
    .Y(_06693_));
 OA21x2_ASAP7_75t_R _13648_ (.A1(_03820_),
    .A2(_03817_),
    .B(_00895_),
    .Y(_06694_));
 OA21x2_ASAP7_75t_R _13649_ (.A1(_06693_),
    .A2(_06694_),
    .B(_04623_),
    .Y(_06695_));
 INVx1_ASAP7_75t_R _13650_ (.A(_00889_),
    .Y(_06696_));
 AND2x2_ASAP7_75t_R _13651_ (.A(_05332_),
    .B(_00894_),
    .Y(_06697_));
 AO21x1_ASAP7_75t_R _13652_ (.A1(_04937_),
    .A2(_00890_),
    .B(_06697_),
    .Y(_06698_));
 AOI22x1_ASAP7_75t_R _13653_ (.A1(_00893_),
    .A2(_04936_),
    .B1(_06698_),
    .B2(_03798_),
    .Y(_06699_));
 OA211x2_ASAP7_75t_R _13654_ (.A1(_04935_),
    .A2(_06699_),
    .B(_03776_),
    .C(_03777_),
    .Y(_06700_));
 OAI22x1_ASAP7_75t_R _13655_ (.A1(_06696_),
    .A2(_04934_),
    .B1(_06700_),
    .B2(_03786_),
    .Y(_06701_));
 OA211x2_ASAP7_75t_R _13656_ (.A1(_06692_),
    .A2(_06695_),
    .B(_03850_),
    .C(_06701_),
    .Y(_06702_));
 OA211x2_ASAP7_75t_R _13657_ (.A1(_03524_),
    .A2(_03880_),
    .B(_03728_),
    .C(_00886_),
    .Y(_06703_));
 AO21x1_ASAP7_75t_R _13658_ (.A1(_00885_),
    .A2(_03586_),
    .B(_06703_),
    .Y(_06704_));
 AND2x2_ASAP7_75t_R _13659_ (.A(_00887_),
    .B(_04236_),
    .Y(_06705_));
 AO221x1_ASAP7_75t_R _13660_ (.A1(_00888_),
    .A2(_03882_),
    .B1(_04592_),
    .B2(_03829_),
    .C(_06705_),
    .Y(_06706_));
 OA21x2_ASAP7_75t_R _13661_ (.A1(_03795_),
    .A2(_06704_),
    .B(_06706_),
    .Y(_06707_));
 INVx1_ASAP7_75t_R _13662_ (.A(_00883_),
    .Y(_06708_));
 INVx1_ASAP7_75t_R _13663_ (.A(_00882_),
    .Y(_06709_));
 NAND2x1_ASAP7_75t_R _13664_ (.A(_03816_),
    .B(_00884_),
    .Y(_06710_));
 OA211x2_ASAP7_75t_R _13665_ (.A1(_03816_),
    .A2(_06709_),
    .B(_06710_),
    .C(_05215_),
    .Y(_06711_));
 AOI21x1_ASAP7_75t_R _13666_ (.A1(_06708_),
    .A2(_04442_),
    .B(_06711_),
    .Y(_06712_));
 OA22x2_ASAP7_75t_R _13667_ (.A1(_00881_),
    .A2(_04344_),
    .B1(_06712_),
    .B2(_03482_),
    .Y(_06713_));
 AO221x2_ASAP7_75t_R _13668_ (.A1(_05403_),
    .A2(_06707_),
    .B1(_06713_),
    .B2(_03773_),
    .C(_03809_),
    .Y(_06714_));
 OAI22x1_ASAP7_75t_R _13669_ (.A1(_06681_),
    .A2(_06691_),
    .B1(_06702_),
    .B2(_06714_),
    .Y(_10072_));
 INVx5_ASAP7_75t_R _13670_ (.A(_10072_),
    .Y(_10074_));
 AND2x2_ASAP7_75t_R _13671_ (.A(_03940_),
    .B(_00913_),
    .Y(_06715_));
 AO21x1_ASAP7_75t_R _13672_ (.A1(_03985_),
    .A2(_00912_),
    .B(_06715_),
    .Y(_06716_));
 AND3x1_ASAP7_75t_R _13673_ (.A(_03940_),
    .B(_03969_),
    .C(_00911_),
    .Y(_06717_));
 AO21x1_ASAP7_75t_R _13674_ (.A1(_00910_),
    .A2(_03548_),
    .B(_06717_),
    .Y(_06718_));
 AO221x1_ASAP7_75t_R _13675_ (.A1(_04075_),
    .A2(_06716_),
    .B1(_06718_),
    .B2(_03937_),
    .C(_03449_),
    .Y(_06719_));
 AND2x2_ASAP7_75t_R _13676_ (.A(_03924_),
    .B(_00908_),
    .Y(_06720_));
 AO21x1_ASAP7_75t_R _13677_ (.A1(_03953_),
    .A2(_00906_),
    .B(_06720_),
    .Y(_06721_));
 AO21x1_ASAP7_75t_R _13678_ (.A1(_00907_),
    .A2(_03963_),
    .B(_03412_),
    .Y(_06722_));
 AO221x1_ASAP7_75t_R _13679_ (.A1(_00909_),
    .A2(_03960_),
    .B1(_06721_),
    .B2(_03929_),
    .C(_06722_),
    .Y(_06723_));
 AND3x1_ASAP7_75t_R _13680_ (.A(_04279_),
    .B(_06719_),
    .C(_06723_),
    .Y(_06724_));
 AO22x1_ASAP7_75t_R _13681_ (.A1(_03928_),
    .A2(_00898_),
    .B1(_00899_),
    .B2(_03988_),
    .Y(_06725_));
 AND2x2_ASAP7_75t_R _13682_ (.A(_03931_),
    .B(_00901_),
    .Y(_06726_));
 AO21x1_ASAP7_75t_R _13683_ (.A1(_03928_),
    .A2(_00900_),
    .B(_06726_),
    .Y(_06727_));
 AO21x1_ASAP7_75t_R _13684_ (.A1(_03973_),
    .A2(_06727_),
    .B(_03412_),
    .Y(_06728_));
 AND2x2_ASAP7_75t_R _13685_ (.A(_03482_),
    .B(_00898_),
    .Y(_06729_));
 AO221x1_ASAP7_75t_R _13686_ (.A1(_03954_),
    .A2(_06725_),
    .B1(_06728_),
    .B2(_03379_),
    .C(_06729_),
    .Y(_06730_));
 AND2x2_ASAP7_75t_R _13687_ (.A(_03940_),
    .B(_00905_),
    .Y(_06731_));
 AO21x1_ASAP7_75t_R _13688_ (.A1(_03985_),
    .A2(_00904_),
    .B(_06731_),
    .Y(_06732_));
 AND3x1_ASAP7_75t_R _13689_ (.A(_03940_),
    .B(_03969_),
    .C(_00903_),
    .Y(_06733_));
 AO21x1_ASAP7_75t_R _13690_ (.A1(_00902_),
    .A2(_03548_),
    .B(_06733_),
    .Y(_06734_));
 AO221x1_ASAP7_75t_R _13691_ (.A1(_04075_),
    .A2(_06732_),
    .B1(_06734_),
    .B2(_03937_),
    .C(_03449_),
    .Y(_06735_));
 AND3x1_ASAP7_75t_R _13692_ (.A(_04097_),
    .B(_06730_),
    .C(_06735_),
    .Y(_06736_));
 OA21x2_ASAP7_75t_R _13693_ (.A1(_06724_),
    .A2(_06736_),
    .B(_03916_),
    .Y(_06737_));
 AND2x2_ASAP7_75t_R _13694_ (.A(_04403_),
    .B(_00921_),
    .Y(_06738_));
 AO21x1_ASAP7_75t_R _13695_ (.A1(_04274_),
    .A2(_00920_),
    .B(_06738_),
    .Y(_06739_));
 AO21x1_ASAP7_75t_R _13696_ (.A1(_04529_),
    .A2(_06739_),
    .B(_04297_),
    .Y(_06740_));
 AND3x1_ASAP7_75t_R _13697_ (.A(_03941_),
    .B(_03970_),
    .C(_00919_),
    .Y(_06741_));
 AO21x1_ASAP7_75t_R _13698_ (.A1(_00918_),
    .A2(_04001_),
    .B(_06741_),
    .Y(_06742_));
 AND2x2_ASAP7_75t_R _13699_ (.A(_04004_),
    .B(_06742_),
    .Y(_06743_));
 AND2x2_ASAP7_75t_R _13700_ (.A(_03940_),
    .B(_00929_),
    .Y(_06744_));
 AO21x1_ASAP7_75t_R _13701_ (.A1(_03985_),
    .A2(_00928_),
    .B(_06744_),
    .Y(_06745_));
 AO21x1_ASAP7_75t_R _13702_ (.A1(_03957_),
    .A2(_06745_),
    .B(_03420_),
    .Y(_06746_));
 AND3x1_ASAP7_75t_R _13703_ (.A(_03940_),
    .B(_03969_),
    .C(_00927_),
    .Y(_06747_));
 AO21x1_ASAP7_75t_R _13704_ (.A1(_00926_),
    .A2(_03548_),
    .B(_06747_),
    .Y(_06748_));
 AND2x2_ASAP7_75t_R _13705_ (.A(_03936_),
    .B(_06748_),
    .Y(_06749_));
 OA21x2_ASAP7_75t_R _13706_ (.A1(_06746_),
    .A2(_06749_),
    .B(_04051_),
    .Y(_06750_));
 AO221x1_ASAP7_75t_R _13707_ (.A1(_03924_),
    .A2(_00925_),
    .B1(_04020_),
    .B2(_00923_),
    .C(_03995_),
    .Y(_06751_));
 AO221x1_ASAP7_75t_R _13708_ (.A1(_03924_),
    .A2(_00917_),
    .B1(_04020_),
    .B2(_00915_),
    .C(_03919_),
    .Y(_06752_));
 AND3x1_ASAP7_75t_R _13709_ (.A(_04033_),
    .B(_06751_),
    .C(_06752_),
    .Y(_06753_));
 AND2x2_ASAP7_75t_R _13710_ (.A(_03923_),
    .B(_00924_),
    .Y(_06754_));
 AO21x1_ASAP7_75t_R _13711_ (.A1(_03953_),
    .A2(_00922_),
    .B(_06754_),
    .Y(_06755_));
 AND2x2_ASAP7_75t_R _13712_ (.A(_03923_),
    .B(_00916_),
    .Y(_06756_));
 AO221x1_ASAP7_75t_R _13713_ (.A1(_03442_),
    .A2(_03969_),
    .B1(_00914_),
    .B2(_03953_),
    .C(_06756_),
    .Y(_06757_));
 OA211x2_ASAP7_75t_R _13714_ (.A1(_03996_),
    .A2(_06755_),
    .B(_06757_),
    .C(_03949_),
    .Y(_06758_));
 OR3x1_ASAP7_75t_R _13715_ (.A(_03966_),
    .B(_06753_),
    .C(_06758_),
    .Y(_06759_));
 OA211x2_ASAP7_75t_R _13716_ (.A1(_06740_),
    .A2(_06743_),
    .B(_06750_),
    .C(_06759_),
    .Y(_06760_));
 OR3x4_ASAP7_75t_R _13717_ (.A(_04055_),
    .B(_06737_),
    .C(_06760_),
    .Y(_06761_));
 INVx11_ASAP7_75t_R _13718_ (.A(_06761_),
    .Y(net126));
 AND3x2_ASAP7_75t_R _13719_ (.A(_03382_),
    .B(net16),
    .C(_06285_),
    .Y(_10118_));
 AND2x2_ASAP7_75t_R _13720_ (.A(_04162_),
    .B(_10118_),
    .Y(_06762_));
 AOI21x1_ASAP7_75t_R _13721_ (.A1(_04065_),
    .A2(net126),
    .B(_06762_),
    .Y(_06763_));
 XNOR2x2_ASAP7_75t_R _13722_ (.A(_03537_),
    .B(_06763_),
    .Y(_10078_));
 INVx1_ASAP7_75t_R _13723_ (.A(_10078_),
    .Y(_10080_));
 AND3x1_ASAP7_75t_R _13724_ (.A(_04916_),
    .B(_03853_),
    .C(_00921_),
    .Y(_06764_));
 AO21x1_ASAP7_75t_R _13725_ (.A1(_00920_),
    .A2(_03891_),
    .B(_06764_),
    .Y(_06765_));
 AND3x1_ASAP7_75t_R _13726_ (.A(_03375_),
    .B(_04435_),
    .C(_00917_),
    .Y(_06766_));
 AO21x1_ASAP7_75t_R _13727_ (.A1(_00916_),
    .A2(_03781_),
    .B(_06766_),
    .Y(_06767_));
 AND2x2_ASAP7_75t_R _13728_ (.A(_00914_),
    .B(_03612_),
    .Y(_06768_));
 AO221x1_ASAP7_75t_R _13729_ (.A1(_03639_),
    .A2(_03816_),
    .B1(_00915_),
    .B2(_03881_),
    .C(_06768_),
    .Y(_06769_));
 OA211x2_ASAP7_75t_R _13730_ (.A1(_04454_),
    .A2(_06767_),
    .B(_06769_),
    .C(_03772_),
    .Y(_06770_));
 AND3x1_ASAP7_75t_R _13731_ (.A(_03843_),
    .B(_03762_),
    .C(_00919_),
    .Y(_06771_));
 AO21x1_ASAP7_75t_R _13732_ (.A1(_00918_),
    .A2(_03761_),
    .B(_06771_),
    .Y(_06772_));
 AO21x1_ASAP7_75t_R _13733_ (.A1(_03721_),
    .A2(_06772_),
    .B(_03723_),
    .Y(_06773_));
 AOI211x1_ASAP7_75t_R _13734_ (.A1(_04440_),
    .A2(_06765_),
    .B(_06770_),
    .C(_06773_),
    .Y(_06774_));
 AND2x2_ASAP7_75t_R _13735_ (.A(_03685_),
    .B(_00927_),
    .Y(_06775_));
 AO21x1_ASAP7_75t_R _13736_ (.A1(_03744_),
    .A2(_00923_),
    .B(_06775_),
    .Y(_06776_));
 AO22x1_ASAP7_75t_R _13737_ (.A1(_00926_),
    .A2(_04456_),
    .B1(_06776_),
    .B2(_03624_),
    .Y(_06777_));
 NAND2x1_ASAP7_75t_R _13738_ (.A(_03663_),
    .B(_06777_),
    .Y(_06778_));
 AO21x1_ASAP7_75t_R _13739_ (.A1(_03824_),
    .A2(_06778_),
    .B(_04163_),
    .Y(_06779_));
 NAND2x1_ASAP7_75t_R _13740_ (.A(_00922_),
    .B(_03750_),
    .Y(_06780_));
 AND3x1_ASAP7_75t_R _13741_ (.A(_00924_),
    .B(_03646_),
    .C(_03830_),
    .Y(_06781_));
 AOI221x1_ASAP7_75t_R _13742_ (.A1(_00929_),
    .A2(_04198_),
    .B1(_04199_),
    .B2(_00928_),
    .C(_06781_),
    .Y(_06782_));
 AOI21x1_ASAP7_75t_R _13743_ (.A1(_00925_),
    .A2(_03834_),
    .B(_04454_),
    .Y(_06783_));
 AO221x2_ASAP7_75t_R _13744_ (.A1(_06779_),
    .A2(_06780_),
    .B1(_06782_),
    .B2(_06783_),
    .C(_03740_),
    .Y(_06784_));
 AND3x1_ASAP7_75t_R _13745_ (.A(_03623_),
    .B(_03624_),
    .C(_00905_),
    .Y(_06785_));
 AO21x1_ASAP7_75t_R _13746_ (.A1(_00904_),
    .A2(_03890_),
    .B(_06785_),
    .Y(_06786_));
 AO21x2_ASAP7_75t_R _13747_ (.A1(_03506_),
    .A2(_03508_),
    .B(_04952_),
    .Y(_06787_));
 OA222x2_ASAP7_75t_R _13748_ (.A1(_00902_),
    .A2(_04492_),
    .B1(_03658_),
    .B2(_06786_),
    .C1(_06787_),
    .C2(_00903_),
    .Y(_06788_));
 AND3x1_ASAP7_75t_R _13749_ (.A(_03843_),
    .B(_04460_),
    .C(_00901_),
    .Y(_06789_));
 AO21x1_ASAP7_75t_R _13750_ (.A1(_00900_),
    .A2(_04236_),
    .B(_06789_),
    .Y(_06790_));
 AND2x2_ASAP7_75t_R _13751_ (.A(_03900_),
    .B(_06790_),
    .Y(_06791_));
 OR3x1_ASAP7_75t_R _13752_ (.A(_04811_),
    .B(_03629_),
    .C(_00899_),
    .Y(_06792_));
 AO21x1_ASAP7_75t_R _13753_ (.A1(_05846_),
    .A2(_06792_),
    .B(_04959_),
    .Y(_06793_));
 AOI211x1_ASAP7_75t_R _13754_ (.A1(_03791_),
    .A2(_06788_),
    .B(_06791_),
    .C(_06793_),
    .Y(_06794_));
 AND2x2_ASAP7_75t_R _13755_ (.A(_03685_),
    .B(_00911_),
    .Y(_06795_));
 AO21x1_ASAP7_75t_R _13756_ (.A1(_03744_),
    .A2(_00907_),
    .B(_06795_),
    .Y(_06796_));
 AO22x1_ASAP7_75t_R _13757_ (.A1(_00910_),
    .A2(_04456_),
    .B1(_06796_),
    .B2(_03624_),
    .Y(_06797_));
 NAND2x1_ASAP7_75t_R _13758_ (.A(_03663_),
    .B(_06797_),
    .Y(_06798_));
 AO21x1_ASAP7_75t_R _13759_ (.A1(_04454_),
    .A2(_06798_),
    .B(_04163_),
    .Y(_06799_));
 NAND2x1_ASAP7_75t_R _13760_ (.A(_00906_),
    .B(_03750_),
    .Y(_06800_));
 AND3x1_ASAP7_75t_R _13761_ (.A(_00908_),
    .B(_03646_),
    .C(_03830_),
    .Y(_06801_));
 AOI221x1_ASAP7_75t_R _13762_ (.A1(_00913_),
    .A2(_04198_),
    .B1(_04199_),
    .B2(_00912_),
    .C(_06801_),
    .Y(_06802_));
 AOI21x1_ASAP7_75t_R _13763_ (.A1(_00909_),
    .A2(_03834_),
    .B(_04454_),
    .Y(_06803_));
 AO221x2_ASAP7_75t_R _13764_ (.A1(_06799_),
    .A2(_06800_),
    .B1(_06802_),
    .B2(_06803_),
    .C(_04468_),
    .Y(_06804_));
 AO22x1_ASAP7_75t_R _13765_ (.A1(_06774_),
    .A2(_06784_),
    .B1(_06794_),
    .B2(_06804_),
    .Y(_06805_));
 BUFx6f_ASAP7_75t_R _13766_ (.A(_06805_),
    .Y(_10077_));
 INVx5_ASAP7_75t_R _13767_ (.A(_10077_),
    .Y(_10079_));
 AOI211x1_ASAP7_75t_R _13768_ (.A1(_03497_),
    .A2(_03503_),
    .B(_03600_),
    .C(_03572_),
    .Y(_06806_));
 AND2x2_ASAP7_75t_R _13769_ (.A(_03797_),
    .B(net3),
    .Y(_06807_));
 AO32x1_ASAP7_75t_R _13770_ (.A1(_04050_),
    .A2(_06806_),
    .A3(_03547_),
    .B1(_06807_),
    .B2(_03503_),
    .Y(_06808_));
 BUFx2_ASAP7_75t_R _13771_ (.A(_06808_),
    .Y(_10116_));
 BUFx4f_ASAP7_75t_R _13772_ (.A(_03396_),
    .Y(_06809_));
 AND3x1_ASAP7_75t_R _13773_ (.A(_06809_),
    .B(_03843_),
    .C(_00962_),
    .Y(_06810_));
 AO21x1_ASAP7_75t_R _13774_ (.A1(_00946_),
    .A2(_03384_),
    .B(_06810_),
    .Y(_06811_));
 AND3x1_ASAP7_75t_R _13775_ (.A(_03396_),
    .B(_03623_),
    .C(_00954_),
    .Y(_06812_));
 AO221x1_ASAP7_75t_R _13776_ (.A1(_03442_),
    .A2(_03639_),
    .B1(_00938_),
    .B2(_03384_),
    .C(_06812_),
    .Y(_06813_));
 BUFx4f_ASAP7_75t_R _13777_ (.A(_03426_),
    .Y(_06814_));
 OA211x2_ASAP7_75t_R _13778_ (.A1(_03995_),
    .A2(_06811_),
    .B(_06813_),
    .C(_06814_),
    .Y(_06815_));
 AND3x1_ASAP7_75t_R _13779_ (.A(_06809_),
    .B(_03843_),
    .C(_00960_),
    .Y(_06816_));
 AO21x1_ASAP7_75t_R _13780_ (.A1(_00944_),
    .A2(_03384_),
    .B(_06816_),
    .Y(_06817_));
 AND3x1_ASAP7_75t_R _13781_ (.A(_03396_),
    .B(_03623_),
    .C(_00952_),
    .Y(_06818_));
 AO221x1_ASAP7_75t_R _13782_ (.A1(_03442_),
    .A2(_03715_),
    .B1(_00936_),
    .B2(_03384_),
    .C(_06818_),
    .Y(_06819_));
 OA211x2_ASAP7_75t_R _13783_ (.A1(_03995_),
    .A2(_06817_),
    .B(_06819_),
    .C(_03953_),
    .Y(_06820_));
 OR3x1_ASAP7_75t_R _13784_ (.A(_03931_),
    .B(_04296_),
    .C(_05417_),
    .Y(_06821_));
 OR3x1_ASAP7_75t_R _13785_ (.A(_03928_),
    .B(_04296_),
    .C(_05417_),
    .Y(_06822_));
 AND2x2_ASAP7_75t_R _13786_ (.A(_03426_),
    .B(_00963_),
    .Y(_06823_));
 AO21x1_ASAP7_75t_R _13787_ (.A1(_03952_),
    .A2(_00961_),
    .B(_06823_),
    .Y(_06824_));
 AO21x1_ASAP7_75t_R _13788_ (.A1(_03386_),
    .A2(_00945_),
    .B(_06809_),
    .Y(_06825_));
 AO22x1_ASAP7_75t_R _13789_ (.A1(_06814_),
    .A2(_00947_),
    .B1(_06825_),
    .B2(_04916_),
    .Y(_06826_));
 OA211x2_ASAP7_75t_R _13790_ (.A1(_03384_),
    .A2(_06824_),
    .B(_06826_),
    .C(_03918_),
    .Y(_06827_));
 AND2x2_ASAP7_75t_R _13791_ (.A(_03922_),
    .B(_00955_),
    .Y(_06828_));
 AO21x1_ASAP7_75t_R _13792_ (.A1(_03952_),
    .A2(_00953_),
    .B(_06828_),
    .Y(_06829_));
 AO21x1_ASAP7_75t_R _13793_ (.A1(_03386_),
    .A2(_00937_),
    .B(_06809_),
    .Y(_06830_));
 AO22x1_ASAP7_75t_R _13794_ (.A1(_06814_),
    .A2(_00939_),
    .B1(_06830_),
    .B2(_04916_),
    .Y(_06831_));
 OA211x2_ASAP7_75t_R _13795_ (.A1(_03916_),
    .A2(_06829_),
    .B(_06831_),
    .C(_03995_),
    .Y(_06832_));
 OA33x2_ASAP7_75t_R _13796_ (.A1(_06815_),
    .A2(_06820_),
    .A3(_06821_),
    .B1(_06822_),
    .B2(_06827_),
    .B3(_06832_),
    .Y(_06833_));
 OR3x1_ASAP7_75t_R _13797_ (.A(_03411_),
    .B(_03429_),
    .C(_03415_),
    .Y(_06834_));
 AND2x2_ASAP7_75t_R _13798_ (.A(_03922_),
    .B(_00950_),
    .Y(_06835_));
 AO21x1_ASAP7_75t_R _13799_ (.A1(_03952_),
    .A2(_00948_),
    .B(_06835_),
    .Y(_06836_));
 AO221x1_ASAP7_75t_R _13800_ (.A1(_06814_),
    .A2(_00951_),
    .B1(_04020_),
    .B2(_00949_),
    .C(_03423_),
    .Y(_06837_));
 OA21x2_ASAP7_75t_R _13801_ (.A1(_03931_),
    .A2(_06836_),
    .B(_06837_),
    .Y(_06838_));
 BUFx4f_ASAP7_75t_R _13802_ (.A(net12),
    .Y(_06839_));
 BUFx4f_ASAP7_75t_R _13803_ (.A(_06839_),
    .Y(_06840_));
 AND2x2_ASAP7_75t_R _13804_ (.A(_06840_),
    .B(_00935_),
    .Y(_06841_));
 AO21x1_ASAP7_75t_R _13805_ (.A1(_03423_),
    .A2(_00934_),
    .B(_06841_),
    .Y(_06842_));
 AO221x1_ASAP7_75t_R _13806_ (.A1(_05417_),
    .A2(_00932_),
    .B1(_04412_),
    .B2(_06842_),
    .C(_04406_),
    .Y(_06843_));
 AND4x1_ASAP7_75t_R _13807_ (.A(_06840_),
    .B(_03952_),
    .C(_03715_),
    .D(_00933_),
    .Y(_06844_));
 AO221x1_ASAP7_75t_R _13808_ (.A1(_06809_),
    .A2(_03797_),
    .B1(_00932_),
    .B2(_03405_),
    .C(_06844_),
    .Y(_06845_));
 OAI22x1_ASAP7_75t_R _13809_ (.A1(_06834_),
    .A2(_06838_),
    .B1(_06843_),
    .B2(_06845_),
    .Y(_06846_));
 AOI22x1_ASAP7_75t_R _13810_ (.A1(_06814_),
    .A2(_00959_),
    .B1(_04020_),
    .B2(_00957_),
    .Y(_06847_));
 INVx1_ASAP7_75t_R _13811_ (.A(_00956_),
    .Y(_06848_));
 NAND2x1_ASAP7_75t_R _13812_ (.A(_03426_),
    .B(_00958_),
    .Y(_06849_));
 BUFx4f_ASAP7_75t_R _13813_ (.A(_03421_),
    .Y(_06850_));
 OA211x2_ASAP7_75t_R _13814_ (.A1(_03922_),
    .A2(_06848_),
    .B(_06849_),
    .C(_06850_),
    .Y(_06851_));
 AO21x1_ASAP7_75t_R _13815_ (.A1(_03931_),
    .A2(_06847_),
    .B(_06851_),
    .Y(_06852_));
 NAND2x1_ASAP7_75t_R _13816_ (.A(_03423_),
    .B(_00940_),
    .Y(_06853_));
 INVx1_ASAP7_75t_R _13817_ (.A(_00941_),
    .Y(_06854_));
 OR3x1_ASAP7_75t_R _13818_ (.A(_06850_),
    .B(_04811_),
    .C(_06854_),
    .Y(_06855_));
 AO21x1_ASAP7_75t_R _13819_ (.A1(_06853_),
    .A2(_06855_),
    .B(_03923_),
    .Y(_06856_));
 AND2x2_ASAP7_75t_R _13820_ (.A(_06840_),
    .B(_00943_),
    .Y(_06857_));
 AO21x1_ASAP7_75t_R _13821_ (.A1(_03423_),
    .A2(_00942_),
    .B(_06857_),
    .Y(_06858_));
 AOI221x1_ASAP7_75t_R _13822_ (.A1(_05417_),
    .A2(_00940_),
    .B1(_06858_),
    .B2(_03923_),
    .C(_04050_),
    .Y(_06859_));
 AO32x1_ASAP7_75t_R _13823_ (.A1(_06809_),
    .A2(_04053_),
    .A3(_06852_),
    .B1(_06856_),
    .B2(_06859_),
    .Y(_06860_));
 AND3x1_ASAP7_75t_R _13824_ (.A(_04296_),
    .B(_03442_),
    .C(_04053_),
    .Y(_06861_));
 AOI22x1_ASAP7_75t_R _13825_ (.A1(_03995_),
    .A2(_06846_),
    .B1(_06860_),
    .B2(_06861_),
    .Y(_06862_));
 AO21x2_ASAP7_75t_R _13826_ (.A1(_06833_),
    .A2(_06862_),
    .B(_04054_),
    .Y(_06863_));
 CKINVDCx12_ASAP7_75t_R _13827_ (.A(_06863_),
    .Y(net125));
 OR2x2_ASAP7_75t_R _13828_ (.A(_04059_),
    .B(_10116_),
    .Y(_06864_));
 OA21x2_ASAP7_75t_R _13829_ (.A1(_03915_),
    .A2(net125),
    .B(_06864_),
    .Y(_06865_));
 BUFx6f_ASAP7_75t_R _13830_ (.A(_06865_),
    .Y(_06866_));
 BUFx4f_ASAP7_75t_R _13831_ (.A(_06866_),
    .Y(_06867_));
 XNOR2x1_ASAP7_75t_R _13832_ (.B(_06867_),
    .Y(_10083_),
    .A(_03913_));
 INVx1_ASAP7_75t_R _13833_ (.A(_10083_),
    .Y(_10085_));
 AND3x1_ASAP7_75t_R _13834_ (.A(_03815_),
    .B(_04930_),
    .C(_00955_),
    .Y(_06868_));
 AO21x1_ASAP7_75t_R _13835_ (.A1(_00954_),
    .A2(_04929_),
    .B(_06868_),
    .Y(_06869_));
 AND3x1_ASAP7_75t_R _13836_ (.A(_03844_),
    .B(_03845_),
    .C(_00953_),
    .Y(_06870_));
 AO21x1_ASAP7_75t_R _13837_ (.A1(_00952_),
    .A2(_03796_),
    .B(_06870_),
    .Y(_06871_));
 AO21x1_ASAP7_75t_R _13838_ (.A1(_03721_),
    .A2(_06871_),
    .B(_04499_),
    .Y(_06872_));
 AND3x1_ASAP7_75t_R _13839_ (.A(_03376_),
    .B(_05215_),
    .C(_00949_),
    .Y(_06873_));
 AO21x1_ASAP7_75t_R _13840_ (.A1(_00948_),
    .A2(_04434_),
    .B(_06873_),
    .Y(_06874_));
 AND2x2_ASAP7_75t_R _13841_ (.A(_00950_),
    .B(_03781_),
    .Y(_06875_));
 AO221x1_ASAP7_75t_R _13842_ (.A1(_00951_),
    .A2(_03882_),
    .B1(_03888_),
    .B2(_03873_),
    .C(_06875_),
    .Y(_06876_));
 OA211x2_ASAP7_75t_R _13843_ (.A1(_03783_),
    .A2(_06874_),
    .B(_06876_),
    .C(_03773_),
    .Y(_06877_));
 AOI211x1_ASAP7_75t_R _13844_ (.A1(_04440_),
    .A2(_06869_),
    .B(_06872_),
    .C(_06877_),
    .Y(_06878_));
 AND2x2_ASAP7_75t_R _13845_ (.A(_04938_),
    .B(_00961_),
    .Y(_06879_));
 AO21x1_ASAP7_75t_R _13846_ (.A1(_04937_),
    .A2(_00957_),
    .B(_06879_),
    .Y(_06880_));
 AO22x1_ASAP7_75t_R _13847_ (.A1(_00960_),
    .A2(_05221_),
    .B1(_06880_),
    .B2(_05215_),
    .Y(_06881_));
 NAND2x1_ASAP7_75t_R _13848_ (.A(_03377_),
    .B(_06881_),
    .Y(_06882_));
 AO21x1_ASAP7_75t_R _13849_ (.A1(_05218_),
    .A2(_06882_),
    .B(_04806_),
    .Y(_06883_));
 NAND2x1_ASAP7_75t_R _13850_ (.A(_00956_),
    .B(_03811_),
    .Y(_06884_));
 AND3x1_ASAP7_75t_R _13851_ (.A(_00958_),
    .B(_03777_),
    .C(_03831_),
    .Y(_06885_));
 AOI221x1_ASAP7_75t_R _13852_ (.A1(_00963_),
    .A2(_05230_),
    .B1(_04476_),
    .B2(_00962_),
    .C(_06885_),
    .Y(_06886_));
 AOI21x1_ASAP7_75t_R _13853_ (.A1(_00959_),
    .A2(_05233_),
    .B(_03826_),
    .Y(_06887_));
 AO221x2_ASAP7_75t_R _13854_ (.A1(_06883_),
    .A2(_06884_),
    .B1(_06886_),
    .B2(_06887_),
    .C(_05235_),
    .Y(_06888_));
 AND3x1_ASAP7_75t_R _13855_ (.A(_04455_),
    .B(_04597_),
    .C(_00939_),
    .Y(_06889_));
 AO21x1_ASAP7_75t_R _13856_ (.A1(_00938_),
    .A2(_03782_),
    .B(_06889_),
    .Y(_06890_));
 OR3x1_ASAP7_75t_R _13857_ (.A(_00937_),
    .B(_03878_),
    .C(_03765_),
    .Y(_06891_));
 OR3x1_ASAP7_75t_R _13858_ (.A(_00936_),
    .B(_03780_),
    .C(_04344_),
    .Y(_06892_));
 OA211x2_ASAP7_75t_R _13859_ (.A1(_04583_),
    .A2(_06890_),
    .B(_06891_),
    .C(_06892_),
    .Y(_06893_));
 AND3x1_ASAP7_75t_R _13860_ (.A(_03844_),
    .B(_03845_),
    .C(_00935_),
    .Y(_06894_));
 AO21x1_ASAP7_75t_R _13861_ (.A1(_00934_),
    .A2(_03796_),
    .B(_06894_),
    .Y(_06895_));
 AO21x1_ASAP7_75t_R _13862_ (.A1(_03901_),
    .A2(_06895_),
    .B(_04959_),
    .Y(_06896_));
 OA21x2_ASAP7_75t_R _13863_ (.A1(_00933_),
    .A2(_04623_),
    .B(_05846_),
    .Y(_06897_));
 AOI211x1_ASAP7_75t_R _13864_ (.A1(_03792_),
    .A2(_06893_),
    .B(_06896_),
    .C(_06897_),
    .Y(_06898_));
 AND2x2_ASAP7_75t_R _13865_ (.A(_04938_),
    .B(_00945_),
    .Y(_06899_));
 AO21x1_ASAP7_75t_R _13866_ (.A1(_04937_),
    .A2(_00941_),
    .B(_06899_),
    .Y(_06900_));
 AO22x1_ASAP7_75t_R _13867_ (.A1(_00944_),
    .A2(_04800_),
    .B1(_06900_),
    .B2(_05215_),
    .Y(_06901_));
 NAND2x1_ASAP7_75t_R _13868_ (.A(_03377_),
    .B(_06901_),
    .Y(_06902_));
 AO21x1_ASAP7_75t_R _13869_ (.A1(_05218_),
    .A2(_06902_),
    .B(_04806_),
    .Y(_06903_));
 NAND2x1_ASAP7_75t_R _13870_ (.A(_00940_),
    .B(_03811_),
    .Y(_06904_));
 AND3x1_ASAP7_75t_R _13871_ (.A(_00942_),
    .B(_03777_),
    .C(_03831_),
    .Y(_06905_));
 AOI221x1_ASAP7_75t_R _13872_ (.A1(_00947_),
    .A2(_05230_),
    .B1(_04476_),
    .B2(_00946_),
    .C(_06905_),
    .Y(_06906_));
 AOI21x1_ASAP7_75t_R _13873_ (.A1(_00943_),
    .A2(_05233_),
    .B(_03826_),
    .Y(_06907_));
 AO221x2_ASAP7_75t_R _13874_ (.A1(_06903_),
    .A2(_06904_),
    .B1(_06906_),
    .B2(_06907_),
    .C(_05235_),
    .Y(_06908_));
 AOI22x1_ASAP7_75t_R _13875_ (.A1(_06878_),
    .A2(_06888_),
    .B1(_06898_),
    .B2(_06908_),
    .Y(_10084_));
 AO32x2_ASAP7_75t_R _13876_ (.A1(_04053_),
    .A2(net2),
    .A3(_03501_),
    .B1(_04172_),
    .B2(_03919_),
    .Y(_06909_));
 NAND2x2_ASAP7_75t_R _13877_ (.A(_04171_),
    .B(_06909_),
    .Y(_06910_));
 NAND2x1_ASAP7_75t_R _13878_ (.A(net2),
    .B(_04166_),
    .Y(_06911_));
 OA21x2_ASAP7_75t_R _13879_ (.A1(_03413_),
    .A2(net64),
    .B(_06911_),
    .Y(_06912_));
 OR4x2_ASAP7_75t_R _13880_ (.A(_03482_),
    .B(_05227_),
    .C(_03542_),
    .D(_06912_),
    .Y(_06913_));
 NAND2x1_ASAP7_75t_R _13881_ (.A(_06910_),
    .B(_06913_),
    .Y(_10114_));
 AO221x1_ASAP7_75t_R _13882_ (.A1(_03423_),
    .A2(_00993_),
    .B1(_00994_),
    .B2(_03988_),
    .C(_06814_),
    .Y(_06914_));
 INVx1_ASAP7_75t_R _13883_ (.A(_00996_),
    .Y(_06915_));
 NOR2x1_ASAP7_75t_R _13884_ (.A(_06840_),
    .B(_00995_),
    .Y(_06916_));
 AO21x1_ASAP7_75t_R _13885_ (.A1(_06840_),
    .A2(_06915_),
    .B(_06916_),
    .Y(_06917_));
 NAND2x1_ASAP7_75t_R _13886_ (.A(_06814_),
    .B(_06917_),
    .Y(_06918_));
 AO21x1_ASAP7_75t_R _13887_ (.A1(_06914_),
    .A2(_06918_),
    .B(_03995_),
    .Y(_06919_));
 AO221x1_ASAP7_75t_R _13888_ (.A1(_06850_),
    .A2(_00985_),
    .B1(_00986_),
    .B2(_03987_),
    .C(_03922_),
    .Y(_06920_));
 AND2x2_ASAP7_75t_R _13889_ (.A(_06839_),
    .B(_00988_),
    .Y(_06921_));
 AO21x1_ASAP7_75t_R _13890_ (.A1(_03422_),
    .A2(_00987_),
    .B(_06921_),
    .Y(_06922_));
 OR2x2_ASAP7_75t_R _13891_ (.A(_03952_),
    .B(_06922_),
    .Y(_06923_));
 AO221x1_ASAP7_75t_R _13892_ (.A1(_03481_),
    .A2(_00985_),
    .B1(_06920_),
    .B2(_06923_),
    .C(_03919_),
    .Y(_06924_));
 AO22x1_ASAP7_75t_R _13893_ (.A1(_03426_),
    .A2(_00992_),
    .B1(_04020_),
    .B2(_00990_),
    .Y(_06925_));
 AND2x2_ASAP7_75t_R _13894_ (.A(_03432_),
    .B(_00984_),
    .Y(_06926_));
 AO221x1_ASAP7_75t_R _13895_ (.A1(_03442_),
    .A2(_03549_),
    .B1(_00982_),
    .B2(_04019_),
    .C(_06926_),
    .Y(_06927_));
 OA211x2_ASAP7_75t_R _13896_ (.A1(_03444_),
    .A2(_06925_),
    .B(_06927_),
    .C(_06840_),
    .Y(_06928_));
 AND2x2_ASAP7_75t_R _13897_ (.A(_03392_),
    .B(_00991_),
    .Y(_06929_));
 AO21x1_ASAP7_75t_R _13898_ (.A1(_03386_),
    .A2(_00989_),
    .B(_06929_),
    .Y(_06930_));
 AND2x2_ASAP7_75t_R _13899_ (.A(_03432_),
    .B(_00983_),
    .Y(_06931_));
 AO221x1_ASAP7_75t_R _13900_ (.A1(_03442_),
    .A2(_03549_),
    .B1(_00981_),
    .B2(_03386_),
    .C(_06931_),
    .Y(_06932_));
 OA211x2_ASAP7_75t_R _13901_ (.A1(_03444_),
    .A2(_06930_),
    .B(_06932_),
    .C(_03423_),
    .Y(_06933_));
 OA21x2_ASAP7_75t_R _13902_ (.A1(_06928_),
    .A2(_06933_),
    .B(_04296_),
    .Y(_06934_));
 AO31x2_ASAP7_75t_R _13903_ (.A1(_03412_),
    .A2(_06919_),
    .A3(_06924_),
    .B(_06934_),
    .Y(_06935_));
 AND2x2_ASAP7_75t_R _13904_ (.A(_03922_),
    .B(_00971_),
    .Y(_06936_));
 AO21x1_ASAP7_75t_R _13905_ (.A1(_03952_),
    .A2(_00969_),
    .B(_06936_),
    .Y(_06937_));
 AO221x1_ASAP7_75t_R _13906_ (.A1(_06814_),
    .A2(_00972_),
    .B1(_04020_),
    .B2(_00970_),
    .C(_03423_),
    .Y(_06938_));
 OA21x2_ASAP7_75t_R _13907_ (.A1(_03931_),
    .A2(_06937_),
    .B(_06938_),
    .Y(_06939_));
 OA21x2_ASAP7_75t_R _13908_ (.A1(_03449_),
    .A2(_06939_),
    .B(_03995_),
    .Y(_06940_));
 AND2x2_ASAP7_75t_R _13909_ (.A(_03400_),
    .B(_00968_),
    .Y(_06941_));
 AO21x1_ASAP7_75t_R _13910_ (.A1(_06850_),
    .A2(_00967_),
    .B(_06941_),
    .Y(_06942_));
 AO21x1_ASAP7_75t_R _13911_ (.A1(_06814_),
    .A2(_06942_),
    .B(_03412_),
    .Y(_06943_));
 AND2x2_ASAP7_75t_R _13912_ (.A(_03815_),
    .B(_06943_),
    .Y(_06944_));
 AO22x1_ASAP7_75t_R _13913_ (.A1(_03423_),
    .A2(_00965_),
    .B1(_00966_),
    .B2(_03988_),
    .Y(_06945_));
 AO22x1_ASAP7_75t_R _13914_ (.A1(_04935_),
    .A2(_00965_),
    .B1(_06945_),
    .B2(_03953_),
    .Y(_06946_));
 OA21x2_ASAP7_75t_R _13915_ (.A1(_06944_),
    .A2(_06946_),
    .B(_03916_),
    .Y(_06947_));
 AND2x2_ASAP7_75t_R _13916_ (.A(_03392_),
    .B(_00975_),
    .Y(_06948_));
 AO21x1_ASAP7_75t_R _13917_ (.A1(_03386_),
    .A2(_00973_),
    .B(_06948_),
    .Y(_06949_));
 AO221x1_ASAP7_75t_R _13918_ (.A1(_03426_),
    .A2(_00976_),
    .B1(_04020_),
    .B2(_00974_),
    .C(_06850_),
    .Y(_06950_));
 OA21x2_ASAP7_75t_R _13919_ (.A1(_03931_),
    .A2(_06949_),
    .B(_06950_),
    .Y(_06951_));
 OR2x2_ASAP7_75t_R _13920_ (.A(_03412_),
    .B(_06951_),
    .Y(_06952_));
 AND2x2_ASAP7_75t_R _13921_ (.A(_03400_),
    .B(_00980_),
    .Y(_06953_));
 AO21x1_ASAP7_75t_R _13922_ (.A1(_06850_),
    .A2(_00979_),
    .B(_06953_),
    .Y(_06954_));
 AO21x1_ASAP7_75t_R _13923_ (.A1(_06814_),
    .A2(_06954_),
    .B(_03449_),
    .Y(_06955_));
 AND3x1_ASAP7_75t_R _13924_ (.A(_06840_),
    .B(_03639_),
    .C(_00978_),
    .Y(_06956_));
 OA21x2_ASAP7_75t_R _13925_ (.A1(_06850_),
    .A2(_03480_),
    .B(_00977_),
    .Y(_06957_));
 OA21x2_ASAP7_75t_R _13926_ (.A1(_06956_),
    .A2(_06957_),
    .B(_03936_),
    .Y(_06958_));
 OA211x2_ASAP7_75t_R _13927_ (.A1(_06955_),
    .A2(_06958_),
    .B(_03916_),
    .C(_03919_),
    .Y(_06959_));
 AO21x1_ASAP7_75t_R _13928_ (.A1(_06952_),
    .A2(_06959_),
    .B(_04054_),
    .Y(_06960_));
 AO221x2_ASAP7_75t_R _13929_ (.A1(_04050_),
    .A2(_06935_),
    .B1(_06940_),
    .B2(_06947_),
    .C(_06960_),
    .Y(_06961_));
 CKINVDCx10_ASAP7_75t_R _13930_ (.A(_06961_),
    .Y(net124));
 AND3x2_ASAP7_75t_R _13931_ (.A(_03915_),
    .B(_06910_),
    .C(_06913_),
    .Y(_06962_));
 AOI21x1_ASAP7_75t_R _13932_ (.A1(_04059_),
    .A2(_06961_),
    .B(_06962_),
    .Y(_06963_));
 BUFx6f_ASAP7_75t_R _13933_ (.A(_06963_),
    .Y(_06964_));
 BUFx4f_ASAP7_75t_R _13934_ (.A(_06964_),
    .Y(_06965_));
 BUFx6f_ASAP7_75t_R _13935_ (.A(_06965_),
    .Y(_06966_));
 XNOR2x1_ASAP7_75t_R _13936_ (.B(_06966_),
    .Y(_10088_),
    .A(_03913_));
 INVx1_ASAP7_75t_R _13937_ (.A(_10088_),
    .Y(_10090_));
 AND2x2_ASAP7_75t_R _13938_ (.A(_05332_),
    .B(_00994_),
    .Y(_06967_));
 AO21x1_ASAP7_75t_R _13939_ (.A1(_05331_),
    .A2(_00990_),
    .B(_06967_),
    .Y(_06968_));
 AO22x1_ASAP7_75t_R _13940_ (.A1(_00993_),
    .A2(_04936_),
    .B1(_06968_),
    .B2(_03798_),
    .Y(_06969_));
 NAND2x1_ASAP7_75t_R _13941_ (.A(_03969_),
    .B(_06969_),
    .Y(_06970_));
 AO21x1_ASAP7_75t_R _13942_ (.A1(_03826_),
    .A2(_06970_),
    .B(_03786_),
    .Y(_06971_));
 NAND2x1_ASAP7_75t_R _13943_ (.A(_00989_),
    .B(_03811_),
    .Y(_06972_));
 AND2x2_ASAP7_75t_R _13944_ (.A(_00995_),
    .B(_03796_),
    .Y(_06973_));
 AND2x2_ASAP7_75t_R _13945_ (.A(_00991_),
    .B(_03714_),
    .Y(_06974_));
 AO32x1_ASAP7_75t_R _13946_ (.A1(_03837_),
    .A2(_03838_),
    .A3(_06974_),
    .B1(_03834_),
    .B2(_00992_),
    .Y(_06975_));
 AOI221x1_ASAP7_75t_R _13947_ (.A1(_00996_),
    .A2(_05230_),
    .B1(_06973_),
    .B2(_03872_),
    .C(_06975_),
    .Y(_06976_));
 AO221x1_ASAP7_75t_R _13948_ (.A1(_06971_),
    .A2(_06972_),
    .B1(_06976_),
    .B2(_03852_),
    .C(_05235_),
    .Y(_06977_));
 AND3x1_ASAP7_75t_R _13949_ (.A(_03377_),
    .B(_04624_),
    .C(_00988_),
    .Y(_06978_));
 AO21x1_ASAP7_75t_R _13950_ (.A1(_00987_),
    .A2(_04929_),
    .B(_06978_),
    .Y(_06979_));
 NAND2x1_ASAP7_75t_R _13951_ (.A(_03852_),
    .B(_06979_),
    .Y(_06980_));
 NAND2x1_ASAP7_75t_R _13952_ (.A(_00986_),
    .B(_03814_),
    .Y(_06981_));
 NAND2x1_ASAP7_75t_R _13953_ (.A(_00985_),
    .B(_03587_),
    .Y(_06982_));
 AO21x1_ASAP7_75t_R _13954_ (.A1(_06981_),
    .A2(_06982_),
    .B(_03852_),
    .Y(_06983_));
 NAND2x1_ASAP7_75t_R _13955_ (.A(_03822_),
    .B(_04920_),
    .Y(_06984_));
 AO21x1_ASAP7_75t_R _13956_ (.A1(_06980_),
    .A2(_06983_),
    .B(_06984_),
    .Y(_06985_));
 INVx1_ASAP7_75t_R _13957_ (.A(_00981_),
    .Y(_06986_));
 INVx1_ASAP7_75t_R _13958_ (.A(_00983_),
    .Y(_06987_));
 INVx1_ASAP7_75t_R _13959_ (.A(_00982_),
    .Y(_06988_));
 NAND2x1_ASAP7_75t_R _13960_ (.A(_03816_),
    .B(_00984_),
    .Y(_06989_));
 OA211x2_ASAP7_75t_R _13961_ (.A1(_03816_),
    .A2(_06988_),
    .B(_06989_),
    .C(_04436_),
    .Y(_06990_));
 AO21x1_ASAP7_75t_R _13962_ (.A1(_06987_),
    .A2(_04442_),
    .B(_06990_),
    .Y(_06991_));
 AO32x1_ASAP7_75t_R _13963_ (.A1(_06986_),
    .A2(_04623_),
    .A3(_03889_),
    .B1(_06991_),
    .B2(_03969_),
    .Y(_06992_));
 OA21x2_ASAP7_75t_R _13964_ (.A1(_05713_),
    .A2(_06992_),
    .B(_03907_),
    .Y(_06993_));
 AND2x2_ASAP7_75t_R _13965_ (.A(_05332_),
    .B(_00978_),
    .Y(_06994_));
 AO21x1_ASAP7_75t_R _13966_ (.A1(_04937_),
    .A2(_00974_),
    .B(_06994_),
    .Y(_06995_));
 AO22x1_ASAP7_75t_R _13967_ (.A1(_00977_),
    .A2(_04936_),
    .B1(_06995_),
    .B2(_03845_),
    .Y(_06996_));
 NAND2x1_ASAP7_75t_R _13968_ (.A(_04053_),
    .B(_06996_),
    .Y(_06997_));
 AO21x1_ASAP7_75t_R _13969_ (.A1(_03826_),
    .A2(_06997_),
    .B(_03786_),
    .Y(_06998_));
 NAND2x1_ASAP7_75t_R _13970_ (.A(_00973_),
    .B(_03811_),
    .Y(_06999_));
 AND3x1_ASAP7_75t_R _13971_ (.A(_00975_),
    .B(_03837_),
    .C(_03831_),
    .Y(_07000_));
 AOI221x1_ASAP7_75t_R _13972_ (.A1(_00980_),
    .A2(_05230_),
    .B1(_04476_),
    .B2(_00979_),
    .C(_07000_),
    .Y(_07001_));
 AOI21x1_ASAP7_75t_R _13973_ (.A1(_00976_),
    .A2(_05233_),
    .B(_04792_),
    .Y(_07002_));
 AO221x1_ASAP7_75t_R _13974_ (.A1(_06998_),
    .A2(_06999_),
    .B1(_07001_),
    .B2(_07002_),
    .C(_05235_),
    .Y(_07003_));
 AND3x1_ASAP7_75t_R _13975_ (.A(_03797_),
    .B(_04930_),
    .C(_00972_),
    .Y(_07004_));
 AO21x1_ASAP7_75t_R _13976_ (.A1(_00971_),
    .A2(_04929_),
    .B(_07004_),
    .Y(_07005_));
 OA222x2_ASAP7_75t_R _13977_ (.A1(_00969_),
    .A2(_04492_),
    .B1(_04583_),
    .B2(_07005_),
    .C1(_06787_),
    .C2(_00970_),
    .Y(_07006_));
 AND3x1_ASAP7_75t_R _13978_ (.A(_03797_),
    .B(_03798_),
    .C(_00968_),
    .Y(_07007_));
 AO21x1_ASAP7_75t_R _13979_ (.A1(_00967_),
    .A2(_04929_),
    .B(_07007_),
    .Y(_07008_));
 OR3x1_ASAP7_75t_R _13980_ (.A(_04935_),
    .B(_03840_),
    .C(_00966_),
    .Y(_07009_));
 AO221x1_ASAP7_75t_R _13981_ (.A1(_03901_),
    .A2(_07008_),
    .B1(_07009_),
    .B2(_05846_),
    .C(_04959_),
    .Y(_07010_));
 AOI21x1_ASAP7_75t_R _13982_ (.A1(_03792_),
    .A2(_07006_),
    .B(_07010_),
    .Y(_07011_));
 AO32x2_ASAP7_75t_R _13983_ (.A1(_06977_),
    .A2(_06985_),
    .A3(_06993_),
    .B1(_07003_),
    .B2(_07011_),
    .Y(_07012_));
 BUFx6f_ASAP7_75t_R _13984_ (.A(_07012_),
    .Y(_10087_));
 INVx1_ASAP7_75t_R _13985_ (.A(_10087_),
    .Y(_10089_));
 NAND3x1_ASAP7_75t_R _13986_ (.A(_03497_),
    .B(_03502_),
    .C(_03557_),
    .Y(_07013_));
 AND3x1_ASAP7_75t_R _13987_ (.A(_03493_),
    .B(_03494_),
    .C(_03563_),
    .Y(_07014_));
 AND4x1_ASAP7_75t_R _13988_ (.A(_03486_),
    .B(_03489_),
    .C(_03754_),
    .D(_07014_),
    .Y(_07015_));
 AO22x1_ASAP7_75t_R _13989_ (.A1(_03375_),
    .A2(net30),
    .B1(_03474_),
    .B2(_03540_),
    .Y(_07016_));
 AO21x1_ASAP7_75t_R _13990_ (.A1(_04406_),
    .A2(_04172_),
    .B(_03501_),
    .Y(_07017_));
 OAI21x1_ASAP7_75t_R _13991_ (.A1(_07015_),
    .A2(_07016_),
    .B(_07017_),
    .Y(_07018_));
 AND2x2_ASAP7_75t_R _13992_ (.A(_03449_),
    .B(_03547_),
    .Y(_07019_));
 NAND2x2_ASAP7_75t_R _13993_ (.A(_03394_),
    .B(net30),
    .Y(_07020_));
 AND2x2_ASAP7_75t_R _13994_ (.A(_04166_),
    .B(_07020_),
    .Y(_07021_));
 OR4x1_ASAP7_75t_R _13995_ (.A(_03599_),
    .B(_03572_),
    .C(_07019_),
    .D(_07021_),
    .Y(_07022_));
 OA22x2_ASAP7_75t_R _13996_ (.A1(_07013_),
    .A2(_07018_),
    .B1(_07022_),
    .B2(_03542_),
    .Y(_07023_));
 BUFx4f_ASAP7_75t_R _13997_ (.A(_07023_),
    .Y(_07024_));
 INVx1_ASAP7_75t_R _13998_ (.A(_07024_),
    .Y(_10108_));
 AND2x2_ASAP7_75t_R _13999_ (.A(_03432_),
    .B(_01013_),
    .Y(_07025_));
 AOI21x1_ASAP7_75t_R _14000_ (.A1(_03386_),
    .A2(_01011_),
    .B(_07025_),
    .Y(_07026_));
 INVx1_ASAP7_75t_R _14001_ (.A(_01010_),
    .Y(_07027_));
 NAND2x1_ASAP7_75t_R _14002_ (.A(_03388_),
    .B(_01012_),
    .Y(_07028_));
 OA211x2_ASAP7_75t_R _14003_ (.A1(_03392_),
    .A2(_07027_),
    .B(_07028_),
    .C(_03407_),
    .Y(_07029_));
 AO21x1_ASAP7_75t_R _14004_ (.A1(_06840_),
    .A2(_07026_),
    .B(_07029_),
    .Y(_07030_));
 NAND2x1_ASAP7_75t_R _14005_ (.A(_06850_),
    .B(_01006_),
    .Y(_07031_));
 INVx1_ASAP7_75t_R _14006_ (.A(_01007_),
    .Y(_07032_));
 OR3x1_ASAP7_75t_R _14007_ (.A(_03407_),
    .B(_03628_),
    .C(_07032_),
    .Y(_07033_));
 AO21x1_ASAP7_75t_R _14008_ (.A1(_07031_),
    .A2(_07033_),
    .B(_03922_),
    .Y(_07034_));
 AND2x2_ASAP7_75t_R _14009_ (.A(_06839_),
    .B(_01009_),
    .Y(_07035_));
 AO21x1_ASAP7_75t_R _14010_ (.A1(_03422_),
    .A2(_01008_),
    .B(_07035_),
    .Y(_07036_));
 AOI221x1_ASAP7_75t_R _14011_ (.A1(_03480_),
    .A2(_01006_),
    .B1(_04412_),
    .B2(_07036_),
    .C(_04406_),
    .Y(_07037_));
 AO221x1_ASAP7_75t_R _14012_ (.A1(_04406_),
    .A2(_07030_),
    .B1(_07034_),
    .B2(_07037_),
    .C(_04050_),
    .Y(_07038_));
 AO221x1_ASAP7_75t_R _14013_ (.A1(_06850_),
    .A2(_01026_),
    .B1(_01027_),
    .B2(_03987_),
    .C(_03922_),
    .Y(_07039_));
 AND2x2_ASAP7_75t_R _14014_ (.A(_06839_),
    .B(_01029_),
    .Y(_07040_));
 AO21x1_ASAP7_75t_R _14015_ (.A1(_03422_),
    .A2(_01028_),
    .B(_07040_),
    .Y(_07041_));
 AND3x1_ASAP7_75t_R _14016_ (.A(_03412_),
    .B(_03396_),
    .C(_03549_),
    .Y(_07042_));
 OA21x2_ASAP7_75t_R _14017_ (.A1(_03952_),
    .A2(_07041_),
    .B(_07042_),
    .Y(_07043_));
 AND2x2_ASAP7_75t_R _14018_ (.A(_03432_),
    .B(_01024_),
    .Y(_07044_));
 AO21x1_ASAP7_75t_R _14019_ (.A1(_03386_),
    .A2(_01022_),
    .B(_07044_),
    .Y(_07045_));
 AO221x1_ASAP7_75t_R _14020_ (.A1(_03392_),
    .A2(_01025_),
    .B1(_04019_),
    .B2(_01023_),
    .C(_03407_),
    .Y(_07046_));
 OA211x2_ASAP7_75t_R _14021_ (.A1(_06840_),
    .A2(_07045_),
    .B(_07046_),
    .C(_03418_),
    .Y(_07047_));
 AOI221x1_ASAP7_75t_R _14022_ (.A1(_07039_),
    .A2(_07043_),
    .B1(_07047_),
    .B2(_04050_),
    .C(_03995_),
    .Y(_07048_));
 NAND2x1_ASAP7_75t_R _14023_ (.A(_03422_),
    .B(_00998_),
    .Y(_07049_));
 INVx1_ASAP7_75t_R _14024_ (.A(_00999_),
    .Y(_07050_));
 OR3x1_ASAP7_75t_R _14025_ (.A(_03407_),
    .B(_03628_),
    .C(_07050_),
    .Y(_07051_));
 AO21x1_ASAP7_75t_R _14026_ (.A1(_07049_),
    .A2(_07051_),
    .B(_03922_),
    .Y(_07052_));
 AND2x2_ASAP7_75t_R _14027_ (.A(_06839_),
    .B(_01001_),
    .Y(_07053_));
 AO21x1_ASAP7_75t_R _14028_ (.A1(_03422_),
    .A2(_01000_),
    .B(_07053_),
    .Y(_07054_));
 AOI221x1_ASAP7_75t_R _14029_ (.A1(_03480_),
    .A2(_00998_),
    .B1(_04412_),
    .B2(_07054_),
    .C(_04406_),
    .Y(_07055_));
 AND2x2_ASAP7_75t_R _14030_ (.A(_03432_),
    .B(_01004_),
    .Y(_07056_));
 AO21x1_ASAP7_75t_R _14031_ (.A1(_03386_),
    .A2(_01002_),
    .B(_07056_),
    .Y(_07057_));
 AND3x1_ASAP7_75t_R _14032_ (.A(_06839_),
    .B(_03432_),
    .C(_01005_),
    .Y(_07058_));
 OR3x1_ASAP7_75t_R _14033_ (.A(_03418_),
    .B(_03628_),
    .C(_07058_),
    .Y(_07059_));
 AOI221x1_ASAP7_75t_R _14034_ (.A1(_01003_),
    .A2(_03963_),
    .B1(_07057_),
    .B2(_06850_),
    .C(_07059_),
    .Y(_07060_));
 AO221x1_ASAP7_75t_R _14035_ (.A1(_06809_),
    .A2(_04596_),
    .B1(_07052_),
    .B2(_07055_),
    .C(_07060_),
    .Y(_07061_));
 AND2x2_ASAP7_75t_R _14036_ (.A(_06839_),
    .B(_01021_),
    .Y(_07062_));
 AO21x1_ASAP7_75t_R _14037_ (.A1(_03422_),
    .A2(_01020_),
    .B(_07062_),
    .Y(_07063_));
 AO21x1_ASAP7_75t_R _14038_ (.A1(_03422_),
    .A2(_01018_),
    .B(_03426_),
    .Y(_07064_));
 AND3x1_ASAP7_75t_R _14039_ (.A(_03400_),
    .B(_03549_),
    .C(_01019_),
    .Y(_07065_));
 OAI22x1_ASAP7_75t_R _14040_ (.A1(_03952_),
    .A2(_07063_),
    .B1(_07064_),
    .B2(_07065_),
    .Y(_07066_));
 AOI221x1_ASAP7_75t_R _14041_ (.A1(_03426_),
    .A2(_01017_),
    .B1(_04019_),
    .B2(_01015_),
    .C(_03422_),
    .Y(_07067_));
 INVx1_ASAP7_75t_R _14042_ (.A(_01014_),
    .Y(_07068_));
 NAND2x1_ASAP7_75t_R _14043_ (.A(_03388_),
    .B(_01016_),
    .Y(_07069_));
 OA211x2_ASAP7_75t_R _14044_ (.A1(_03392_),
    .A2(_07068_),
    .B(_07069_),
    .C(_03421_),
    .Y(_07070_));
 OR3x1_ASAP7_75t_R _14045_ (.A(_06834_),
    .B(_07067_),
    .C(_07070_),
    .Y(_07071_));
 AND3x1_ASAP7_75t_R _14046_ (.A(_03413_),
    .B(_03623_),
    .C(_03445_),
    .Y(_07072_));
 OA211x2_ASAP7_75t_R _14047_ (.A1(_06548_),
    .A2(_07066_),
    .B(_07071_),
    .C(_07072_),
    .Y(_07073_));
 AOI22x1_ASAP7_75t_R _14048_ (.A1(_07038_),
    .A2(_07048_),
    .B1(_07061_),
    .B2(_07073_),
    .Y(_07074_));
 BUFx12_ASAP7_75t_R _14049_ (.A(_07074_),
    .Y(_07075_));
 CKINVDCx10_ASAP7_75t_R _14050_ (.A(_07075_),
    .Y(net121));
 AND2x2_ASAP7_75t_R _14051_ (.A(_04058_),
    .B(_07074_),
    .Y(_07076_));
 AOI21x1_ASAP7_75t_R _14052_ (.A1(_03915_),
    .A2(_07024_),
    .B(_07076_),
    .Y(_07077_));
 BUFx4f_ASAP7_75t_R _14053_ (.A(_07077_),
    .Y(_07078_));
 BUFx4f_ASAP7_75t_R _14054_ (.A(_07078_),
    .Y(_07079_));
 BUFx6f_ASAP7_75t_R _14055_ (.A(_07079_),
    .Y(_07080_));
 BUFx6f_ASAP7_75t_R _14056_ (.A(_07080_),
    .Y(_07081_));
 XNOR2x1_ASAP7_75t_R _14057_ (.B(_07081_),
    .Y(_10093_),
    .A(_03913_));
 INVx1_ASAP7_75t_R _14058_ (.A(_10093_),
    .Y(_10095_));
 INVx1_ASAP7_75t_R _14059_ (.A(_01006_),
    .Y(_07082_));
 NAND2x1_ASAP7_75t_R _14060_ (.A(_01011_),
    .B(_05640_),
    .Y(_07083_));
 OA21x2_ASAP7_75t_R _14061_ (.A1(_07027_),
    .A2(_05640_),
    .B(_07083_),
    .Y(_07084_));
 AND2x2_ASAP7_75t_R _14062_ (.A(_05224_),
    .B(_01009_),
    .Y(_07085_));
 AO21x1_ASAP7_75t_R _14063_ (.A1(_03840_),
    .A2(_01008_),
    .B(_07085_),
    .Y(_07086_));
 AND2x2_ASAP7_75t_R _14064_ (.A(_05224_),
    .B(_01013_),
    .Y(_07087_));
 AO21x1_ASAP7_75t_R _14065_ (.A1(_03840_),
    .A2(_01012_),
    .B(_07087_),
    .Y(_07088_));
 OAI22x1_ASAP7_75t_R _14066_ (.A1(_04948_),
    .A2(_07086_),
    .B1(_07088_),
    .B2(_03707_),
    .Y(_07089_));
 AND4x1_ASAP7_75t_R _14067_ (.A(_05331_),
    .B(_07032_),
    .C(_03814_),
    .D(_03803_),
    .Y(_07090_));
 OR3x1_ASAP7_75t_R _14068_ (.A(_05235_),
    .B(_07089_),
    .C(_07090_),
    .Y(_07091_));
 AO221x2_ASAP7_75t_R _14069_ (.A1(_07082_),
    .A2(_06578_),
    .B1(_07084_),
    .B2(_06575_),
    .C(_07091_),
    .Y(_07092_));
 OA211x2_ASAP7_75t_R _14070_ (.A1(_03524_),
    .A2(_03880_),
    .B(_03887_),
    .C(_00999_),
    .Y(_07093_));
 AO21x1_ASAP7_75t_R _14071_ (.A1(_00998_),
    .A2(_03587_),
    .B(_07093_),
    .Y(_07094_));
 AND3x1_ASAP7_75t_R _14072_ (.A(_03844_),
    .B(_03845_),
    .C(_01001_),
    .Y(_07095_));
 AO21x1_ASAP7_75t_R _14073_ (.A1(_01000_),
    .A2(_04434_),
    .B(_07095_),
    .Y(_07096_));
 AND4x1_ASAP7_75t_R _14074_ (.A(_06285_),
    .B(_03557_),
    .C(_03783_),
    .D(_07096_),
    .Y(_07097_));
 AO21x1_ASAP7_75t_R _14075_ (.A1(_03889_),
    .A2(_07094_),
    .B(_07097_),
    .Y(_07098_));
 NAND2x2_ASAP7_75t_R _14076_ (.A(_03773_),
    .B(_07098_),
    .Y(_07099_));
 OA211x2_ASAP7_75t_R _14077_ (.A1(_03524_),
    .A2(_03880_),
    .B(_03887_),
    .C(_01003_),
    .Y(_07100_));
 AO21x1_ASAP7_75t_R _14078_ (.A1(_01002_),
    .A2(_03587_),
    .B(_07100_),
    .Y(_07101_));
 OA222x2_ASAP7_75t_R _14079_ (.A1(_01004_),
    .A2(_05640_),
    .B1(_03587_),
    .B2(_01005_),
    .C1(_03783_),
    .C2(_03820_),
    .Y(_07102_));
 AO21x1_ASAP7_75t_R _14080_ (.A1(_04792_),
    .A2(_07101_),
    .B(_07102_),
    .Y(_07103_));
 AOI21x1_ASAP7_75t_R _14081_ (.A1(_03792_),
    .A2(_07103_),
    .B(_04452_),
    .Y(_07104_));
 AO32x1_ASAP7_75t_R _14082_ (.A1(_01024_),
    .A2(_03862_),
    .A3(_03831_),
    .B1(_05233_),
    .B2(_01025_),
    .Y(_07105_));
 AO21x1_ASAP7_75t_R _14083_ (.A1(_03844_),
    .A2(_05224_),
    .B(_01028_),
    .Y(_07106_));
 OA21x2_ASAP7_75t_R _14084_ (.A1(_01029_),
    .A2(_04595_),
    .B(_07106_),
    .Y(_07107_));
 OA21x2_ASAP7_75t_R _14085_ (.A1(_03820_),
    .A2(_03817_),
    .B(_07107_),
    .Y(_07108_));
 OAI21x1_ASAP7_75t_R _14086_ (.A1(_07105_),
    .A2(_07108_),
    .B(_06606_),
    .Y(_07109_));
 OA211x2_ASAP7_75t_R _14087_ (.A1(_03524_),
    .A2(_03880_),
    .B(_04921_),
    .C(_01023_),
    .Y(_07110_));
 AOI21x1_ASAP7_75t_R _14088_ (.A1(_01022_),
    .A2(_03879_),
    .B(_07110_),
    .Y(_07111_));
 NAND2x1_ASAP7_75t_R _14089_ (.A(_01027_),
    .B(_03886_),
    .Y(_07112_));
 NAND2x1_ASAP7_75t_R _14090_ (.A(_01026_),
    .B(_03805_),
    .Y(_07113_));
 AND5x1_ASAP7_75t_R _14091_ (.A(_03742_),
    .B(_03678_),
    .C(_06097_),
    .D(_07112_),
    .E(_07113_),
    .Y(_07114_));
 AO211x2_ASAP7_75t_R _14092_ (.A1(_06094_),
    .A2(_07111_),
    .B(_07114_),
    .C(_06101_),
    .Y(_07115_));
 OAI22x1_ASAP7_75t_R _14093_ (.A1(_04930_),
    .A2(_01014_),
    .B1(_01015_),
    .B2(_03711_),
    .Y(_07116_));
 AO22x1_ASAP7_75t_R _14094_ (.A1(_04935_),
    .A2(_07068_),
    .B1(_07116_),
    .B2(_03632_),
    .Y(_07117_));
 AND2x2_ASAP7_75t_R _14095_ (.A(_01016_),
    .B(_03711_),
    .Y(_07118_));
 AOI221x1_ASAP7_75t_R _14096_ (.A1(_01017_),
    .A2(_03887_),
    .B1(_03803_),
    .B2(_03862_),
    .C(_07118_),
    .Y(_07119_));
 OR3x1_ASAP7_75t_R _14097_ (.A(_05713_),
    .B(_07117_),
    .C(_07119_),
    .Y(_07120_));
 NAND2x1_ASAP7_75t_R _14098_ (.A(_01019_),
    .B(_03886_),
    .Y(_07121_));
 NAND2x1_ASAP7_75t_R _14099_ (.A(_01018_),
    .B(_03761_),
    .Y(_07122_));
 AND4x1_ASAP7_75t_R _14100_ (.A(_03705_),
    .B(_03888_),
    .C(_07121_),
    .D(_07122_),
    .Y(_07123_));
 AND2x2_ASAP7_75t_R _14101_ (.A(_01020_),
    .B(_03761_),
    .Y(_07124_));
 AOI221x1_ASAP7_75t_R _14102_ (.A1(_01021_),
    .A2(_03774_),
    .B1(_03776_),
    .B2(_03804_),
    .C(_07124_),
    .Y(_07125_));
 OR4x1_ASAP7_75t_R _14103_ (.A(_05227_),
    .B(_05698_),
    .C(_07123_),
    .D(_07125_),
    .Y(_07126_));
 AND5x2_ASAP7_75t_R _14104_ (.A(_03907_),
    .B(_07109_),
    .C(_07115_),
    .D(_07120_),
    .E(_07126_),
    .Y(_07127_));
 AO31x2_ASAP7_75t_R _14105_ (.A1(_07092_),
    .A2(_07099_),
    .A3(_07104_),
    .B(_07127_),
    .Y(_07128_));
 BUFx6f_ASAP7_75t_R _14106_ (.A(_07128_),
    .Y(_10092_));
 INVx1_ASAP7_75t_R _14107_ (.A(_10092_),
    .Y(_10094_));
 AND3x1_ASAP7_75t_R _14108_ (.A(_03509_),
    .B(_03557_),
    .C(_03547_),
    .Y(_07129_));
 INVx2_ASAP7_75t_R _14109_ (.A(net29),
    .Y(_07130_));
 OAI21x1_ASAP7_75t_R _14110_ (.A1(_03415_),
    .A2(_07130_),
    .B(_03566_),
    .Y(_07131_));
 AO32x1_ASAP7_75t_R _14111_ (.A1(_03504_),
    .A2(_04412_),
    .A3(_07129_),
    .B1(_07131_),
    .B2(_03503_),
    .Y(_07132_));
 BUFx4f_ASAP7_75t_R _14112_ (.A(_07132_),
    .Y(_09945_));
 AND2x2_ASAP7_75t_R _14113_ (.A(_03387_),
    .B(_01061_),
    .Y(_07133_));
 AO21x1_ASAP7_75t_R _14114_ (.A1(_03424_),
    .A2(_01059_),
    .B(_07133_),
    .Y(_07134_));
 AO221x1_ASAP7_75t_R _14115_ (.A1(_03391_),
    .A2(_01062_),
    .B1(_04019_),
    .B2(_01060_),
    .C(_03421_),
    .Y(_07135_));
 OA211x2_ASAP7_75t_R _14116_ (.A1(_03400_),
    .A2(_07134_),
    .B(_07135_),
    .C(_03411_),
    .Y(_07136_));
 AND2x2_ASAP7_75t_R _14117_ (.A(_03387_),
    .B(_01057_),
    .Y(_07137_));
 AO21x1_ASAP7_75t_R _14118_ (.A1(_03424_),
    .A2(_01055_),
    .B(_07137_),
    .Y(_07138_));
 AO221x1_ASAP7_75t_R _14119_ (.A1(_03391_),
    .A2(_01058_),
    .B1(_04019_),
    .B2(_01056_),
    .C(_03406_),
    .Y(_07139_));
 OA211x2_ASAP7_75t_R _14120_ (.A1(_06839_),
    .A2(_07138_),
    .B(_07139_),
    .C(_03418_),
    .Y(_07140_));
 OA21x2_ASAP7_75t_R _14121_ (.A1(_07136_),
    .A2(_07140_),
    .B(_06809_),
    .Y(_07141_));
 AND2x2_ASAP7_75t_R _14122_ (.A(_03387_),
    .B(_01045_),
    .Y(_07142_));
 AO21x1_ASAP7_75t_R _14123_ (.A1(_03424_),
    .A2(_01043_),
    .B(_07142_),
    .Y(_07143_));
 AO22x1_ASAP7_75t_R _14124_ (.A1(_01046_),
    .A2(_03960_),
    .B1(_07143_),
    .B2(_03407_),
    .Y(_07144_));
 AO21x1_ASAP7_75t_R _14125_ (.A1(_01044_),
    .A2(_03963_),
    .B(_03449_),
    .Y(_07145_));
 OR2x2_ASAP7_75t_R _14126_ (.A(_03387_),
    .B(_03411_),
    .Y(_07146_));
 AO221x1_ASAP7_75t_R _14127_ (.A1(_03421_),
    .A2(_01039_),
    .B1(_01040_),
    .B2(_03987_),
    .C(_07146_),
    .Y(_07147_));
 AND2x2_ASAP7_75t_R _14128_ (.A(net12),
    .B(_01042_),
    .Y(_07148_));
 AO21x1_ASAP7_75t_R _14129_ (.A1(_03421_),
    .A2(_01041_),
    .B(_07148_),
    .Y(_07149_));
 NAND2x1_ASAP7_75t_R _14130_ (.A(_03388_),
    .B(_03418_),
    .Y(_07150_));
 OA21x2_ASAP7_75t_R _14131_ (.A1(_07149_),
    .A2(_07150_),
    .B(_03383_),
    .Y(_07151_));
 OA211x2_ASAP7_75t_R _14132_ (.A1(_07144_),
    .A2(_07145_),
    .B(_07147_),
    .C(_07151_),
    .Y(_07152_));
 OR3x4_ASAP7_75t_R _14133_ (.A(_03995_),
    .B(_07141_),
    .C(_07152_),
    .Y(_07153_));
 AND2x2_ASAP7_75t_R _14134_ (.A(_03388_),
    .B(_01049_),
    .Y(_07154_));
 AO21x1_ASAP7_75t_R _14135_ (.A1(_03386_),
    .A2(_01047_),
    .B(_07154_),
    .Y(_07155_));
 AO221x1_ASAP7_75t_R _14136_ (.A1(_03392_),
    .A2(_01050_),
    .B1(_04019_),
    .B2(_01048_),
    .C(_03407_),
    .Y(_07156_));
 OAI21x1_ASAP7_75t_R _14137_ (.A1(_06840_),
    .A2(_07155_),
    .B(_07156_),
    .Y(_07157_));
 INVx2_ASAP7_75t_R _14138_ (.A(_01054_),
    .Y(_07158_));
 NOR2x1_ASAP7_75t_R _14139_ (.A(_03388_),
    .B(_01052_),
    .Y(_07159_));
 AO21x1_ASAP7_75t_R _14140_ (.A1(_03392_),
    .A2(_07158_),
    .B(_07159_),
    .Y(_07160_));
 INVx2_ASAP7_75t_R _14141_ (.A(_01051_),
    .Y(_07161_));
 NAND2x1_ASAP7_75t_R _14142_ (.A(_03391_),
    .B(_01053_),
    .Y(_07162_));
 OA211x2_ASAP7_75t_R _14143_ (.A1(_03432_),
    .A2(_07161_),
    .B(_07162_),
    .C(_03421_),
    .Y(_07163_));
 AO21x1_ASAP7_75t_R _14144_ (.A1(_03400_),
    .A2(_07160_),
    .B(_07163_),
    .Y(_07164_));
 AO32x1_ASAP7_75t_R _14145_ (.A1(_04296_),
    .A2(_06809_),
    .A3(_07157_),
    .B1(_07164_),
    .B2(_07042_),
    .Y(_07165_));
 NOR2x1_ASAP7_75t_R _14146_ (.A(_03412_),
    .B(_06809_),
    .Y(_07166_));
 AND2x2_ASAP7_75t_R _14147_ (.A(_03399_),
    .B(_01034_),
    .Y(_07167_));
 AO21x1_ASAP7_75t_R _14148_ (.A1(_03407_),
    .A2(_01033_),
    .B(_07167_),
    .Y(_07168_));
 AND4x1_ASAP7_75t_R _14149_ (.A(_06839_),
    .B(_03424_),
    .C(_03374_),
    .D(_01032_),
    .Y(_07169_));
 AOI221x1_ASAP7_75t_R _14150_ (.A1(_01031_),
    .A2(_03405_),
    .B1(_04412_),
    .B2(_07168_),
    .C(_07169_),
    .Y(_07170_));
 AND3x1_ASAP7_75t_R _14151_ (.A(_03400_),
    .B(_03443_),
    .C(_01036_),
    .Y(_07171_));
 AO21x1_ASAP7_75t_R _14152_ (.A1(_03407_),
    .A2(_01035_),
    .B(_03426_),
    .Y(_07172_));
 AND2x2_ASAP7_75t_R _14153_ (.A(_06839_),
    .B(_01038_),
    .Y(_07173_));
 AO21x1_ASAP7_75t_R _14154_ (.A1(_03422_),
    .A2(_01037_),
    .B(_07173_),
    .Y(_07174_));
 OAI22x1_ASAP7_75t_R _14155_ (.A1(_07171_),
    .A2(_07172_),
    .B1(_07174_),
    .B2(_03952_),
    .Y(_07175_));
 AND2x2_ASAP7_75t_R _14156_ (.A(_03412_),
    .B(_03429_),
    .Y(_07176_));
 AO22x1_ASAP7_75t_R _14157_ (.A1(_07166_),
    .A2(_07170_),
    .B1(_07175_),
    .B2(_07176_),
    .Y(_07177_));
 OAI21x1_ASAP7_75t_R _14158_ (.A1(_07165_),
    .A2(_07177_),
    .B(_07072_),
    .Y(_07178_));
 AND2x6_ASAP7_75t_R _14159_ (.A(_07153_),
    .B(_07178_),
    .Y(_07179_));
 CKINVDCx9p33_ASAP7_75t_R _14160_ (.A(_07179_),
    .Y(net110));
 NAND3x2_ASAP7_75t_R _14161_ (.B(_07153_),
    .C(_07178_),
    .Y(_07180_),
    .A(_04058_));
 OR2x2_ASAP7_75t_R _14162_ (.A(_04057_),
    .B(_09945_),
    .Y(_07181_));
 BUFx6f_ASAP7_75t_R _14163_ (.A(_07181_),
    .Y(_07182_));
 AND2x6_ASAP7_75t_R _14164_ (.A(_07180_),
    .B(_07182_),
    .Y(_07183_));
 BUFx10_ASAP7_75t_R _14165_ (.A(_07183_),
    .Y(_07184_));
 BUFx6f_ASAP7_75t_R _14166_ (.A(_07184_),
    .Y(_07185_));
 BUFx6f_ASAP7_75t_R _14167_ (.A(_07185_),
    .Y(_07186_));
 XNOR2x2_ASAP7_75t_R _14168_ (.A(_03913_),
    .B(_07186_),
    .Y(_09942_));
 INVx1_ASAP7_75t_R _14169_ (.A(_09942_),
    .Y(_10098_));
 NOR2x1_ASAP7_75t_R _14170_ (.A(_01034_),
    .B(_03587_),
    .Y(_07187_));
 OAI21x1_ASAP7_75t_R _14171_ (.A1(_01033_),
    .A2(_05640_),
    .B(_03901_),
    .Y(_07188_));
 OAI21x1_ASAP7_75t_R _14172_ (.A1(_01032_),
    .A2(_03587_),
    .B(_03601_),
    .Y(_07189_));
 OA21x2_ASAP7_75t_R _14173_ (.A1(_07187_),
    .A2(_07188_),
    .B(_07189_),
    .Y(_07190_));
 AND2x2_ASAP7_75t_R _14174_ (.A(_04938_),
    .B(_01060_),
    .Y(_07191_));
 AO21x1_ASAP7_75t_R _14175_ (.A1(_04831_),
    .A2(_01056_),
    .B(_07191_),
    .Y(_07192_));
 AO22x1_ASAP7_75t_R _14176_ (.A1(_01059_),
    .A2(_04800_),
    .B1(_07192_),
    .B2(_05215_),
    .Y(_07193_));
 NAND2x1_ASAP7_75t_R _14177_ (.A(_03377_),
    .B(_07193_),
    .Y(_07194_));
 AO21x1_ASAP7_75t_R _14178_ (.A1(_03825_),
    .A2(_07194_),
    .B(_04806_),
    .Y(_07195_));
 NAND2x1_ASAP7_75t_R _14179_ (.A(_01055_),
    .B(_03811_),
    .Y(_07196_));
 AND3x1_ASAP7_75t_R _14180_ (.A(_01057_),
    .B(_03777_),
    .C(_03831_),
    .Y(_07197_));
 AOI221x1_ASAP7_75t_R _14181_ (.A1(_01062_),
    .A2(_05230_),
    .B1(_04476_),
    .B2(_01061_),
    .C(_07197_),
    .Y(_07198_));
 AOI21x1_ASAP7_75t_R _14182_ (.A1(_01058_),
    .A2(_05233_),
    .B(_03826_),
    .Y(_07199_));
 AO221x2_ASAP7_75t_R _14183_ (.A1(_07195_),
    .A2(_07196_),
    .B1(_07198_),
    .B2(_07199_),
    .C(_04468_),
    .Y(_07200_));
 OA21x2_ASAP7_75t_R _14184_ (.A1(_04806_),
    .A2(_05698_),
    .B(_03907_),
    .Y(_07201_));
 OR3x1_ASAP7_75t_R _14185_ (.A(_07161_),
    .B(_03780_),
    .C(_03765_),
    .Y(_07202_));
 OAI21x1_ASAP7_75t_R _14186_ (.A1(_03820_),
    .A2(_03783_),
    .B(_01053_),
    .Y(_07203_));
 AND4x1_ASAP7_75t_R _14187_ (.A(_04929_),
    .B(_03907_),
    .C(_07202_),
    .D(_07203_),
    .Y(_07204_));
 NAND2x1_ASAP7_75t_R _14188_ (.A(_01052_),
    .B(_04804_),
    .Y(_07205_));
 OA211x2_ASAP7_75t_R _14189_ (.A1(_03756_),
    .A2(_07205_),
    .B(_03906_),
    .C(_03882_),
    .Y(_07206_));
 OA21x2_ASAP7_75t_R _14190_ (.A1(_07158_),
    .A2(_05218_),
    .B(_07206_),
    .Y(_07207_));
 NOR2x1_ASAP7_75t_R _14191_ (.A(_01048_),
    .B(_03781_),
    .Y(_07208_));
 OR4x1_ASAP7_75t_R _14192_ (.A(_03780_),
    .B(_03765_),
    .C(_03611_),
    .D(_07208_),
    .Y(_07209_));
 AND3x1_ASAP7_75t_R _14193_ (.A(_03623_),
    .B(_03624_),
    .C(_01050_),
    .Y(_07210_));
 AOI21x1_ASAP7_75t_R _14194_ (.A1(_01049_),
    .A2(_03781_),
    .B(_07210_),
    .Y(_07211_));
 OR4x1_ASAP7_75t_R _14195_ (.A(_03780_),
    .B(_03802_),
    .C(_03611_),
    .D(_07211_),
    .Y(_07212_));
 INVx1_ASAP7_75t_R _14196_ (.A(_01047_),
    .Y(_07213_));
 AO32x1_ASAP7_75t_R _14197_ (.A1(_03655_),
    .A2(_07209_),
    .A3(_07212_),
    .B1(_03703_),
    .B2(_07213_),
    .Y(_07214_));
 OA31x2_ASAP7_75t_R _14198_ (.A1(_07201_),
    .A2(_07204_),
    .A3(_07207_),
    .B1(_07214_),
    .Y(_07215_));
 AND3x1_ASAP7_75t_R _14199_ (.A(_03844_),
    .B(_03845_),
    .C(_01036_),
    .Y(_07216_));
 AO21x1_ASAP7_75t_R _14200_ (.A1(_01035_),
    .A2(_04434_),
    .B(_07216_),
    .Y(_07217_));
 AND2x2_ASAP7_75t_R _14201_ (.A(_01037_),
    .B(_03761_),
    .Y(_07218_));
 AO221x1_ASAP7_75t_R _14202_ (.A1(_01038_),
    .A2(_03774_),
    .B1(_03776_),
    .B2(_03777_),
    .C(_07218_),
    .Y(_07219_));
 OA21x2_ASAP7_75t_R _14203_ (.A1(_03795_),
    .A2(_07217_),
    .B(_07219_),
    .Y(_07220_));
 OR3x1_ASAP7_75t_R _14204_ (.A(_01042_),
    .B(_03782_),
    .C(_04948_),
    .Y(_07221_));
 OR3x1_ASAP7_75t_R _14205_ (.A(_01041_),
    .B(_03774_),
    .C(_04948_),
    .Y(_07222_));
 AND2x2_ASAP7_75t_R _14206_ (.A(_01045_),
    .B(_03781_),
    .Y(_07223_));
 AO221x1_ASAP7_75t_R _14207_ (.A1(_01046_),
    .A2(_03882_),
    .B1(_03707_),
    .B2(_03873_),
    .C(_07223_),
    .Y(_07224_));
 AND4x1_ASAP7_75t_R _14208_ (.A(_03868_),
    .B(_07221_),
    .C(_07222_),
    .D(_07224_),
    .Y(_07225_));
 AND2x2_ASAP7_75t_R _14209_ (.A(_03610_),
    .B(_01044_),
    .Y(_07226_));
 AO21x1_ASAP7_75t_R _14210_ (.A1(_04609_),
    .A2(_01040_),
    .B(_07226_),
    .Y(_07227_));
 AO21x1_ASAP7_75t_R _14211_ (.A1(_05332_),
    .A2(_01043_),
    .B(_04460_),
    .Y(_07228_));
 OA211x2_ASAP7_75t_R _14212_ (.A1(_03629_),
    .A2(_07227_),
    .B(_07228_),
    .C(_04916_),
    .Y(_07229_));
 OR3x1_ASAP7_75t_R _14213_ (.A(_03820_),
    .B(_03783_),
    .C(_07229_),
    .Y(_07230_));
 AO32x1_ASAP7_75t_R _14214_ (.A1(_06285_),
    .A2(_03678_),
    .A3(_07230_),
    .B1(_03750_),
    .B2(_01039_),
    .Y(_07231_));
 AOI221x1_ASAP7_75t_R _14215_ (.A1(_03792_),
    .A2(_07220_),
    .B1(_07225_),
    .B2(_07231_),
    .C(_03907_),
    .Y(_07232_));
 AO21x2_ASAP7_75t_R _14216_ (.A1(_07200_),
    .A2(_07215_),
    .B(_07232_),
    .Y(_07233_));
 AND2x4_ASAP7_75t_R _14217_ (.A(_07190_),
    .B(_07233_),
    .Y(_09941_));
 INVx1_ASAP7_75t_R _14218_ (.A(_09941_),
    .Y(_10097_));
 NAND2x2_ASAP7_75t_R _14219_ (.A(_03576_),
    .B(_03577_),
    .Y(_07234_));
 BUFx4f_ASAP7_75t_R _14220_ (.A(_07234_),
    .Y(_07235_));
 AND3x1_ASAP7_75t_R _14221_ (.A(_07235_),
    .B(_03602_),
    .C(_03770_),
    .Y(_07236_));
 AO21x2_ASAP7_75t_R _14222_ (.A1(_03537_),
    .A2(_03579_),
    .B(_07236_),
    .Y(_09940_));
 INVx1_ASAP7_75t_R _14223_ (.A(_09949_),
    .Y(_09947_));
 INVx1_ASAP7_75t_R _14224_ (.A(_09984_),
    .Y(_09982_));
 INVx1_ASAP7_75t_R _14225_ (.A(_09969_),
    .Y(_09967_));
 BUFx6f_ASAP7_75t_R _14226_ (.A(_03910_),
    .Y(_09955_));
 INVx1_ASAP7_75t_R _14227_ (.A(_10084_),
    .Y(_10082_));
 INVx1_ASAP7_75t_R _14228_ (.A(_10064_),
    .Y(_10062_));
 INVx2_ASAP7_75t_R _14229_ (.A(_10059_),
    .Y(_10057_));
 INVx1_ASAP7_75t_R _14230_ (.A(_10102_),
    .Y(_10100_));
 INVx2_ASAP7_75t_R _14231_ (.A(_10054_),
    .Y(_10052_));
 INVx3_ASAP7_75t_R _14232_ (.A(_10034_),
    .Y(_10032_));
 INVx1_ASAP7_75t_R _14233_ (.A(_10024_),
    .Y(_10022_));
 INVx1_ASAP7_75t_R _14234_ (.A(_10019_),
    .Y(_10017_));
 INVx1_ASAP7_75t_R _14235_ (.A(_09946_),
    .Y(_09943_));
 INVx3_ASAP7_75t_R _14236_ (.A(_10110_),
    .Y(net90));
 INVx4_ASAP7_75t_R _14237_ (.A(_10109_),
    .Y(net87));
 AO21x1_ASAP7_75t_R _14238_ (.A1(_04059_),
    .A2(_06961_),
    .B(_06962_),
    .Y(_07237_));
 BUFx4f_ASAP7_75t_R _14239_ (.A(_07237_),
    .Y(_07238_));
 NAND2x2_ASAP7_75t_R _14240_ (.A(_04596_),
    .B(_03483_),
    .Y(_07239_));
 INVx1_ASAP7_75t_R _14241_ (.A(net4),
    .Y(_07240_));
 OR2x2_ASAP7_75t_R _14242_ (.A(net5),
    .B(_07240_),
    .Y(_07241_));
 OR3x2_ASAP7_75t_R _14243_ (.A(_03526_),
    .B(_07239_),
    .C(_07241_),
    .Y(_07242_));
 BUFx6f_ASAP7_75t_R _14244_ (.A(_07242_),
    .Y(_07243_));
 NAND2x2_ASAP7_75t_R _14245_ (.A(_07238_),
    .B(_07243_),
    .Y(_07244_));
 OAI22x1_ASAP7_75t_R _14246_ (.A1(_03401_),
    .A2(_03417_),
    .B1(_03420_),
    .B2(_03440_),
    .Y(_07245_));
 NOR3x2_ASAP7_75t_R _14247_ (.B(_03462_),
    .C(_03476_),
    .Y(_07246_),
    .A(_03448_));
 OR4x2_ASAP7_75t_R _14248_ (.A(_07245_),
    .B(_07246_),
    .C(_03575_),
    .D(_07074_),
    .Y(_07247_));
 OR3x2_ASAP7_75t_R _14249_ (.A(_10106_),
    .B(_04058_),
    .C(_07024_),
    .Y(_07248_));
 NAND2x2_ASAP7_75t_R _14250_ (.A(_07247_),
    .B(_07248_),
    .Y(_07249_));
 NAND3x2_ASAP7_75t_R _14251_ (.B(_07190_),
    .C(_07233_),
    .Y(_07250_),
    .A(_07183_));
 BUFx6f_ASAP7_75t_R _14252_ (.A(_07180_),
    .Y(_07251_));
 NAND2x2_ASAP7_75t_R _14253_ (.A(_07251_),
    .B(_07182_),
    .Y(_07252_));
 NAND2x2_ASAP7_75t_R _14254_ (.A(_07012_),
    .B(_07252_),
    .Y(_07253_));
 AND3x4_ASAP7_75t_R _14255_ (.A(_04058_),
    .B(_07153_),
    .C(_07178_),
    .Y(_07254_));
 NOR2x2_ASAP7_75t_R _14256_ (.A(_04058_),
    .B(_09945_),
    .Y(_07255_));
 OA222x2_ASAP7_75t_R _14257_ (.A1(_06588_),
    .A2(_06601_),
    .B1(_06607_),
    .B2(_06624_),
    .C1(_07254_),
    .C2(_07255_),
    .Y(_07256_));
 AO21x1_ASAP7_75t_R _14258_ (.A1(_10079_),
    .A2(_07183_),
    .B(_07256_),
    .Y(_07257_));
 AND2x2_ASAP7_75t_R _14259_ (.A(_03552_),
    .B(_03575_),
    .Y(_07258_));
 AO32x2_ASAP7_75t_R _14260_ (.A1(_03478_),
    .A2(_04059_),
    .A3(_07075_),
    .B1(_07258_),
    .B2(_07024_),
    .Y(_07259_));
 AO32x1_ASAP7_75t_R _14261_ (.A1(_07249_),
    .A2(_07250_),
    .A3(_07253_),
    .B1(_07257_),
    .B2(_07259_),
    .Y(_07260_));
 OA21x2_ASAP7_75t_R _14262_ (.A1(_07245_),
    .A2(_07246_),
    .B(_04058_),
    .Y(_07261_));
 AND3x1_ASAP7_75t_R _14263_ (.A(_10106_),
    .B(_03575_),
    .C(_07024_),
    .Y(_07262_));
 AO21x2_ASAP7_75t_R _14264_ (.A1(_07261_),
    .A2(_07074_),
    .B(_07262_),
    .Y(_07263_));
 OA222x2_ASAP7_75t_R _14265_ (.A1(_06681_),
    .A2(_06691_),
    .B1(_06702_),
    .B2(_06714_),
    .C1(_07254_),
    .C2(_07255_),
    .Y(_07264_));
 AO21x2_ASAP7_75t_R _14266_ (.A1(_10084_),
    .A2(_07183_),
    .B(_07264_),
    .Y(_07265_));
 AO211x2_ASAP7_75t_R _14267_ (.A1(_03441_),
    .A2(_03477_),
    .B(_03915_),
    .C(_07074_),
    .Y(_07266_));
 OR3x2_ASAP7_75t_R _14268_ (.A(_03552_),
    .B(_04058_),
    .C(_07024_),
    .Y(_07267_));
 AND2x2_ASAP7_75t_R _14269_ (.A(_07266_),
    .B(_07267_),
    .Y(_07268_));
 NOR3x1_ASAP7_75t_R _14270_ (.A(_07128_),
    .B(_07184_),
    .C(_07268_),
    .Y(_07269_));
 BUFx6f_ASAP7_75t_R _14271_ (.A(_07252_),
    .Y(_07270_));
 AOI211x1_ASAP7_75t_R _14272_ (.A1(_03602_),
    .A2(_03770_),
    .B(_07270_),
    .C(_07268_),
    .Y(_07271_));
 AO211x2_ASAP7_75t_R _14273_ (.A1(_07263_),
    .A2(_07265_),
    .B(_07269_),
    .C(_07271_),
    .Y(_07272_));
 OR2x2_ASAP7_75t_R _14274_ (.A(_07260_),
    .B(_07272_),
    .Y(_07273_));
 INVx2_ASAP7_75t_R _14275_ (.A(_07241_),
    .Y(_07274_));
 AND3x4_ASAP7_75t_R _14276_ (.A(_03559_),
    .B(_05755_),
    .C(_07274_),
    .Y(_07275_));
 BUFx6f_ASAP7_75t_R _14277_ (.A(_07275_),
    .Y(_07276_));
 AND2x4_ASAP7_75t_R _14278_ (.A(_04169_),
    .B(_07276_),
    .Y(_07277_));
 NAND2x1_ASAP7_75t_R _14279_ (.A(_03911_),
    .B(_07277_),
    .Y(_07278_));
 AND2x2_ASAP7_75t_R _14280_ (.A(_06865_),
    .B(_07278_),
    .Y(_07279_));
 OAI21x1_ASAP7_75t_R _14281_ (.A1(_07244_),
    .A2(_07273_),
    .B(_07279_),
    .Y(_07280_));
 OA21x2_ASAP7_75t_R _14282_ (.A1(_05342_),
    .A2(_05345_),
    .B(_07263_),
    .Y(_07281_));
 AO32x1_ASAP7_75t_R _14283_ (.A1(_07235_),
    .A2(_10029_),
    .A3(_07077_),
    .B1(_07259_),
    .B2(_10002_),
    .Y(_07282_));
 AO221x1_ASAP7_75t_R _14284_ (.A1(_09997_),
    .A2(_07263_),
    .B1(_07259_),
    .B2(_09994_),
    .C(_07183_),
    .Y(_07283_));
 OA31x2_ASAP7_75t_R _14285_ (.A1(_07270_),
    .A2(_07281_),
    .A3(_07282_),
    .B1(_07283_),
    .Y(_07284_));
 AO21x1_ASAP7_75t_R _14286_ (.A1(_03441_),
    .A2(_03477_),
    .B(_07074_),
    .Y(_07285_));
 OA22x2_ASAP7_75t_R _14287_ (.A1(_07013_),
    .A2(_07018_),
    .B1(_07019_),
    .B2(_07021_),
    .Y(_07286_));
 OR4x1_ASAP7_75t_R _14288_ (.A(_03552_),
    .B(_04058_),
    .C(_09945_),
    .D(_07286_),
    .Y(_07287_));
 OAI21x1_ASAP7_75t_R _14289_ (.A1(_07251_),
    .A2(_07285_),
    .B(_07287_),
    .Y(_07288_));
 OA211x2_ASAP7_75t_R _14290_ (.A1(_07254_),
    .A2(_07255_),
    .B(_03576_),
    .C(_03577_),
    .Y(_07289_));
 BUFx3_ASAP7_75t_R _14291_ (.A(_07289_),
    .Y(_07290_));
 AO32x1_ASAP7_75t_R _14292_ (.A1(_03478_),
    .A2(_04058_),
    .A3(net110),
    .B1(_07258_),
    .B2(_09945_),
    .Y(_07291_));
 AO32x1_ASAP7_75t_R _14293_ (.A1(_05424_),
    .A2(_05446_),
    .A3(_07290_),
    .B1(_07291_),
    .B2(_10024_),
    .Y(_07292_));
 AO221x1_ASAP7_75t_R _14294_ (.A1(_10019_),
    .A2(_07288_),
    .B1(_07292_),
    .B2(_07077_),
    .C(_06963_),
    .Y(_07293_));
 AOI211x1_ASAP7_75t_R _14295_ (.A1(_07266_),
    .A2(_07267_),
    .B(_07254_),
    .C(_07255_),
    .Y(_07294_));
 AO32x1_ASAP7_75t_R _14296_ (.A1(_10049_),
    .A2(_07183_),
    .A3(_07263_),
    .B1(_07294_),
    .B2(_06524_),
    .Y(_07295_));
 NAND2x2_ASAP7_75t_R _14297_ (.A(_06037_),
    .B(_06026_),
    .Y(_07296_));
 NAND3x2_ASAP7_75t_R _14298_ (.B(_06013_),
    .C(_06017_),
    .Y(_07297_),
    .A(_06002_));
 AO21x2_ASAP7_75t_R _14299_ (.A1(_03915_),
    .A2(_07024_),
    .B(_07076_),
    .Y(_07298_));
 AND4x1_ASAP7_75t_R _14300_ (.A(_07296_),
    .B(_07297_),
    .C(_07298_),
    .D(_07291_),
    .Y(_07299_));
 OA211x2_ASAP7_75t_R _14301_ (.A1(_06207_),
    .A2(_06238_),
    .B(_07252_),
    .C(_07249_),
    .Y(_07300_));
 OR3x4_ASAP7_75t_R _14302_ (.A(_06301_),
    .B(_06307_),
    .C(_06312_),
    .Y(_07301_));
 OR4x2_ASAP7_75t_R _14303_ (.A(_04452_),
    .B(_06290_),
    .C(_06326_),
    .D(_06330_),
    .Y(_07302_));
 AO33x2_ASAP7_75t_R _14304_ (.A1(_06431_),
    .A2(_07183_),
    .A3(_07249_),
    .B1(_07288_),
    .B2(_07301_),
    .B3(_07302_),
    .Y(_07303_));
 OR4x2_ASAP7_75t_R _14305_ (.A(_07295_),
    .B(_07299_),
    .C(_07300_),
    .D(_07303_),
    .Y(_07304_));
 AND2x2_ASAP7_75t_R _14306_ (.A(_07298_),
    .B(_07290_),
    .Y(_07305_));
 AOI21x1_ASAP7_75t_R _14307_ (.A1(_07261_),
    .A2(_07075_),
    .B(_07262_),
    .Y(_07306_));
 NOR3x2_ASAP7_75t_R _14308_ (.B(_07184_),
    .C(_07306_),
    .Y(_07307_),
    .A(_10037_));
 AO211x2_ASAP7_75t_R _14309_ (.A1(_05851_),
    .A2(_07305_),
    .B(_07307_),
    .C(_07238_),
    .Y(_07308_));
 OAI22x1_ASAP7_75t_R _14310_ (.A1(_07284_),
    .A2(_07293_),
    .B1(_07304_),
    .B2(_07308_),
    .Y(_07309_));
 NAND2x2_ASAP7_75t_R _14311_ (.A(_04315_),
    .B(net22),
    .Y(_07310_));
 AND2x6_ASAP7_75t_R _14312_ (.A(_07310_),
    .B(_07275_),
    .Y(_07311_));
 AND2x4_ASAP7_75t_R _14313_ (.A(_07238_),
    .B(_07311_),
    .Y(_07312_));
 AOI211x1_ASAP7_75t_R _14314_ (.A1(_04601_),
    .A2(_04621_),
    .B(_04630_),
    .C(_07183_),
    .Y(_07313_));
 NAND2x1_ASAP7_75t_R _14315_ (.A(_07266_),
    .B(_07267_),
    .Y(_07314_));
 AO22x1_ASAP7_75t_R _14316_ (.A1(_09964_),
    .A2(_07249_),
    .B1(_07314_),
    .B2(_09959_),
    .Y(_07315_));
 AND2x2_ASAP7_75t_R _14317_ (.A(_09969_),
    .B(_07288_),
    .Y(_07316_));
 AO221x1_ASAP7_75t_R _14318_ (.A1(_07249_),
    .A2(_07313_),
    .B1(_07315_),
    .B2(_07183_),
    .C(_07316_),
    .Y(_07317_));
 AO21x1_ASAP7_75t_R _14319_ (.A1(_04809_),
    .A2(_04847_),
    .B(_07252_),
    .Y(_07318_));
 NAND2x2_ASAP7_75t_R _14320_ (.A(_09994_),
    .B(_07252_),
    .Y(_07319_));
 AO221x1_ASAP7_75t_R _14321_ (.A1(_04914_),
    .A2(_04928_),
    .B1(_07251_),
    .B2(_07182_),
    .C(_04961_),
    .Y(_07320_));
 OA21x2_ASAP7_75t_R _14322_ (.A1(_09979_),
    .A2(_07252_),
    .B(_07320_),
    .Y(_07321_));
 AO32x1_ASAP7_75t_R _14323_ (.A1(_07259_),
    .A2(_07318_),
    .A3(_07319_),
    .B1(_07321_),
    .B2(_07263_),
    .Y(_07322_));
 OR2x2_ASAP7_75t_R _14324_ (.A(_07317_),
    .B(_07322_),
    .Y(_07323_));
 AND2x2_ASAP7_75t_R _14325_ (.A(_03911_),
    .B(_06963_),
    .Y(_07324_));
 AND3x1_ASAP7_75t_R _14326_ (.A(_07298_),
    .B(_07290_),
    .C(_07311_),
    .Y(_07325_));
 AO21x1_ASAP7_75t_R _14327_ (.A1(_07324_),
    .A2(_07325_),
    .B(_06865_),
    .Y(_07326_));
 AO221x1_ASAP7_75t_R _14328_ (.A1(_07243_),
    .A2(_07309_),
    .B1(_07312_),
    .B2(_07323_),
    .C(_07326_),
    .Y(_07327_));
 OAI21x1_ASAP7_75t_R _14329_ (.A1(_03915_),
    .A2(net125),
    .B(_06864_),
    .Y(_07328_));
 AND2x2_ASAP7_75t_R _14330_ (.A(_07328_),
    .B(_07238_),
    .Y(_07329_));
 OA21x2_ASAP7_75t_R _14331_ (.A1(_03911_),
    .A2(_07329_),
    .B(_07277_),
    .Y(_07330_));
 OR3x1_ASAP7_75t_R _14332_ (.A(_06963_),
    .B(_07317_),
    .C(_07322_),
    .Y(_07331_));
 INVx1_ASAP7_75t_R _14333_ (.A(_03483_),
    .Y(_07332_));
 NAND2x1_ASAP7_75t_R _14334_ (.A(_07332_),
    .B(net22),
    .Y(_07333_));
 AND4x2_ASAP7_75t_R _14335_ (.A(_03972_),
    .B(_03559_),
    .C(_07274_),
    .D(_07333_),
    .Y(_07334_));
 NAND2x2_ASAP7_75t_R _14336_ (.A(_03822_),
    .B(_07334_),
    .Y(_07335_));
 BUFx6f_ASAP7_75t_R _14337_ (.A(_07335_),
    .Y(_07336_));
 AO21x1_ASAP7_75t_R _14338_ (.A1(_07330_),
    .A2(_07331_),
    .B(_07336_),
    .Y(_07337_));
 AO21x1_ASAP7_75t_R _14339_ (.A1(_07280_),
    .A2(_07327_),
    .B(_07337_),
    .Y(_07338_));
 BUFx6f_ASAP7_75t_R _14340_ (.A(_07338_),
    .Y(_07339_));
 INVx1_ASAP7_75t_R _14341_ (.A(_00997_),
    .Y(_07340_));
 NOR2x1_ASAP7_75t_R _14342_ (.A(_01030_),
    .B(_01063_),
    .Y(_07341_));
 AND2x2_ASAP7_75t_R _14343_ (.A(_07340_),
    .B(_07341_),
    .Y(_07342_));
 AND2x2_ASAP7_75t_R _14344_ (.A(_07234_),
    .B(_07342_),
    .Y(_07343_));
 OAI21x1_ASAP7_75t_R _14345_ (.A1(_01030_),
    .A2(_01213_),
    .B(_01211_),
    .Y(_07344_));
 AO32x1_ASAP7_75t_R _14346_ (.A1(_03537_),
    .A2(_03578_),
    .A3(_07342_),
    .B1(_07344_),
    .B2(_07340_),
    .Y(_07345_));
 AOI21x1_ASAP7_75t_R _14347_ (.A1(_09949_),
    .A2(_07343_),
    .B(_07345_),
    .Y(_07346_));
 OR3x1_ASAP7_75t_R _14348_ (.A(_00532_),
    .B(_00565_),
    .C(_00599_),
    .Y(_07347_));
 OR2x2_ASAP7_75t_R _14349_ (.A(_00499_),
    .B(_07347_),
    .Y(_07348_));
 OR3x2_ASAP7_75t_R _14350_ (.A(_00433_),
    .B(_00466_),
    .C(_07348_),
    .Y(_07349_));
 OR2x2_ASAP7_75t_R _14351_ (.A(_00632_),
    .B(_00665_),
    .Y(_07350_));
 OR2x2_ASAP7_75t_R _14352_ (.A(_00797_),
    .B(_01067_),
    .Y(_07351_));
 OR4x1_ASAP7_75t_R _14353_ (.A(_00698_),
    .B(_00731_),
    .C(_07350_),
    .D(_07351_),
    .Y(_07352_));
 BUFx3_ASAP7_75t_R _14354_ (.A(_00964_),
    .Y(_07353_));
 OR2x4_ASAP7_75t_R _14355_ (.A(_00897_),
    .B(_00931_),
    .Y(_07354_));
 OR4x1_ASAP7_75t_R _14356_ (.A(_00830_),
    .B(_00864_),
    .C(_07353_),
    .D(_07354_),
    .Y(_07355_));
 OR2x2_ASAP7_75t_R _14357_ (.A(_07352_),
    .B(_07355_),
    .Y(_07356_));
 OR2x2_ASAP7_75t_R _14358_ (.A(_07349_),
    .B(_07356_),
    .Y(_07357_));
 OA21x2_ASAP7_75t_R _14359_ (.A1(_00830_),
    .A2(_00863_),
    .B(_01201_),
    .Y(_07358_));
 OA21x2_ASAP7_75t_R _14360_ (.A1(_00797_),
    .A2(_07358_),
    .B(_00796_),
    .Y(_07359_));
 OA21x2_ASAP7_75t_R _14361_ (.A1(_01067_),
    .A2(_07359_),
    .B(_01215_),
    .Y(_07360_));
 OA21x2_ASAP7_75t_R _14362_ (.A1(_00731_),
    .A2(_07360_),
    .B(_01198_),
    .Y(_07361_));
 OA21x2_ASAP7_75t_R _14363_ (.A1(_00698_),
    .A2(_07361_),
    .B(_01196_),
    .Y(_07362_));
 OA21x2_ASAP7_75t_R _14364_ (.A1(_00632_),
    .A2(_01194_),
    .B(_01192_),
    .Y(_07363_));
 OA21x2_ASAP7_75t_R _14365_ (.A1(_07350_),
    .A2(_07362_),
    .B(_07363_),
    .Y(_07364_));
 OA21x2_ASAP7_75t_R _14366_ (.A1(_07353_),
    .A2(_01209_),
    .B(_01207_),
    .Y(_07365_));
 OA21x2_ASAP7_75t_R _14367_ (.A1(_00897_),
    .A2(_00930_),
    .B(_01204_),
    .Y(_07366_));
 OA21x2_ASAP7_75t_R _14368_ (.A1(_07354_),
    .A2(_07365_),
    .B(_07366_),
    .Y(_07367_));
 OR3x1_ASAP7_75t_R _14369_ (.A(_00830_),
    .B(_00864_),
    .C(_07367_),
    .Y(_07368_));
 OR2x2_ASAP7_75t_R _14370_ (.A(_07368_),
    .B(_07352_),
    .Y(_07369_));
 AO21x2_ASAP7_75t_R _14371_ (.A1(_07364_),
    .A2(_07369_),
    .B(_07349_),
    .Y(_07370_));
 OAI21x1_ASAP7_75t_R _14372_ (.A1(_07346_),
    .A2(_07357_),
    .B(_07370_),
    .Y(_07371_));
 INVx1_ASAP7_75t_R _14373_ (.A(_03501_),
    .Y(_07372_));
 AO21x1_ASAP7_75t_R _14374_ (.A1(_03530_),
    .A2(_03557_),
    .B(_07372_),
    .Y(_07373_));
 XOR2x1_ASAP7_75t_R _14375_ (.A(net6),
    .Y(_07374_),
    .B(net4));
 OA21x2_ASAP7_75t_R _14376_ (.A1(_03483_),
    .A2(net22),
    .B(_04596_),
    .Y(_07375_));
 OA21x2_ASAP7_75t_R _14377_ (.A1(_03528_),
    .A2(_07374_),
    .B(_07375_),
    .Y(_07376_));
 NOR2x1_ASAP7_75t_R _14378_ (.A(_07373_),
    .B(_07376_),
    .Y(_07377_));
 OA211x2_ASAP7_75t_R _14379_ (.A1(_07239_),
    .A2(_07274_),
    .B(_03559_),
    .C(_07373_),
    .Y(_07378_));
 NOR2x1_ASAP7_75t_R _14380_ (.A(_03483_),
    .B(_03534_),
    .Y(_07379_));
 OA21x2_ASAP7_75t_R _14381_ (.A1(_05852_),
    .A2(_07379_),
    .B(_03526_),
    .Y(_07380_));
 OR4x2_ASAP7_75t_R _14382_ (.A(_03519_),
    .B(_07377_),
    .C(_07378_),
    .D(_07380_),
    .Y(_07381_));
 NAND2x1_ASAP7_75t_R _14383_ (.A(_03483_),
    .B(net4),
    .Y(_07382_));
 AND5x2_ASAP7_75t_R _14384_ (.A(_06806_),
    .B(_03559_),
    .C(_03532_),
    .D(_05853_),
    .E(_07382_),
    .Y(_07383_));
 INVx1_ASAP7_75t_R _14385_ (.A(_07383_),
    .Y(_07384_));
 AND2x2_ASAP7_75t_R _14386_ (.A(_07381_),
    .B(_07384_),
    .Y(_07385_));
 BUFx4f_ASAP7_75t_R _14387_ (.A(_07385_),
    .Y(_07386_));
 OR2x2_ASAP7_75t_R _14388_ (.A(_00367_),
    .B(_00400_),
    .Y(_07387_));
 BUFx3_ASAP7_75t_R _14389_ (.A(_07387_),
    .Y(_07388_));
 INVx1_ASAP7_75t_R _14390_ (.A(_07388_),
    .Y(_07389_));
 AND3x1_ASAP7_75t_R _14391_ (.A(_00334_),
    .B(_07386_),
    .C(_07389_),
    .Y(_07390_));
 INVx1_ASAP7_75t_R _14392_ (.A(_00334_),
    .Y(_07391_));
 NOR2x1_ASAP7_75t_R _14393_ (.A(_03528_),
    .B(_03534_),
    .Y(_07392_));
 AND5x2_ASAP7_75t_R _14394_ (.A(_06806_),
    .B(_03559_),
    .C(_03532_),
    .D(_07392_),
    .E(_05755_),
    .Y(_07393_));
 OA21x2_ASAP7_75t_R _14395_ (.A1(_00565_),
    .A2(_00598_),
    .B(_01189_),
    .Y(_07394_));
 OA21x2_ASAP7_75t_R _14396_ (.A1(_00532_),
    .A2(_07394_),
    .B(_01187_),
    .Y(_07395_));
 OA21x2_ASAP7_75t_R _14397_ (.A1(_00499_),
    .A2(_07395_),
    .B(_01185_),
    .Y(_07396_));
 OA21x2_ASAP7_75t_R _14398_ (.A1(_00466_),
    .A2(_07396_),
    .B(_01183_),
    .Y(_07397_));
 OA21x2_ASAP7_75t_R _14399_ (.A1(_00433_),
    .A2(_07397_),
    .B(_01181_),
    .Y(_07398_));
 OA21x2_ASAP7_75t_R _14400_ (.A1(_00400_),
    .A2(_07398_),
    .B(_01180_),
    .Y(_07399_));
 OA21x2_ASAP7_75t_R _14401_ (.A1(_00367_),
    .A2(_07399_),
    .B(_01178_),
    .Y(_07400_));
 AND3x1_ASAP7_75t_R _14402_ (.A(_07391_),
    .B(_07385_),
    .C(_07388_),
    .Y(_07401_));
 INVx1_ASAP7_75t_R _14403_ (.A(_07400_),
    .Y(_07402_));
 AND3x1_ASAP7_75t_R _14404_ (.A(_00334_),
    .B(_07386_),
    .C(_07402_),
    .Y(_07403_));
 AO221x1_ASAP7_75t_R _14405_ (.A1(_07391_),
    .A2(_07393_),
    .B1(_07400_),
    .B2(_07401_),
    .C(_07403_),
    .Y(_07404_));
 AND3x1_ASAP7_75t_R _14406_ (.A(_07391_),
    .B(_07385_),
    .C(_07400_),
    .Y(_07405_));
 OA211x2_ASAP7_75t_R _14407_ (.A1(_07346_),
    .A2(_07357_),
    .B(_07405_),
    .C(_07370_),
    .Y(_07406_));
 AO211x2_ASAP7_75t_R _14408_ (.A1(_07371_),
    .A2(_07390_),
    .B(_07404_),
    .C(_07406_),
    .Y(_07407_));
 INVx3_ASAP7_75t_R _14409_ (.A(_07381_),
    .Y(_07408_));
 NOR2x2_ASAP7_75t_R _14410_ (.A(_07383_),
    .B(_07393_),
    .Y(_07409_));
 INVx1_ASAP7_75t_R _14411_ (.A(_00333_),
    .Y(_07410_));
 AO22x1_ASAP7_75t_R _14412_ (.A1(_01176_),
    .A2(_07383_),
    .B1(_07409_),
    .B2(_07410_),
    .Y(_07411_));
 AND2x6_ASAP7_75t_R _14413_ (.A(_03822_),
    .B(_07334_),
    .Y(_07412_));
 AO21x2_ASAP7_75t_R _14414_ (.A1(_07408_),
    .A2(_07411_),
    .B(_07412_),
    .Y(_07413_));
 OR2x2_ASAP7_75t_R _14415_ (.A(_07407_),
    .B(_07413_),
    .Y(_07414_));
 BUFx6f_ASAP7_75t_R _14416_ (.A(_07414_),
    .Y(_07415_));
 NAND2x2_ASAP7_75t_R _14417_ (.A(_07339_),
    .B(_07415_),
    .Y(_07416_));
 INVx5_ASAP7_75t_R _14418_ (.A(_07416_),
    .Y(_07417_));
 BUFx6f_ASAP7_75t_R _14419_ (.A(_07417_),
    .Y(net47));
 INVx1_ASAP7_75t_R _14420_ (.A(_00599_),
    .Y(_07418_));
 OA211x2_ASAP7_75t_R _14421_ (.A1(_07346_),
    .A2(_07356_),
    .B(_07364_),
    .C(_07369_),
    .Y(_07419_));
 AND3x1_ASAP7_75t_R _14422_ (.A(_07418_),
    .B(_07386_),
    .C(_07419_),
    .Y(_07420_));
 OA21x2_ASAP7_75t_R _14423_ (.A1(_07346_),
    .A2(_07356_),
    .B(_07369_),
    .Y(_07421_));
 NAND2x1_ASAP7_75t_R _14424_ (.A(_00599_),
    .B(_07386_),
    .Y(_07422_));
 BUFx4f_ASAP7_75t_R _14425_ (.A(_07381_),
    .Y(_07423_));
 OR2x6_ASAP7_75t_R _14426_ (.A(_07383_),
    .B(_07393_),
    .Y(_07424_));
 NAND2x1_ASAP7_75t_R _14427_ (.A(_01191_),
    .B(_07383_),
    .Y(_07425_));
 OA21x2_ASAP7_75t_R _14428_ (.A1(_00598_),
    .A2(_07424_),
    .B(_07425_),
    .Y(_07426_));
 NAND2x1_ASAP7_75t_R _14429_ (.A(_03559_),
    .B(_03532_),
    .Y(_07427_));
 OR5x2_ASAP7_75t_R _14430_ (.A(_03528_),
    .B(_03534_),
    .C(_03519_),
    .D(_07239_),
    .E(_07427_),
    .Y(_07428_));
 OA21x2_ASAP7_75t_R _14431_ (.A1(_00599_),
    .A2(_07428_),
    .B(_07335_),
    .Y(_07429_));
 NAND2x2_ASAP7_75t_R _14432_ (.A(_07381_),
    .B(_07384_),
    .Y(_07430_));
 OR3x1_ASAP7_75t_R _14433_ (.A(_07418_),
    .B(_07430_),
    .C(_07364_),
    .Y(_07431_));
 OA211x2_ASAP7_75t_R _14434_ (.A1(_07423_),
    .A2(_07426_),
    .B(_07429_),
    .C(_07431_),
    .Y(_07432_));
 OAI21x1_ASAP7_75t_R _14435_ (.A1(_07421_),
    .A2(_07422_),
    .B(_07432_),
    .Y(_07433_));
 AND2x2_ASAP7_75t_R _14436_ (.A(_07328_),
    .B(_06963_),
    .Y(_07434_));
 OA211x2_ASAP7_75t_R _14437_ (.A1(_07317_),
    .A2(_07322_),
    .B(_07434_),
    .C(_07276_),
    .Y(_07435_));
 OR3x1_ASAP7_75t_R _14438_ (.A(_06865_),
    .B(_06963_),
    .C(_07276_),
    .Y(_07436_));
 AO211x2_ASAP7_75t_R _14439_ (.A1(_05851_),
    .A2(_07305_),
    .B(_07436_),
    .C(_07307_),
    .Y(_07437_));
 BUFx6f_ASAP7_75t_R _14440_ (.A(_07298_),
    .Y(_07438_));
 AO32x1_ASAP7_75t_R _14441_ (.A1(_07238_),
    .A2(_07438_),
    .A3(_07290_),
    .B1(_07276_),
    .B2(_04169_),
    .Y(_07439_));
 AND3x1_ASAP7_75t_R _14442_ (.A(_03911_),
    .B(_06865_),
    .C(_07276_),
    .Y(_07440_));
 AOI21x1_ASAP7_75t_R _14443_ (.A1(_07439_),
    .A2(_07440_),
    .B(_07335_),
    .Y(_07441_));
 OAI21x1_ASAP7_75t_R _14444_ (.A1(_07304_),
    .A2(_07437_),
    .B(_07441_),
    .Y(_07442_));
 AND3x1_ASAP7_75t_R _14445_ (.A(_07328_),
    .B(_06963_),
    .C(_07243_),
    .Y(_07443_));
 INVx1_ASAP7_75t_R _14446_ (.A(_07443_),
    .Y(_07444_));
 NOR3x1_ASAP7_75t_R _14447_ (.A(_07260_),
    .B(_07272_),
    .C(_07444_),
    .Y(_07445_));
 NAND2x2_ASAP7_75t_R _14448_ (.A(_10002_),
    .B(_07184_),
    .Y(_07446_));
 OA211x2_ASAP7_75t_R _14449_ (.A1(_10012_),
    .A2(_07184_),
    .B(_07249_),
    .C(_07446_),
    .Y(_07447_));
 OA21x2_ASAP7_75t_R _14450_ (.A1(_05529_),
    .A2(_05545_),
    .B(_07184_),
    .Y(_07448_));
 AND2x4_ASAP7_75t_R _14451_ (.A(_10029_),
    .B(_07270_),
    .Y(_07449_));
 NOR3x2_ASAP7_75t_R _14452_ (.B(_07448_),
    .C(_07449_),
    .Y(_07450_),
    .A(_07306_));
 AOI21x1_ASAP7_75t_R _14453_ (.A1(_07251_),
    .A2(_07182_),
    .B(_05345_),
    .Y(_07451_));
 AOI21x1_ASAP7_75t_R _14454_ (.A1(_03792_),
    .A2(_05308_),
    .B(_03809_),
    .Y(_07452_));
 OAI21x1_ASAP7_75t_R _14455_ (.A1(_05312_),
    .A2(_05313_),
    .B(_04915_),
    .Y(_07453_));
 AO221x1_ASAP7_75t_R _14456_ (.A1(_05319_),
    .A2(_05320_),
    .B1(_05322_),
    .B2(_05323_),
    .C(_05235_),
    .Y(_07454_));
 NOR2x1_ASAP7_75t_R _14457_ (.A(_04452_),
    .B(_05329_),
    .Y(_07455_));
 NAND2x1_ASAP7_75t_R _14458_ (.A(_05337_),
    .B(_05340_),
    .Y(_07456_));
 AO32x2_ASAP7_75t_R _14459_ (.A1(_07452_),
    .A2(_07453_),
    .A3(_07454_),
    .B1(_07455_),
    .B2(_07456_),
    .Y(_07457_));
 AO32x2_ASAP7_75t_R _14460_ (.A1(_09999_),
    .A2(_07251_),
    .A3(_07182_),
    .B1(_07451_),
    .B2(_07457_),
    .Y(_07458_));
 OA22x2_ASAP7_75t_R _14461_ (.A1(_05850_),
    .A2(_05825_),
    .B1(_07254_),
    .B2(_07255_),
    .Y(_07459_));
 AOI22x1_ASAP7_75t_R _14462_ (.A1(_10024_),
    .A2(_07184_),
    .B1(_07459_),
    .B2(_05845_),
    .Y(_07460_));
 AO32x2_ASAP7_75t_R _14463_ (.A1(_07235_),
    .A2(_07077_),
    .A3(_07458_),
    .B1(_07460_),
    .B2(_07259_),
    .Y(_07461_));
 AND3x1_ASAP7_75t_R _14464_ (.A(_07328_),
    .B(_07238_),
    .C(_07276_),
    .Y(_07462_));
 OA31x2_ASAP7_75t_R _14465_ (.A1(_07447_),
    .A2(_07450_),
    .A3(_07461_),
    .B1(_07462_),
    .Y(_07463_));
 OR4x2_ASAP7_75t_R _14466_ (.A(_07435_),
    .B(_07442_),
    .C(_07445_),
    .D(_07463_),
    .Y(_07464_));
 OAI21x1_ASAP7_75t_R _14467_ (.A1(_07420_),
    .A2(_07433_),
    .B(_07464_),
    .Y(_07465_));
 CKINVDCx6p67_ASAP7_75t_R _14468_ (.A(_07465_),
    .Y(net38));
 INVx1_ASAP7_75t_R _14469_ (.A(_01163_),
    .Y(_07466_));
 INVx1_ASAP7_75t_R _14470_ (.A(_01162_),
    .Y(_07467_));
 AO22x1_ASAP7_75t_R _14471_ (.A1(_01164_),
    .A2(_07383_),
    .B1(_07409_),
    .B2(_07467_),
    .Y(_07468_));
 AOI221x1_ASAP7_75t_R _14472_ (.A1(_07466_),
    .A2(_07393_),
    .B1(_07468_),
    .B2(_07408_),
    .C(_07412_),
    .Y(_07469_));
 OR2x2_ASAP7_75t_R _14473_ (.A(_00300_),
    .B(_00334_),
    .Y(_07470_));
 OR3x1_ASAP7_75t_R _14474_ (.A(_00234_),
    .B(_00267_),
    .C(_07470_),
    .Y(_07471_));
 OR5x2_ASAP7_75t_R _14475_ (.A(_00100_),
    .B(_00134_),
    .C(_00167_),
    .D(_00201_),
    .E(_07471_),
    .Y(_07472_));
 NOR2x1_ASAP7_75t_R _14476_ (.A(_07388_),
    .B(_07472_),
    .Y(_07473_));
 OA21x2_ASAP7_75t_R _14477_ (.A1(_00300_),
    .A2(_00333_),
    .B(_01174_),
    .Y(_07474_));
 OA21x2_ASAP7_75t_R _14478_ (.A1(_00267_),
    .A2(_07474_),
    .B(_01173_),
    .Y(_07475_));
 OA21x2_ASAP7_75t_R _14479_ (.A1(_00234_),
    .A2(_07475_),
    .B(_01171_),
    .Y(_07476_));
 OA21x2_ASAP7_75t_R _14480_ (.A1(_00201_),
    .A2(_07476_),
    .B(_00200_),
    .Y(_07477_));
 OA21x2_ASAP7_75t_R _14481_ (.A1(_00167_),
    .A2(_07477_),
    .B(_01168_),
    .Y(_07478_));
 OA21x2_ASAP7_75t_R _14482_ (.A1(_00134_),
    .A2(_07478_),
    .B(_00133_),
    .Y(_07479_));
 OA21x2_ASAP7_75t_R _14483_ (.A1(_00100_),
    .A2(_07479_),
    .B(_00099_),
    .Y(_07480_));
 OAI21x1_ASAP7_75t_R _14484_ (.A1(_07400_),
    .A2(_07472_),
    .B(_07480_),
    .Y(_07481_));
 AOI21x1_ASAP7_75t_R _14485_ (.A1(_07371_),
    .A2(_07473_),
    .B(_07481_),
    .Y(_07482_));
 OR3x1_ASAP7_75t_R _14486_ (.A(_07466_),
    .B(_07430_),
    .C(_07482_),
    .Y(_07483_));
 AO21x1_ASAP7_75t_R _14487_ (.A1(_07371_),
    .A2(_07473_),
    .B(_07481_),
    .Y(_07484_));
 OR3x1_ASAP7_75t_R _14488_ (.A(_01163_),
    .B(_07430_),
    .C(_07484_),
    .Y(_07485_));
 AOI221x1_ASAP7_75t_R _14489_ (.A1(_10019_),
    .A2(_07288_),
    .B1(_07292_),
    .B2(_07078_),
    .C(_07284_),
    .Y(_07486_));
 NAND2x2_ASAP7_75t_R _14490_ (.A(_06866_),
    .B(_07243_),
    .Y(_07487_));
 INVx1_ASAP7_75t_R _14491_ (.A(_07487_),
    .Y(_07488_));
 BUFx6f_ASAP7_75t_R _14492_ (.A(_07238_),
    .Y(_07489_));
 AO21x1_ASAP7_75t_R _14493_ (.A1(_05851_),
    .A2(_07305_),
    .B(_07307_),
    .Y(_07490_));
 OR2x2_ASAP7_75t_R _14494_ (.A(_06963_),
    .B(_07490_),
    .Y(_07491_));
 OAI22x1_ASAP7_75t_R _14495_ (.A1(_07489_),
    .A2(_07273_),
    .B1(_07304_),
    .B2(_07491_),
    .Y(_07492_));
 AND2x2_ASAP7_75t_R _14496_ (.A(_07247_),
    .B(_07248_),
    .Y(_07493_));
 AND3x1_ASAP7_75t_R _14497_ (.A(_04809_),
    .B(_04847_),
    .C(_07184_),
    .Y(_07494_));
 OR2x2_ASAP7_75t_R _14498_ (.A(_07313_),
    .B(_07494_),
    .Y(_07495_));
 NAND2x1_ASAP7_75t_R _14499_ (.A(_09977_),
    .B(_07270_),
    .Y(_07496_));
 OA21x2_ASAP7_75t_R _14500_ (.A1(_09987_),
    .A2(_07270_),
    .B(_07496_),
    .Y(_07497_));
 OA22x2_ASAP7_75t_R _14501_ (.A1(_07493_),
    .A2(_07495_),
    .B1(_07497_),
    .B2(_07268_),
    .Y(_07498_));
 INVx1_ASAP7_75t_R _14502_ (.A(_07259_),
    .Y(_07499_));
 BUFx6f_ASAP7_75t_R _14503_ (.A(_07184_),
    .Y(_07500_));
 NAND2x1_ASAP7_75t_R _14504_ (.A(_09962_),
    .B(_07184_),
    .Y(_07501_));
 OA21x2_ASAP7_75t_R _14505_ (.A1(_03911_),
    .A2(_07500_),
    .B(_07501_),
    .Y(_07502_));
 OR2x2_ASAP7_75t_R _14506_ (.A(_09969_),
    .B(_07270_),
    .Y(_07503_));
 NAND2x1_ASAP7_75t_R _14507_ (.A(_09957_),
    .B(_07270_),
    .Y(_07504_));
 AO21x1_ASAP7_75t_R _14508_ (.A1(_07503_),
    .A2(_07504_),
    .B(_07306_),
    .Y(_07505_));
 BUFx6f_ASAP7_75t_R _14509_ (.A(_07328_),
    .Y(_07506_));
 AND3x2_ASAP7_75t_R _14510_ (.A(_07506_),
    .B(_07238_),
    .C(_07243_),
    .Y(_07507_));
 OA211x2_ASAP7_75t_R _14511_ (.A1(_07499_),
    .A2(_07502_),
    .B(_07505_),
    .C(_07507_),
    .Y(_07508_));
 AND3x2_ASAP7_75t_R _14512_ (.A(_07328_),
    .B(_07238_),
    .C(_07311_),
    .Y(_07509_));
 AO21x1_ASAP7_75t_R _14513_ (.A1(_07305_),
    .A2(_07509_),
    .B(_07277_),
    .Y(_07510_));
 AO21x1_ASAP7_75t_R _14514_ (.A1(_03911_),
    .A2(_07510_),
    .B(_07336_),
    .Y(_07511_));
 AO21x1_ASAP7_75t_R _14515_ (.A1(_07498_),
    .A2(_07508_),
    .B(_07511_),
    .Y(_07512_));
 AOI221x1_ASAP7_75t_R _14516_ (.A1(_07486_),
    .A2(_07443_),
    .B1(_07488_),
    .B2(_07492_),
    .C(_07512_),
    .Y(_07513_));
 AO31x2_ASAP7_75t_R _14517_ (.A1(_07469_),
    .A2(_07483_),
    .A3(_07485_),
    .B(_07513_),
    .Y(_07514_));
 CKINVDCx5p33_ASAP7_75t_R _14518_ (.A(_07514_),
    .Y(_07515_));
 BUFx10_ASAP7_75t_R _14519_ (.A(_07515_),
    .Y(\dmem.ce_mem[3] ));
 BUFx4f_ASAP7_75t_R _14520_ (.A(_07276_),
    .Y(_07516_));
 BUFx6f_ASAP7_75t_R _14521_ (.A(_07516_),
    .Y(_07517_));
 BUFx6f_ASAP7_75t_R _14522_ (.A(_07270_),
    .Y(_07518_));
 OR3x2_ASAP7_75t_R _14523_ (.A(_06290_),
    .B(_06331_),
    .C(_07518_),
    .Y(_07519_));
 OA21x2_ASAP7_75t_R _14524_ (.A1(_10064_),
    .A2(_07186_),
    .B(_07519_),
    .Y(_07520_));
 BUFx4f_ASAP7_75t_R _14525_ (.A(_07235_),
    .Y(_07521_));
 BUFx6f_ASAP7_75t_R _14526_ (.A(_07270_),
    .Y(_07522_));
 OR3x2_ASAP7_75t_R _14527_ (.A(_06207_),
    .B(_06238_),
    .C(_07522_),
    .Y(_07523_));
 OR2x2_ASAP7_75t_R _14528_ (.A(_10059_),
    .B(_07185_),
    .Y(_07524_));
 AND3x1_ASAP7_75t_R _14529_ (.A(_07521_),
    .B(_07523_),
    .C(_07524_),
    .Y(_07525_));
 AO21x1_ASAP7_75t_R _14530_ (.A1(_03581_),
    .A2(_07520_),
    .B(_07525_),
    .Y(_07526_));
 NOR2x2_ASAP7_75t_R _14531_ (.A(_10037_),
    .B(_07522_),
    .Y(_07527_));
 AND2x2_ASAP7_75t_R _14532_ (.A(_10049_),
    .B(_07522_),
    .Y(_07528_));
 OR3x1_ASAP7_75t_R _14533_ (.A(_07521_),
    .B(_07527_),
    .C(_07528_),
    .Y(_07529_));
 BUFx6f_ASAP7_75t_R _14534_ (.A(_07500_),
    .Y(_07530_));
 NOR2x1_ASAP7_75t_R _14535_ (.A(_10042_),
    .B(_07530_),
    .Y(_07531_));
 AO221x1_ASAP7_75t_R _14536_ (.A1(_03576_),
    .A2(_03577_),
    .B1(_10034_),
    .B2(_07186_),
    .C(_07531_),
    .Y(_07532_));
 BUFx6f_ASAP7_75t_R _14537_ (.A(_07438_),
    .Y(_07533_));
 BUFx6f_ASAP7_75t_R _14538_ (.A(_07533_),
    .Y(_07534_));
 BUFx6f_ASAP7_75t_R _14539_ (.A(_07534_),
    .Y(_07535_));
 AO21x1_ASAP7_75t_R _14540_ (.A1(_07529_),
    .A2(_07532_),
    .B(_07535_),
    .Y(_07536_));
 OAI21x1_ASAP7_75t_R _14541_ (.A1(_07081_),
    .A2(_07526_),
    .B(_07536_),
    .Y(_07537_));
 BUFx4f_ASAP7_75t_R _14542_ (.A(_06964_),
    .Y(_07538_));
 BUFx6f_ASAP7_75t_R _14543_ (.A(_07533_),
    .Y(_07539_));
 BUFx4f_ASAP7_75t_R _14544_ (.A(_07539_),
    .Y(_07540_));
 BUFx4f_ASAP7_75t_R _14545_ (.A(_03579_),
    .Y(_07541_));
 AO211x2_ASAP7_75t_R _14546_ (.A1(_04601_),
    .A2(_04621_),
    .B(_04630_),
    .C(_07522_),
    .Y(_07542_));
 NAND3x1_ASAP7_75t_R _14547_ (.A(_04809_),
    .B(_04847_),
    .C(_07518_),
    .Y(_07543_));
 NAND2x1_ASAP7_75t_R _14548_ (.A(_07542_),
    .B(_07543_),
    .Y(_07544_));
 BUFx4f_ASAP7_75t_R _14549_ (.A(_07235_),
    .Y(_07545_));
 OR2x2_ASAP7_75t_R _14550_ (.A(_07545_),
    .B(_07321_),
    .Y(_07546_));
 OA21x2_ASAP7_75t_R _14551_ (.A1(_07541_),
    .A2(_07544_),
    .B(_07546_),
    .Y(_07547_));
 BUFx4f_ASAP7_75t_R _14552_ (.A(_07235_),
    .Y(_07548_));
 BUFx4f_ASAP7_75t_R _14553_ (.A(_07270_),
    .Y(_07549_));
 BUFx4f_ASAP7_75t_R _14554_ (.A(_07549_),
    .Y(_07550_));
 NAND2x1_ASAP7_75t_R _14555_ (.A(_09962_),
    .B(_07550_),
    .Y(_07551_));
 BUFx6f_ASAP7_75t_R _14556_ (.A(_07500_),
    .Y(_07552_));
 NAND2x1_ASAP7_75t_R _14557_ (.A(_09955_),
    .B(_07552_),
    .Y(_07553_));
 AO222x2_ASAP7_75t_R _14558_ (.A1(_04453_),
    .A2(_04469_),
    .B1(_04484_),
    .B2(_04500_),
    .C1(_07251_),
    .C2(_07182_),
    .Y(_07554_));
 OA211x2_ASAP7_75t_R _14559_ (.A1(_09959_),
    .A2(_07518_),
    .B(_07554_),
    .C(_03579_),
    .Y(_07555_));
 AO31x2_ASAP7_75t_R _14560_ (.A1(_07548_),
    .A2(_07551_),
    .A3(_07553_),
    .B(_07555_),
    .Y(_07556_));
 AND2x2_ASAP7_75t_R _14561_ (.A(_07080_),
    .B(_07556_),
    .Y(_07557_));
 AOI21x1_ASAP7_75t_R _14562_ (.A1(_07540_),
    .A2(_07547_),
    .B(_07557_),
    .Y(_07558_));
 BUFx4f_ASAP7_75t_R _14563_ (.A(_07489_),
    .Y(_07559_));
 OR3x1_ASAP7_75t_R _14564_ (.A(_07548_),
    .B(_07448_),
    .C(_07449_),
    .Y(_07560_));
 AND3x1_ASAP7_75t_R _14565_ (.A(_05424_),
    .B(_05446_),
    .C(_07185_),
    .Y(_07561_));
 AND2x2_ASAP7_75t_R _14566_ (.A(_10024_),
    .B(_07522_),
    .Y(_07562_));
 OR3x1_ASAP7_75t_R _14567_ (.A(_03580_),
    .B(_07561_),
    .C(_07562_),
    .Y(_07563_));
 AO222x2_ASAP7_75t_R _14568_ (.A1(_05220_),
    .A2(_05236_),
    .B1(_05247_),
    .B2(_05256_),
    .C1(_07251_),
    .C2(_07182_),
    .Y(_07564_));
 OA211x2_ASAP7_75t_R _14569_ (.A1(_09992_),
    .A2(_07549_),
    .B(_07564_),
    .C(_07235_),
    .Y(_07565_));
 AOI211x1_ASAP7_75t_R _14570_ (.A1(_07541_),
    .A2(_07458_),
    .B(_07565_),
    .C(_07533_),
    .Y(_07566_));
 AO31x2_ASAP7_75t_R _14571_ (.A1(_07539_),
    .A2(_07560_),
    .A3(_07563_),
    .B(_07566_),
    .Y(_07567_));
 AND2x2_ASAP7_75t_R _14572_ (.A(_07559_),
    .B(_07567_),
    .Y(_07568_));
 AOI21x1_ASAP7_75t_R _14573_ (.A1(_07538_),
    .A2(_07558_),
    .B(_07568_),
    .Y(_07569_));
 BUFx6f_ASAP7_75t_R _14574_ (.A(_07545_),
    .Y(_07570_));
 NAND2x1_ASAP7_75t_R _14575_ (.A(_10069_),
    .B(_07185_),
    .Y(_07571_));
 AO222x2_ASAP7_75t_R _14576_ (.A1(_06774_),
    .A2(_06784_),
    .B1(_06794_),
    .B2(_06804_),
    .C1(_07251_),
    .C2(_07182_),
    .Y(_07572_));
 AND2x2_ASAP7_75t_R _14577_ (.A(_07571_),
    .B(_07572_),
    .Y(_07573_));
 NAND2x2_ASAP7_75t_R _14578_ (.A(_10074_),
    .B(_07500_),
    .Y(_07574_));
 AO222x2_ASAP7_75t_R _14579_ (.A1(_06878_),
    .A2(_06888_),
    .B1(_06898_),
    .B2(_06908_),
    .C1(_07251_),
    .C2(_07182_),
    .Y(_07575_));
 AND3x1_ASAP7_75t_R _14580_ (.A(_03580_),
    .B(_07574_),
    .C(_07575_),
    .Y(_07576_));
 AO21x1_ASAP7_75t_R _14581_ (.A1(_07570_),
    .A2(_07573_),
    .B(_07576_),
    .Y(_07577_));
 BUFx4f_ASAP7_75t_R _14582_ (.A(_07079_),
    .Y(_07578_));
 BUFx6f_ASAP7_75t_R _14583_ (.A(_07548_),
    .Y(_07579_));
 BUFx4f_ASAP7_75t_R _14584_ (.A(_07522_),
    .Y(_07580_));
 AND2x2_ASAP7_75t_R _14585_ (.A(_10087_),
    .B(_07530_),
    .Y(_07581_));
 AO21x1_ASAP7_75t_R _14586_ (.A1(_07580_),
    .A2(_09941_),
    .B(_07581_),
    .Y(_07582_));
 OR2x2_ASAP7_75t_R _14587_ (.A(_10092_),
    .B(_07522_),
    .Y(_07583_));
 OA211x2_ASAP7_75t_R _14588_ (.A1(_09949_),
    .A2(_07186_),
    .B(_07583_),
    .C(_03580_),
    .Y(_07584_));
 AO21x1_ASAP7_75t_R _14589_ (.A1(_07579_),
    .A2(_07582_),
    .B(_07584_),
    .Y(_07585_));
 OR2x2_ASAP7_75t_R _14590_ (.A(_07578_),
    .B(_07585_),
    .Y(_07586_));
 OA211x2_ASAP7_75t_R _14591_ (.A1(_07535_),
    .A2(_07577_),
    .B(_07586_),
    .C(_07329_),
    .Y(_07587_));
 AO221x1_ASAP7_75t_R _14592_ (.A1(_07434_),
    .A2(_07537_),
    .B1(_07569_),
    .B2(_06867_),
    .C(_07587_),
    .Y(_07588_));
 AND2x2_ASAP7_75t_R _14593_ (.A(_07517_),
    .B(_07588_),
    .Y(_07589_));
 AND2x2_ASAP7_75t_R _14594_ (.A(_09949_),
    .B(_07305_),
    .Y(_07590_));
 BUFx6f_ASAP7_75t_R _14595_ (.A(_07336_),
    .Y(_07591_));
 BUFx6f_ASAP7_75t_R _14596_ (.A(_07591_),
    .Y(_07592_));
 AO21x1_ASAP7_75t_R _14597_ (.A1(_07507_),
    .A2(_07590_),
    .B(_07592_),
    .Y(_07593_));
 BUFx4f_ASAP7_75t_R _14598_ (.A(_07423_),
    .Y(_07594_));
 BUFx6f_ASAP7_75t_R _14599_ (.A(_07383_),
    .Y(_07595_));
 BUFx6f_ASAP7_75t_R _14600_ (.A(_07595_),
    .Y(_07596_));
 AND2x2_ASAP7_75t_R _14601_ (.A(_07594_),
    .B(_07596_),
    .Y(_07597_));
 OA21x2_ASAP7_75t_R _14602_ (.A1(_01030_),
    .A2(_01064_),
    .B(_01211_),
    .Y(_07598_));
 OA21x2_ASAP7_75t_R _14603_ (.A1(_00997_),
    .A2(_07598_),
    .B(_01209_),
    .Y(_07599_));
 OA211x2_ASAP7_75t_R _14604_ (.A1(_07353_),
    .A2(_07599_),
    .B(_07366_),
    .C(_01207_),
    .Y(_07600_));
 OR4x1_ASAP7_75t_R _14605_ (.A(_00731_),
    .B(_00830_),
    .C(_00864_),
    .D(_07351_),
    .Y(_07601_));
 AO21x1_ASAP7_75t_R _14606_ (.A1(_07366_),
    .A2(_07354_),
    .B(_07601_),
    .Y(_07602_));
 OR2x2_ASAP7_75t_R _14607_ (.A(_07600_),
    .B(_07602_),
    .Y(_07603_));
 OA211x2_ASAP7_75t_R _14608_ (.A1(_00731_),
    .A2(_07360_),
    .B(_01198_),
    .C(_01196_),
    .Y(_07604_));
 AO221x2_ASAP7_75t_R _14609_ (.A1(_00698_),
    .A2(_01196_),
    .B1(_07603_),
    .B2(_07604_),
    .C(_07350_),
    .Y(_07605_));
 OR2x2_ASAP7_75t_R _14610_ (.A(_07349_),
    .B(_07388_),
    .Y(_07606_));
 OA211x2_ASAP7_75t_R _14611_ (.A1(_00367_),
    .A2(_01180_),
    .B(_01178_),
    .C(_00333_),
    .Y(_07607_));
 OA21x2_ASAP7_75t_R _14612_ (.A1(_00599_),
    .A2(_07363_),
    .B(_00598_),
    .Y(_07608_));
 AND3x1_ASAP7_75t_R _14613_ (.A(_01185_),
    .B(_01187_),
    .C(_01189_),
    .Y(_07609_));
 OA21x2_ASAP7_75t_R _14614_ (.A1(_00565_),
    .A2(_07608_),
    .B(_07609_),
    .Y(_07610_));
 AND3x1_ASAP7_75t_R _14615_ (.A(_00532_),
    .B(_01185_),
    .C(_01187_),
    .Y(_07611_));
 AO21x1_ASAP7_75t_R _14616_ (.A1(_00499_),
    .A2(_01185_),
    .B(_07611_),
    .Y(_07612_));
 OR5x1_ASAP7_75t_R _14617_ (.A(_00433_),
    .B(_00466_),
    .C(_07388_),
    .D(_07610_),
    .E(_07612_),
    .Y(_07613_));
 OR3x1_ASAP7_75t_R _14618_ (.A(_00433_),
    .B(_01183_),
    .C(_07388_),
    .Y(_07614_));
 OA211x2_ASAP7_75t_R _14619_ (.A1(_01181_),
    .A2(_07388_),
    .B(_07613_),
    .C(_07614_),
    .Y(_07615_));
 OA211x2_ASAP7_75t_R _14620_ (.A1(_07605_),
    .A2(_07606_),
    .B(_07607_),
    .C(_07615_),
    .Y(_07616_));
 AO21x1_ASAP7_75t_R _14621_ (.A1(_00334_),
    .A2(_00333_),
    .B(_00300_),
    .Y(_07617_));
 AND3x1_ASAP7_75t_R _14622_ (.A(_01171_),
    .B(_01173_),
    .C(_01174_),
    .Y(_07618_));
 OA21x2_ASAP7_75t_R _14623_ (.A1(_07616_),
    .A2(_07617_),
    .B(_07618_),
    .Y(_07619_));
 AND3x1_ASAP7_75t_R _14624_ (.A(_00267_),
    .B(_01171_),
    .C(_01173_),
    .Y(_07620_));
 AO21x1_ASAP7_75t_R _14625_ (.A1(_00234_),
    .A2(_01171_),
    .B(_07620_),
    .Y(_07621_));
 OR3x1_ASAP7_75t_R _14626_ (.A(_00134_),
    .B(_00167_),
    .C(_00201_),
    .Y(_07622_));
 OR3x1_ASAP7_75t_R _14627_ (.A(_00134_),
    .B(_00167_),
    .C(_00200_),
    .Y(_07623_));
 OA21x2_ASAP7_75t_R _14628_ (.A1(_00134_),
    .A2(_01168_),
    .B(_07623_),
    .Y(_07624_));
 OA31x2_ASAP7_75t_R _14629_ (.A1(_07619_),
    .A2(_07621_),
    .A3(_07622_),
    .B1(_07624_),
    .Y(_07625_));
 AND2x2_ASAP7_75t_R _14630_ (.A(_00133_),
    .B(_07625_),
    .Y(_07626_));
 OA21x2_ASAP7_75t_R _14631_ (.A1(_00100_),
    .A2(_07626_),
    .B(_00099_),
    .Y(_07627_));
 OA21x2_ASAP7_75t_R _14632_ (.A1(_01163_),
    .A2(_07627_),
    .B(_01162_),
    .Y(_07628_));
 OR4x2_ASAP7_75t_R _14633_ (.A(_03483_),
    .B(_07240_),
    .C(_05852_),
    .D(_07427_),
    .Y(_07629_));
 XNOR2x1_ASAP7_75t_R _14634_ (.B(_04064_),
    .Y(_07630_),
    .A(_09955_));
 AND2x2_ASAP7_75t_R _14635_ (.A(_07629_),
    .B(_07630_),
    .Y(_07631_));
 XNOR2x2_ASAP7_75t_R _14636_ (.A(_03913_),
    .B(_07631_),
    .Y(_07632_));
 XNOR2x1_ASAP7_75t_R _14637_ (.B(_07632_),
    .Y(_07633_),
    .A(_07628_));
 BUFx4f_ASAP7_75t_R _14638_ (.A(_07408_),
    .Y(_07634_));
 BUFx4f_ASAP7_75t_R _14639_ (.A(_07409_),
    .Y(_07635_));
 INVx1_ASAP7_75t_R _14640_ (.A(_01161_),
    .Y(_07636_));
 AO22x1_ASAP7_75t_R _14641_ (.A1(_01065_),
    .A2(_07596_),
    .B1(_07635_),
    .B2(_07636_),
    .Y(_07637_));
 INVx1_ASAP7_75t_R _14642_ (.A(_00034_),
    .Y(_07638_));
 BUFx4f_ASAP7_75t_R _14643_ (.A(_07393_),
    .Y(_07639_));
 AO21x1_ASAP7_75t_R _14644_ (.A1(_03913_),
    .A2(_07386_),
    .B(_07639_),
    .Y(_07640_));
 AND2x2_ASAP7_75t_R _14645_ (.A(_00034_),
    .B(_03537_),
    .Y(_07641_));
 BUFx4f_ASAP7_75t_R _14646_ (.A(_07386_),
    .Y(_07642_));
 BUFx6f_ASAP7_75t_R _14647_ (.A(_07412_),
    .Y(_07643_));
 AO221x1_ASAP7_75t_R _14648_ (.A1(_07638_),
    .A2(_07640_),
    .B1(_07641_),
    .B2(_07642_),
    .C(_07643_),
    .Y(_07644_));
 AO21x1_ASAP7_75t_R _14649_ (.A1(_07634_),
    .A2(_07637_),
    .B(_07644_),
    .Y(_07645_));
 AO21x1_ASAP7_75t_R _14650_ (.A1(_07597_),
    .A2(_07633_),
    .B(_07645_),
    .Y(_07646_));
 OA21x2_ASAP7_75t_R _14651_ (.A1(_07589_),
    .A2(_07593_),
    .B(_07646_),
    .Y(net32));
 BUFx4f_ASAP7_75t_R _14652_ (.A(_07243_),
    .Y(_07647_));
 BUFx4f_ASAP7_75t_R _14653_ (.A(_07647_),
    .Y(_07648_));
 BUFx4f_ASAP7_75t_R _14654_ (.A(_07648_),
    .Y(_07649_));
 AND3x1_ASAP7_75t_R _14655_ (.A(_03579_),
    .B(_07190_),
    .C(_07233_),
    .Y(_07650_));
 AO32x1_ASAP7_75t_R _14656_ (.A1(_04059_),
    .A2(_07075_),
    .A3(_07179_),
    .B1(_07255_),
    .B2(_07024_),
    .Y(_07651_));
 OA21x2_ASAP7_75t_R _14657_ (.A1(_07236_),
    .A2(_07650_),
    .B(_07651_),
    .Y(_07652_));
 NAND2x1_ASAP7_75t_R _14658_ (.A(_10084_),
    .B(_07186_),
    .Y(_07653_));
 OR2x4_ASAP7_75t_R _14659_ (.A(_07128_),
    .B(_07500_),
    .Y(_07654_));
 AND3x1_ASAP7_75t_R _14660_ (.A(_07579_),
    .B(_07653_),
    .C(_07654_),
    .Y(_07655_));
 AO21x1_ASAP7_75t_R _14661_ (.A1(_03581_),
    .A2(_07582_),
    .B(_07655_),
    .Y(_07656_));
 BUFx4f_ASAP7_75t_R _14662_ (.A(_07533_),
    .Y(_07657_));
 NAND2x1_ASAP7_75t_R _14663_ (.A(_10074_),
    .B(_07550_),
    .Y(_07658_));
 NAND2x1_ASAP7_75t_R _14664_ (.A(_10064_),
    .B(_07552_),
    .Y(_07659_));
 OA211x2_ASAP7_75t_R _14665_ (.A1(_10067_),
    .A2(_07518_),
    .B(_07572_),
    .C(_03579_),
    .Y(_07660_));
 AO31x2_ASAP7_75t_R _14666_ (.A1(_07521_),
    .A2(_07658_),
    .A3(_07659_),
    .B(_07660_),
    .Y(_07661_));
 OR2x2_ASAP7_75t_R _14667_ (.A(_07657_),
    .B(_07661_),
    .Y(_07662_));
 OA211x2_ASAP7_75t_R _14668_ (.A1(_07081_),
    .A2(_07656_),
    .B(_07662_),
    .C(_07516_),
    .Y(_07663_));
 AOI21x1_ASAP7_75t_R _14669_ (.A1(_07649_),
    .A2(_07652_),
    .B(_07663_),
    .Y(_07664_));
 BUFx4f_ASAP7_75t_R _14670_ (.A(_07489_),
    .Y(_07665_));
 BUFx4f_ASAP7_75t_R _14671_ (.A(_07665_),
    .Y(_07666_));
 AND2x2_ASAP7_75t_R _14672_ (.A(_10049_),
    .B(_07185_),
    .Y(_07667_));
 AO21x1_ASAP7_75t_R _14673_ (.A1(_10102_),
    .A2(_07550_),
    .B(_07667_),
    .Y(_07668_));
 AO21x1_ASAP7_75t_R _14674_ (.A1(_07523_),
    .A2(_07524_),
    .B(_07548_),
    .Y(_07669_));
 OA21x2_ASAP7_75t_R _14675_ (.A1(_07541_),
    .A2(_07668_),
    .B(_07669_),
    .Y(_07670_));
 BUFx4f_ASAP7_75t_R _14676_ (.A(_07545_),
    .Y(_07671_));
 AO21x1_ASAP7_75t_R _14677_ (.A1(_10034_),
    .A2(_07552_),
    .B(_07531_),
    .Y(_07672_));
 BUFx4f_ASAP7_75t_R _14678_ (.A(_03579_),
    .Y(_07673_));
 AND2x2_ASAP7_75t_R _14679_ (.A(_10029_),
    .B(_07500_),
    .Y(_07674_));
 NOR2x2_ASAP7_75t_R _14680_ (.A(_10037_),
    .B(_07185_),
    .Y(_07675_));
 OR3x1_ASAP7_75t_R _14681_ (.A(_07673_),
    .B(_07674_),
    .C(_07675_),
    .Y(_07676_));
 BUFx6f_ASAP7_75t_R _14682_ (.A(_07078_),
    .Y(_07677_));
 OA211x2_ASAP7_75t_R _14683_ (.A1(_07671_),
    .A2(_07672_),
    .B(_07676_),
    .C(_07677_),
    .Y(_07678_));
 AO21x1_ASAP7_75t_R _14684_ (.A1(_07535_),
    .A2(_07670_),
    .B(_07678_),
    .Y(_07679_));
 OR3x1_ASAP7_75t_R _14685_ (.A(_07666_),
    .B(_07648_),
    .C(_07679_),
    .Y(_07680_));
 AND2x2_ASAP7_75t_R _14686_ (.A(_07506_),
    .B(_07412_),
    .Y(_07681_));
 BUFx4f_ASAP7_75t_R _14687_ (.A(_07681_),
    .Y(_07682_));
 OA211x2_ASAP7_75t_R _14688_ (.A1(_06966_),
    .A2(_07664_),
    .B(_07680_),
    .C(_07682_),
    .Y(_07683_));
 BUFx4f_ASAP7_75t_R _14689_ (.A(_07424_),
    .Y(_07684_));
 NAND2x1_ASAP7_75t_R _14690_ (.A(_01214_),
    .B(_07596_),
    .Y(_07685_));
 OA21x2_ASAP7_75t_R _14691_ (.A1(_01213_),
    .A2(_07684_),
    .B(_07685_),
    .Y(_07686_));
 BUFx4f_ASAP7_75t_R _14692_ (.A(_07430_),
    .Y(_07687_));
 BUFx4f_ASAP7_75t_R _14693_ (.A(_07428_),
    .Y(_07688_));
 OA21x2_ASAP7_75t_R _14694_ (.A1(_01063_),
    .A2(_07688_),
    .B(_07591_),
    .Y(_07689_));
 OA21x2_ASAP7_75t_R _14695_ (.A1(_01066_),
    .A2(_07687_),
    .B(_07689_),
    .Y(_07690_));
 OA21x2_ASAP7_75t_R _14696_ (.A1(_07594_),
    .A2(_07686_),
    .B(_07690_),
    .Y(_07691_));
 AND2x2_ASAP7_75t_R _14697_ (.A(_06866_),
    .B(_07412_),
    .Y(_07692_));
 OR3x1_ASAP7_75t_R _14698_ (.A(_07545_),
    .B(_07561_),
    .C(_07562_),
    .Y(_07693_));
 OA21x2_ASAP7_75t_R _14699_ (.A1(_05529_),
    .A2(_05545_),
    .B(_07522_),
    .Y(_07694_));
 AO221x1_ASAP7_75t_R _14700_ (.A1(_03576_),
    .A2(_03577_),
    .B1(_10009_),
    .B2(_07552_),
    .C(_07694_),
    .Y(_07695_));
 OAI21x1_ASAP7_75t_R _14701_ (.A1(_09992_),
    .A2(_07518_),
    .B(_07564_),
    .Y(_07696_));
 OA222x2_ASAP7_75t_R _14702_ (.A1(_05119_),
    .A2(_05131_),
    .B1(_05143_),
    .B2(_05155_),
    .C1(_07254_),
    .C2(_07255_),
    .Y(_07697_));
 AO221x1_ASAP7_75t_R _14703_ (.A1(_03576_),
    .A2(_03577_),
    .B1(_09989_),
    .B2(_07185_),
    .C(_07697_),
    .Y(_07698_));
 OA211x2_ASAP7_75t_R _14704_ (.A1(_07548_),
    .A2(_07696_),
    .B(_07698_),
    .C(_07078_),
    .Y(_07699_));
 AO31x2_ASAP7_75t_R _14705_ (.A1(_07539_),
    .A2(_07693_),
    .A3(_07695_),
    .B(_07699_),
    .Y(_07700_));
 OR2x2_ASAP7_75t_R _14706_ (.A(_06965_),
    .B(_07700_),
    .Y(_07701_));
 BUFx4f_ASAP7_75t_R _14707_ (.A(_07438_),
    .Y(_07702_));
 AO21x1_ASAP7_75t_R _14708_ (.A1(_07542_),
    .A2(_07543_),
    .B(_07545_),
    .Y(_07703_));
 AND2x2_ASAP7_75t_R _14709_ (.A(_09977_),
    .B(_07549_),
    .Y(_07704_));
 NOR2x1_ASAP7_75t_R _14710_ (.A(_09969_),
    .B(_07518_),
    .Y(_07705_));
 OR3x1_ASAP7_75t_R _14711_ (.A(_07673_),
    .B(_07704_),
    .C(_07705_),
    .Y(_07706_));
 AND2x2_ASAP7_75t_R _14712_ (.A(_07235_),
    .B(_09957_),
    .Y(_07707_));
 AO221x1_ASAP7_75t_R _14713_ (.A1(_07673_),
    .A2(_09962_),
    .B1(_07251_),
    .B2(_07182_),
    .C(_07707_),
    .Y(_07708_));
 OA21x2_ASAP7_75t_R _14714_ (.A1(_09955_),
    .A2(_07580_),
    .B(_07078_),
    .Y(_07709_));
 AO32x2_ASAP7_75t_R _14715_ (.A1(_07702_),
    .A2(_07703_),
    .A3(_07706_),
    .B1(_07708_),
    .B2(_07709_),
    .Y(_07710_));
 OR2x2_ASAP7_75t_R _14716_ (.A(_07665_),
    .B(_07710_),
    .Y(_07711_));
 NAND2x2_ASAP7_75t_R _14717_ (.A(_04169_),
    .B(_07276_),
    .Y(_07712_));
 AO21x1_ASAP7_75t_R _14718_ (.A1(_07701_),
    .A2(_07711_),
    .B(_07712_),
    .Y(_07713_));
 AND2x2_ASAP7_75t_R _14719_ (.A(_07538_),
    .B(_07311_),
    .Y(_07714_));
 OR3x4_ASAP7_75t_R _14720_ (.A(_09955_),
    .B(_07438_),
    .C(_07550_),
    .Y(_07715_));
 INVx1_ASAP7_75t_R _14721_ (.A(_07715_),
    .Y(_07716_));
 AO21x1_ASAP7_75t_R _14722_ (.A1(_07702_),
    .A2(_07544_),
    .B(_07716_),
    .Y(_07717_));
 BUFx4f_ASAP7_75t_R _14723_ (.A(_03579_),
    .Y(_07718_));
 AOI211x1_ASAP7_75t_R _14724_ (.A1(_07718_),
    .A2(_09962_),
    .B(_07552_),
    .C(_07707_),
    .Y(_07719_));
 AO32x1_ASAP7_75t_R _14725_ (.A1(_07263_),
    .A2(_07496_),
    .A3(_07503_),
    .B1(_07719_),
    .B2(_07677_),
    .Y(_07720_));
 AO21x2_ASAP7_75t_R _14726_ (.A1(_03581_),
    .A2(_07717_),
    .B(_07720_),
    .Y(_07721_));
 NAND2x1_ASAP7_75t_R _14727_ (.A(_07559_),
    .B(_07311_),
    .Y(_07722_));
 NOR2x1_ASAP7_75t_R _14728_ (.A(_07722_),
    .B(_07700_),
    .Y(_07723_));
 AOI21x1_ASAP7_75t_R _14729_ (.A1(_07714_),
    .A2(_07721_),
    .B(_07723_),
    .Y(_07724_));
 AND3x1_ASAP7_75t_R _14730_ (.A(_07692_),
    .B(_07713_),
    .C(_07724_),
    .Y(_07725_));
 OR3x4_ASAP7_75t_R _14731_ (.A(_07683_),
    .B(_07691_),
    .C(_07725_),
    .Y(_07726_));
 INVx5_ASAP7_75t_R _14732_ (.A(_07726_),
    .Y(net43));
 BUFx6f_ASAP7_75t_R _14733_ (.A(_06964_),
    .Y(_07727_));
 BUFx6f_ASAP7_75t_R _14734_ (.A(_07727_),
    .Y(_07728_));
 BUFx6f_ASAP7_75t_R _14735_ (.A(_07718_),
    .Y(_07729_));
 OR3x2_ASAP7_75t_R _14736_ (.A(_06207_),
    .B(_06238_),
    .C(_07500_),
    .Y(_07730_));
 NAND2x1_ASAP7_75t_R _14737_ (.A(_10042_),
    .B(_07552_),
    .Y(_07731_));
 AND3x1_ASAP7_75t_R _14738_ (.A(_07521_),
    .B(_07730_),
    .C(_07731_),
    .Y(_07732_));
 AO21x1_ASAP7_75t_R _14739_ (.A1(_07729_),
    .A2(_07668_),
    .B(_07732_),
    .Y(_07733_));
 AO221x1_ASAP7_75t_R _14740_ (.A1(_10024_),
    .A2(_07530_),
    .B1(_07459_),
    .B2(_05845_),
    .C(_07673_),
    .Y(_07734_));
 OA31x2_ASAP7_75t_R _14741_ (.A1(_07521_),
    .A2(_07674_),
    .A3(_07675_),
    .B1(_07734_),
    .Y(_07735_));
 OR2x2_ASAP7_75t_R _14742_ (.A(_07539_),
    .B(_07735_),
    .Y(_07736_));
 OA21x2_ASAP7_75t_R _14743_ (.A1(_07578_),
    .A2(_07733_),
    .B(_07736_),
    .Y(_07737_));
 AO21x1_ASAP7_75t_R _14744_ (.A1(_10059_),
    .A2(_07530_),
    .B(_07256_),
    .Y(_07738_));
 AND2x2_ASAP7_75t_R _14745_ (.A(_10064_),
    .B(_07185_),
    .Y(_07739_));
 OR3x1_ASAP7_75t_R _14746_ (.A(_07671_),
    .B(_07264_),
    .C(_07739_),
    .Y(_07740_));
 OA21x2_ASAP7_75t_R _14747_ (.A1(_03581_),
    .A2(_07738_),
    .B(_07740_),
    .Y(_07741_));
 NAND3x1_ASAP7_75t_R _14748_ (.A(_07729_),
    .B(_07653_),
    .C(_07654_),
    .Y(_07742_));
 NOR2x1_ASAP7_75t_R _14749_ (.A(_10087_),
    .B(_07530_),
    .Y(_07743_));
 AND2x2_ASAP7_75t_R _14750_ (.A(_10079_),
    .B(_07530_),
    .Y(_07744_));
 OR3x1_ASAP7_75t_R _14751_ (.A(_07729_),
    .B(_07743_),
    .C(_07744_),
    .Y(_07745_));
 AO21x1_ASAP7_75t_R _14752_ (.A1(_07742_),
    .A2(_07745_),
    .B(_07080_),
    .Y(_07746_));
 OA211x2_ASAP7_75t_R _14753_ (.A1(_07540_),
    .A2(_07741_),
    .B(_07746_),
    .C(_07665_),
    .Y(_07747_));
 AOI211x1_ASAP7_75t_R _14754_ (.A1(_07728_),
    .A2(_07737_),
    .B(_07747_),
    .C(_07648_),
    .Y(_07748_));
 AND2x6_ASAP7_75t_R _14755_ (.A(_07489_),
    .B(_07243_),
    .Y(_07749_));
 AO21x1_ASAP7_75t_R _14756_ (.A1(_03602_),
    .A2(_03770_),
    .B(_07518_),
    .Y(_07750_));
 AND4x1_ASAP7_75t_R _14757_ (.A(_07545_),
    .B(_07550_),
    .C(_07190_),
    .D(_07233_),
    .Y(_07751_));
 AO31x2_ASAP7_75t_R _14758_ (.A1(_07541_),
    .A2(_07654_),
    .A3(_07750_),
    .B(_07751_),
    .Y(_07752_));
 NAND3x2_ASAP7_75t_R _14759_ (.B(_07749_),
    .C(_07752_),
    .Y(_07753_),
    .A(_07535_));
 NAND2x1_ASAP7_75t_R _14760_ (.A(_07682_),
    .B(_07753_),
    .Y(_07754_));
 AND2x2_ASAP7_75t_R _14761_ (.A(_07718_),
    .B(_09957_),
    .Y(_07755_));
 AO21x1_ASAP7_75t_R _14762_ (.A1(_07671_),
    .A2(_09955_),
    .B(_07755_),
    .Y(_07756_));
 AND2x2_ASAP7_75t_R _14763_ (.A(_07078_),
    .B(_07522_),
    .Y(_07757_));
 INVx1_ASAP7_75t_R _14764_ (.A(_07757_),
    .Y(_07758_));
 AOI21x1_ASAP7_75t_R _14765_ (.A1(_09964_),
    .A2(_07530_),
    .B(_07313_),
    .Y(_07759_));
 OA21x2_ASAP7_75t_R _14766_ (.A1(_07704_),
    .A2(_07705_),
    .B(_07718_),
    .Y(_07760_));
 AO211x2_ASAP7_75t_R _14767_ (.A1(_07671_),
    .A2(_07759_),
    .B(_07760_),
    .C(_07079_),
    .Y(_07761_));
 OA211x2_ASAP7_75t_R _14768_ (.A1(_07756_),
    .A2(_07758_),
    .B(_07761_),
    .C(_06964_),
    .Y(_07762_));
 OAI21x1_ASAP7_75t_R _14769_ (.A1(_07310_),
    .A2(_07715_),
    .B(_07762_),
    .Y(_07763_));
 AND2x2_ASAP7_75t_R _14770_ (.A(_10002_),
    .B(_07185_),
    .Y(_07764_));
 AND3x2_ASAP7_75t_R _14771_ (.A(_05424_),
    .B(_05446_),
    .C(_07549_),
    .Y(_07765_));
 OR2x2_ASAP7_75t_R _14772_ (.A(_07764_),
    .B(_07765_),
    .Y(_07766_));
 OR3x1_ASAP7_75t_R _14773_ (.A(_05342_),
    .B(_05345_),
    .C(_07549_),
    .Y(_07767_));
 OA211x2_ASAP7_75t_R _14774_ (.A1(_10019_),
    .A2(_07552_),
    .B(_07767_),
    .C(_07673_),
    .Y(_07768_));
 AO21x1_ASAP7_75t_R _14775_ (.A1(_07671_),
    .A2(_07766_),
    .B(_07768_),
    .Y(_07769_));
 AND3x1_ASAP7_75t_R _14776_ (.A(_07545_),
    .B(_07318_),
    .C(_07319_),
    .Y(_07770_));
 AOI211x1_ASAP7_75t_R _14777_ (.A1(_09989_),
    .A2(_07186_),
    .B(_07697_),
    .C(_07521_),
    .Y(_07771_));
 OAI21x1_ASAP7_75t_R _14778_ (.A1(_07770_),
    .A2(_07771_),
    .B(_07677_),
    .Y(_07772_));
 OA211x2_ASAP7_75t_R _14779_ (.A1(_07080_),
    .A2(_07769_),
    .B(_07772_),
    .C(_07489_),
    .Y(_07773_));
 NOR2x1_ASAP7_75t_R _14780_ (.A(_07647_),
    .B(_07773_),
    .Y(_07774_));
 NAND2x2_ASAP7_75t_R _14781_ (.A(_06866_),
    .B(_07412_),
    .Y(_07775_));
 AO21x1_ASAP7_75t_R _14782_ (.A1(_07763_),
    .A2(_07774_),
    .B(_07775_),
    .Y(_07776_));
 BUFx6f_ASAP7_75t_R _14783_ (.A(_07383_),
    .Y(_07777_));
 INVx1_ASAP7_75t_R _14784_ (.A(_01211_),
    .Y(_07778_));
 AO22x1_ASAP7_75t_R _14785_ (.A1(_01212_),
    .A2(_07777_),
    .B1(_07635_),
    .B2(_07778_),
    .Y(_07779_));
 AO21x1_ASAP7_75t_R _14786_ (.A1(_01064_),
    .A2(_07386_),
    .B(_07639_),
    .Y(_07780_));
 OAI21x1_ASAP7_75t_R _14787_ (.A1(_01064_),
    .A2(_07430_),
    .B(_01030_),
    .Y(_07781_));
 OA21x2_ASAP7_75t_R _14788_ (.A1(_01030_),
    .A2(_07780_),
    .B(_07781_),
    .Y(_07782_));
 AOI211x1_ASAP7_75t_R _14789_ (.A1(_07634_),
    .A2(_07779_),
    .B(_07782_),
    .C(_07643_),
    .Y(_07783_));
 INVx1_ASAP7_75t_R _14790_ (.A(_07783_),
    .Y(_07784_));
 OA211x2_ASAP7_75t_R _14791_ (.A1(_07748_),
    .A2(_07754_),
    .B(_07776_),
    .C(_07784_),
    .Y(_07785_));
 BUFx6f_ASAP7_75t_R _14792_ (.A(_07785_),
    .Y(net54));
 NAND2x2_ASAP7_75t_R _14793_ (.A(_07506_),
    .B(_07643_),
    .Y(_07786_));
 AO21x1_ASAP7_75t_R _14794_ (.A1(_07730_),
    .A2(_07731_),
    .B(_07521_),
    .Y(_07787_));
 OR3x1_ASAP7_75t_R _14795_ (.A(_03580_),
    .B(_07527_),
    .C(_07528_),
    .Y(_07788_));
 AND2x2_ASAP7_75t_R _14796_ (.A(_07787_),
    .B(_07788_),
    .Y(_07789_));
 AND2x2_ASAP7_75t_R _14797_ (.A(_10024_),
    .B(_07500_),
    .Y(_07790_));
 AO21x1_ASAP7_75t_R _14798_ (.A1(_10034_),
    .A2(_07580_),
    .B(_07790_),
    .Y(_07791_));
 OR3x1_ASAP7_75t_R _14799_ (.A(_07718_),
    .B(_07448_),
    .C(_07449_),
    .Y(_07792_));
 OA211x2_ASAP7_75t_R _14800_ (.A1(_07570_),
    .A2(_07791_),
    .B(_07792_),
    .C(_07677_),
    .Y(_07793_));
 AOI21x1_ASAP7_75t_R _14801_ (.A1(_07657_),
    .A2(_07789_),
    .B(_07793_),
    .Y(_07794_));
 AND2x2_ASAP7_75t_R _14802_ (.A(_03580_),
    .B(_07738_),
    .Y(_07795_));
 AO21x1_ASAP7_75t_R _14803_ (.A1(_07579_),
    .A2(_07520_),
    .B(_07795_),
    .Y(_07796_));
 NAND2x1_ASAP7_75t_R _14804_ (.A(_07574_),
    .B(_07575_),
    .Y(_07797_));
 OR3x1_ASAP7_75t_R _14805_ (.A(_07548_),
    .B(_07743_),
    .C(_07744_),
    .Y(_07798_));
 OA211x2_ASAP7_75t_R _14806_ (.A1(_07729_),
    .A2(_07797_),
    .B(_07798_),
    .C(_07702_),
    .Y(_07799_));
 AOI211x1_ASAP7_75t_R _14807_ (.A1(_07578_),
    .A2(_07796_),
    .B(_07799_),
    .C(_07727_),
    .Y(_07800_));
 AO21x1_ASAP7_75t_R _14808_ (.A1(_06965_),
    .A2(_07794_),
    .B(_07800_),
    .Y(_07801_));
 NAND2x1_ASAP7_75t_R _14809_ (.A(_07654_),
    .B(_07750_),
    .Y(_07802_));
 AND2x2_ASAP7_75t_R _14810_ (.A(_07673_),
    .B(_07253_),
    .Y(_07803_));
 AOI22x1_ASAP7_75t_R _14811_ (.A1(_07579_),
    .A2(_07802_),
    .B1(_07803_),
    .B2(_07250_),
    .Y(_07804_));
 AND3x1_ASAP7_75t_R _14812_ (.A(_07540_),
    .B(_07749_),
    .C(_07804_),
    .Y(_07805_));
 AO21x1_ASAP7_75t_R _14813_ (.A1(_07516_),
    .A2(_07801_),
    .B(_07805_),
    .Y(_07806_));
 OAI21x1_ASAP7_75t_R _14814_ (.A1(_07764_),
    .A2(_07765_),
    .B(_07533_),
    .Y(_07807_));
 AO21x1_ASAP7_75t_R _14815_ (.A1(_07318_),
    .A2(_07319_),
    .B(_07533_),
    .Y(_07808_));
 AO221x1_ASAP7_75t_R _14816_ (.A1(_09999_),
    .A2(_07500_),
    .B1(_07451_),
    .B2(_07457_),
    .C(_07077_),
    .Y(_07809_));
 OA211x2_ASAP7_75t_R _14817_ (.A1(_07438_),
    .A2(_07321_),
    .B(_07809_),
    .C(_07545_),
    .Y(_07810_));
 AO31x2_ASAP7_75t_R _14818_ (.A1(_07729_),
    .A2(_07807_),
    .A3(_07808_),
    .B(_07810_),
    .Y(_07811_));
 OA21x2_ASAP7_75t_R _14819_ (.A1(_09959_),
    .A2(_07549_),
    .B(_07554_),
    .Y(_07812_));
 OAI21x1_ASAP7_75t_R _14820_ (.A1(_07673_),
    .A2(_07812_),
    .B(_07438_),
    .Y(_07813_));
 AOI21x1_ASAP7_75t_R _14821_ (.A1(_07718_),
    .A2(_07759_),
    .B(_07813_),
    .Y(_07814_));
 AND2x2_ASAP7_75t_R _14822_ (.A(_03911_),
    .B(_07077_),
    .Y(_07815_));
 OA21x2_ASAP7_75t_R _14823_ (.A1(_07277_),
    .A2(_07290_),
    .B(_07815_),
    .Y(_07816_));
 OR3x1_ASAP7_75t_R _14824_ (.A(_07489_),
    .B(_07814_),
    .C(_07816_),
    .Y(_07817_));
 OA211x2_ASAP7_75t_R _14825_ (.A1(_06964_),
    .A2(_07811_),
    .B(_07817_),
    .C(_07516_),
    .Y(_07818_));
 OR2x2_ASAP7_75t_R _14826_ (.A(_07775_),
    .B(_07818_),
    .Y(_07819_));
 AO21x1_ASAP7_75t_R _14827_ (.A1(_09940_),
    .A2(_07341_),
    .B(_07344_),
    .Y(_07820_));
 XNOR2x1_ASAP7_75t_R _14828_ (.B(_07820_),
    .Y(_07821_),
    .A(_07340_));
 NAND2x1_ASAP7_75t_R _14829_ (.A(_01210_),
    .B(_07595_),
    .Y(_07822_));
 OA21x2_ASAP7_75t_R _14830_ (.A1(_01209_),
    .A2(_07424_),
    .B(_07822_),
    .Y(_07823_));
 OA222x2_ASAP7_75t_R _14831_ (.A1(_00997_),
    .A2(_07428_),
    .B1(_07430_),
    .B2(_07821_),
    .C1(_07823_),
    .C2(_07423_),
    .Y(_07824_));
 NAND2x1_ASAP7_75t_R _14832_ (.A(_07591_),
    .B(_07824_),
    .Y(_07825_));
 OA211x2_ASAP7_75t_R _14833_ (.A1(_07786_),
    .A2(_07806_),
    .B(_07819_),
    .C(_07825_),
    .Y(_07826_));
 BUFx4f_ASAP7_75t_R _14834_ (.A(_07826_),
    .Y(net57));
 BUFx6f_ASAP7_75t_R _14835_ (.A(_07386_),
    .Y(_07827_));
 BUFx6f_ASAP7_75t_R _14836_ (.A(_07639_),
    .Y(_07828_));
 AOI211x1_ASAP7_75t_R _14837_ (.A1(_07827_),
    .A2(_07599_),
    .B(_07353_),
    .C(_07828_),
    .Y(_07829_));
 BUFx4f_ASAP7_75t_R _14838_ (.A(_07430_),
    .Y(_07830_));
 OA21x2_ASAP7_75t_R _14839_ (.A1(_07830_),
    .A2(_07599_),
    .B(_07353_),
    .Y(_07831_));
 INVx1_ASAP7_75t_R _14840_ (.A(_01207_),
    .Y(_07832_));
 AOI22x1_ASAP7_75t_R _14841_ (.A1(_01208_),
    .A2(_07777_),
    .B1(_07635_),
    .B2(_07832_),
    .Y(_07833_));
 OA21x2_ASAP7_75t_R _14842_ (.A1(_07594_),
    .A2(_07833_),
    .B(_07591_),
    .Y(_07834_));
 OAI21x1_ASAP7_75t_R _14843_ (.A1(_07829_),
    .A2(_07831_),
    .B(_07834_),
    .Y(_07835_));
 AO21x1_ASAP7_75t_R _14844_ (.A1(_07718_),
    .A2(_07458_),
    .B(_07565_),
    .Y(_07836_));
 OR2x2_ASAP7_75t_R _14845_ (.A(_07079_),
    .B(_07836_),
    .Y(_07837_));
 OA211x2_ASAP7_75t_R _14846_ (.A1(_07657_),
    .A2(_07547_),
    .B(_07837_),
    .C(_07489_),
    .Y(_07838_));
 AND3x1_ASAP7_75t_R _14847_ (.A(_07727_),
    .B(_07657_),
    .C(_07556_),
    .Y(_07839_));
 OA21x2_ASAP7_75t_R _14848_ (.A1(_07838_),
    .A2(_07839_),
    .B(_07311_),
    .Y(_07840_));
 AO21x1_ASAP7_75t_R _14849_ (.A1(_07539_),
    .A2(_07556_),
    .B(_07815_),
    .Y(_07841_));
 AND2x2_ASAP7_75t_R _14850_ (.A(_07727_),
    .B(_07841_),
    .Y(_07842_));
 OA21x2_ASAP7_75t_R _14851_ (.A1(_07838_),
    .A2(_07842_),
    .B(_07277_),
    .Y(_07843_));
 OR3x1_ASAP7_75t_R _14852_ (.A(_07775_),
    .B(_07840_),
    .C(_07843_),
    .Y(_07844_));
 AOI211x1_ASAP7_75t_R _14853_ (.A1(_03581_),
    .A2(_07520_),
    .B(_07525_),
    .C(_07534_),
    .Y(_07845_));
 AO21x1_ASAP7_75t_R _14854_ (.A1(_07657_),
    .A2(_07577_),
    .B(_07845_),
    .Y(_07846_));
 AO21x1_ASAP7_75t_R _14855_ (.A1(_07250_),
    .A2(_07253_),
    .B(_07078_),
    .Y(_07847_));
 OA211x2_ASAP7_75t_R _14856_ (.A1(_10092_),
    .A2(_07518_),
    .B(_07575_),
    .C(_07438_),
    .Y(_07848_));
 AOI211x1_ASAP7_75t_R _14857_ (.A1(_09949_),
    .A2(_07757_),
    .B(_07848_),
    .C(_07548_),
    .Y(_07849_));
 AOI21x1_ASAP7_75t_R _14858_ (.A1(_07671_),
    .A2(_07847_),
    .B(_07849_),
    .Y(_07850_));
 OR2x2_ASAP7_75t_R _14859_ (.A(_07276_),
    .B(_07850_),
    .Y(_07851_));
 OA211x2_ASAP7_75t_R _14860_ (.A1(_07647_),
    .A2(_07846_),
    .B(_07851_),
    .C(_07665_),
    .Y(_07852_));
 BUFx6f_ASAP7_75t_R _14861_ (.A(_07559_),
    .Y(_07853_));
 AND3x1_ASAP7_75t_R _14862_ (.A(_07080_),
    .B(_07560_),
    .C(_07563_),
    .Y(_07854_));
 AND3x1_ASAP7_75t_R _14863_ (.A(_07539_),
    .B(_07529_),
    .C(_07532_),
    .Y(_07855_));
 OR3x2_ASAP7_75t_R _14864_ (.A(_07647_),
    .B(_07854_),
    .C(_07855_),
    .Y(_07856_));
 NOR2x1_ASAP7_75t_R _14865_ (.A(_07853_),
    .B(_07856_),
    .Y(_07857_));
 OR3x1_ASAP7_75t_R _14866_ (.A(_07786_),
    .B(_07852_),
    .C(_07857_),
    .Y(_07858_));
 AND3x4_ASAP7_75t_R _14867_ (.A(_07835_),
    .B(_07844_),
    .C(_07858_),
    .Y(net58));
 INVx1_ASAP7_75t_R _14868_ (.A(_00931_),
    .Y(_07859_));
 INVx1_ASAP7_75t_R _14869_ (.A(_07353_),
    .Y(_07860_));
 NAND2x1_ASAP7_75t_R _14870_ (.A(_01209_),
    .B(_07346_),
    .Y(_07861_));
 AO21x1_ASAP7_75t_R _14871_ (.A1(_07860_),
    .A2(_07861_),
    .B(_07832_),
    .Y(_07862_));
 XNOR2x1_ASAP7_75t_R _14872_ (.B(_07862_),
    .Y(_07863_),
    .A(_00931_));
 INVx1_ASAP7_75t_R _14873_ (.A(_00930_),
    .Y(_07864_));
 AO22x1_ASAP7_75t_R _14874_ (.A1(_01206_),
    .A2(_07595_),
    .B1(_07635_),
    .B2(_07864_),
    .Y(_07865_));
 AO222x2_ASAP7_75t_R _14875_ (.A1(_07859_),
    .A2(_07639_),
    .B1(_07642_),
    .B2(_07863_),
    .C1(_07865_),
    .C2(_07634_),
    .Y(_07866_));
 OA211x2_ASAP7_75t_R _14876_ (.A1(_10087_),
    .A2(_07549_),
    .B(_07572_),
    .C(_03579_),
    .Y(_07867_));
 OA211x2_ASAP7_75t_R _14877_ (.A1(_07128_),
    .A2(_07549_),
    .B(_07575_),
    .C(_07235_),
    .Y(_07868_));
 OR2x2_ASAP7_75t_R _14878_ (.A(_07867_),
    .B(_07868_),
    .Y(_07869_));
 OA21x2_ASAP7_75t_R _14879_ (.A1(_07236_),
    .A2(_07650_),
    .B(_07757_),
    .Y(_07870_));
 AO21x2_ASAP7_75t_R _14880_ (.A1(_07702_),
    .A2(_07869_),
    .B(_07870_),
    .Y(_07871_));
 NAND2x1_ASAP7_75t_R _14881_ (.A(_07749_),
    .B(_07871_),
    .Y(_07872_));
 NAND2x1_ASAP7_75t_R _14882_ (.A(_07702_),
    .B(_07661_),
    .Y(_07873_));
 OA211x2_ASAP7_75t_R _14883_ (.A1(_07534_),
    .A2(_07670_),
    .B(_07873_),
    .C(_07489_),
    .Y(_07874_));
 AND3x1_ASAP7_75t_R _14884_ (.A(_07677_),
    .B(_07693_),
    .C(_07695_),
    .Y(_07875_));
 OA211x2_ASAP7_75t_R _14885_ (.A1(_07671_),
    .A2(_07672_),
    .B(_07676_),
    .C(_07533_),
    .Y(_07876_));
 OA21x2_ASAP7_75t_R _14886_ (.A1(_07875_),
    .A2(_07876_),
    .B(_06964_),
    .Y(_07877_));
 OR3x2_ASAP7_75t_R _14887_ (.A(_07647_),
    .B(_07874_),
    .C(_07877_),
    .Y(_07878_));
 NAND2x1_ASAP7_75t_R _14888_ (.A(_07872_),
    .B(_07878_),
    .Y(_07879_));
 OA211x2_ASAP7_75t_R _14889_ (.A1(_07548_),
    .A2(_07696_),
    .B(_07698_),
    .C(_07533_),
    .Y(_07880_));
 AO31x2_ASAP7_75t_R _14890_ (.A1(_07080_),
    .A2(_07703_),
    .A3(_07706_),
    .B(_07880_),
    .Y(_07881_));
 NOR2x1_ASAP7_75t_R _14891_ (.A(_06965_),
    .B(_07881_),
    .Y(_07882_));
 AND3x1_ASAP7_75t_R _14892_ (.A(_07718_),
    .B(_09953_),
    .C(_07186_),
    .Y(_07883_));
 OA21x2_ASAP7_75t_R _14893_ (.A1(_07719_),
    .A2(_07883_),
    .B(_07702_),
    .Y(_07884_));
 AOI22x1_ASAP7_75t_R _14894_ (.A1(_07076_),
    .A2(_07179_),
    .B1(_07255_),
    .B2(_07024_),
    .Y(_07885_));
 AOI22x1_ASAP7_75t_R _14895_ (.A1(_09953_),
    .A2(_07885_),
    .B1(_07719_),
    .B2(_07539_),
    .Y(_07886_));
 NAND2x1_ASAP7_75t_R _14896_ (.A(_04169_),
    .B(_07886_),
    .Y(_07887_));
 OA211x2_ASAP7_75t_R _14897_ (.A1(_04169_),
    .A2(_07884_),
    .B(_07887_),
    .C(_07727_),
    .Y(_07888_));
 NAND2x1_ASAP7_75t_R _14898_ (.A(_06866_),
    .B(_07516_),
    .Y(_07889_));
 INVx1_ASAP7_75t_R _14899_ (.A(_07889_),
    .Y(_07890_));
 OA21x2_ASAP7_75t_R _14900_ (.A1(_07882_),
    .A2(_07888_),
    .B(_07890_),
    .Y(_07891_));
 AO221x1_ASAP7_75t_R _14901_ (.A1(_07591_),
    .A2(_07866_),
    .B1(_07879_),
    .B2(_07682_),
    .C(_07891_),
    .Y(_07892_));
 BUFx4f_ASAP7_75t_R _14902_ (.A(_07892_),
    .Y(net59));
 BUFx4f_ASAP7_75t_R _14903_ (.A(_07506_),
    .Y(_07893_));
 NAND2x1_ASAP7_75t_R _14904_ (.A(_07578_),
    .B(_07752_),
    .Y(_07894_));
 AND2x2_ASAP7_75t_R _14905_ (.A(_03580_),
    .B(_07265_),
    .Y(_07895_));
 AOI211x1_ASAP7_75t_R _14906_ (.A1(_10077_),
    .A2(_07580_),
    .B(_07581_),
    .C(_07541_),
    .Y(_07896_));
 OR3x1_ASAP7_75t_R _14907_ (.A(_07080_),
    .B(_07895_),
    .C(_07896_),
    .Y(_07897_));
 AND3x1_ASAP7_75t_R _14908_ (.A(_07648_),
    .B(_07894_),
    .C(_07897_),
    .Y(_07898_));
 OR2x2_ASAP7_75t_R _14909_ (.A(_07657_),
    .B(_07733_),
    .Y(_07899_));
 OA211x2_ASAP7_75t_R _14910_ (.A1(_07081_),
    .A2(_07741_),
    .B(_07899_),
    .C(_07516_),
    .Y(_07900_));
 OR3x1_ASAP7_75t_R _14911_ (.A(_06966_),
    .B(_07898_),
    .C(_07900_),
    .Y(_07901_));
 AND2x2_ASAP7_75t_R _14912_ (.A(_07534_),
    .B(_07735_),
    .Y(_07902_));
 AO21x1_ASAP7_75t_R _14913_ (.A1(_07578_),
    .A2(_07769_),
    .B(_07902_),
    .Y(_07903_));
 OR3x1_ASAP7_75t_R _14914_ (.A(_07666_),
    .B(_07649_),
    .C(_07903_),
    .Y(_07904_));
 AOI21x1_ASAP7_75t_R _14915_ (.A1(_07579_),
    .A2(_07759_),
    .B(_07760_),
    .Y(_07905_));
 OR3x1_ASAP7_75t_R _14916_ (.A(_07677_),
    .B(_07770_),
    .C(_07771_),
    .Y(_07906_));
 OA211x2_ASAP7_75t_R _14917_ (.A1(_07540_),
    .A2(_07905_),
    .B(_07906_),
    .C(_07559_),
    .Y(_07907_));
 NOR2x2_ASAP7_75t_R _14918_ (.A(_07885_),
    .B(_07756_),
    .Y(_07908_));
 AND2x2_ASAP7_75t_R _14919_ (.A(_07538_),
    .B(_07908_),
    .Y(_07909_));
 OA21x2_ASAP7_75t_R _14920_ (.A1(_07907_),
    .A2(_07909_),
    .B(_07311_),
    .Y(_07910_));
 INVx1_ASAP7_75t_R _14921_ (.A(_07910_),
    .Y(_07911_));
 AO21x1_ASAP7_75t_R _14922_ (.A1(_09953_),
    .A2(_07885_),
    .B(_07908_),
    .Y(_07912_));
 AO21x1_ASAP7_75t_R _14923_ (.A1(_07538_),
    .A2(_07912_),
    .B(_07907_),
    .Y(_07913_));
 AOI21x1_ASAP7_75t_R _14924_ (.A1(_07277_),
    .A2(_07913_),
    .B(_07893_),
    .Y(_07914_));
 AO32x2_ASAP7_75t_R _14925_ (.A1(_07893_),
    .A2(_07901_),
    .A3(_07904_),
    .B1(_07911_),
    .B2(_07914_),
    .Y(_07915_));
 INVx1_ASAP7_75t_R _14926_ (.A(_01204_),
    .Y(_07916_));
 AO22x1_ASAP7_75t_R _14927_ (.A1(_01205_),
    .A2(_07596_),
    .B1(_07635_),
    .B2(_07916_),
    .Y(_07917_));
 AND2x2_ASAP7_75t_R _14928_ (.A(_07634_),
    .B(_07917_),
    .Y(_07918_));
 OA21x2_ASAP7_75t_R _14929_ (.A1(_07353_),
    .A2(_07599_),
    .B(_01207_),
    .Y(_07919_));
 OA21x2_ASAP7_75t_R _14930_ (.A1(_00931_),
    .A2(_07919_),
    .B(_00930_),
    .Y(_07920_));
 AO21x1_ASAP7_75t_R _14931_ (.A1(_07827_),
    .A2(_07920_),
    .B(_07828_),
    .Y(_07921_));
 OAI21x1_ASAP7_75t_R _14932_ (.A1(_07687_),
    .A2(_07920_),
    .B(_00897_),
    .Y(_07922_));
 OA21x2_ASAP7_75t_R _14933_ (.A1(_00897_),
    .A2(_07921_),
    .B(_07922_),
    .Y(_07923_));
 OAI21x1_ASAP7_75t_R _14934_ (.A1(_07918_),
    .A2(_07923_),
    .B(_07592_),
    .Y(_07924_));
 OAI21x1_ASAP7_75t_R _14935_ (.A1(_07592_),
    .A2(_07915_),
    .B(_07924_),
    .Y(net60));
 OA21x2_ASAP7_75t_R _14936_ (.A1(_04169_),
    .A2(_07305_),
    .B(_07324_),
    .Y(_07925_));
 AO21x1_ASAP7_75t_R _14937_ (.A1(_07666_),
    .A2(_07323_),
    .B(_07925_),
    .Y(_07926_));
 AO21x1_ASAP7_75t_R _14938_ (.A1(_07787_),
    .A2(_07788_),
    .B(_07540_),
    .Y(_07927_));
 OA211x2_ASAP7_75t_R _14939_ (.A1(_07081_),
    .A2(_07796_),
    .B(_07927_),
    .C(_07516_),
    .Y(_07928_));
 AO21x1_ASAP7_75t_R _14940_ (.A1(_07649_),
    .A2(_07273_),
    .B(_07928_),
    .Y(_07929_));
 NOR3x1_ASAP7_75t_R _14941_ (.A(_07447_),
    .B(_07450_),
    .C(_07461_),
    .Y(_07930_));
 OR3x1_ASAP7_75t_R _14942_ (.A(_07666_),
    .B(_07649_),
    .C(_07930_),
    .Y(_07931_));
 OAI21x1_ASAP7_75t_R _14943_ (.A1(_06966_),
    .A2(_07929_),
    .B(_07931_),
    .Y(_07932_));
 BUFx4f_ASAP7_75t_R _14944_ (.A(_07643_),
    .Y(_07933_));
 NOR2x1_ASAP7_75t_R _14945_ (.A(_07353_),
    .B(_07354_),
    .Y(_07934_));
 OAI21x1_ASAP7_75t_R _14946_ (.A1(_01207_),
    .A2(_07354_),
    .B(_07366_),
    .Y(_07935_));
 AO21x1_ASAP7_75t_R _14947_ (.A1(_07934_),
    .A2(_07861_),
    .B(_07935_),
    .Y(_07936_));
 XOR2x1_ASAP7_75t_R _14948_ (.A(_00864_),
    .Y(_07937_),
    .B(_07936_));
 NAND2x1_ASAP7_75t_R _14949_ (.A(_01203_),
    .B(_07777_),
    .Y(_07938_));
 OA21x2_ASAP7_75t_R _14950_ (.A1(_00863_),
    .A2(_07684_),
    .B(_07938_),
    .Y(_07939_));
 OA222x2_ASAP7_75t_R _14951_ (.A1(_00864_),
    .A2(_07688_),
    .B1(_07687_),
    .B2(_07937_),
    .C1(_07939_),
    .C2(_07594_),
    .Y(_07940_));
 NOR2x1_ASAP7_75t_R _14952_ (.A(_07933_),
    .B(_07940_),
    .Y(_07941_));
 AO221x2_ASAP7_75t_R _14953_ (.A1(_07890_),
    .A2(_07926_),
    .B1(_07932_),
    .B2(_07682_),
    .C(_07941_),
    .Y(net61));
 NAND2x1_ASAP7_75t_R _14954_ (.A(_07728_),
    .B(_07567_),
    .Y(_07942_));
 OAI21x1_ASAP7_75t_R _14955_ (.A1(_06966_),
    .A2(_07537_),
    .B(_07942_),
    .Y(_07943_));
 NAND2x1_ASAP7_75t_R _14956_ (.A(_10064_),
    .B(_07522_),
    .Y(_07944_));
 AOI211x1_ASAP7_75t_R _14957_ (.A1(_10079_),
    .A2(_07530_),
    .B(_07256_),
    .C(_07673_),
    .Y(_07945_));
 AO31x2_ASAP7_75t_R _14958_ (.A1(_03580_),
    .A2(_07574_),
    .A3(_07944_),
    .B(_07945_),
    .Y(_07946_));
 NOR2x2_ASAP7_75t_R _14959_ (.A(_07677_),
    .B(_07946_),
    .Y(_07947_));
 NAND2x1_ASAP7_75t_R _14960_ (.A(_07575_),
    .B(_07583_),
    .Y(_07948_));
 AO21x1_ASAP7_75t_R _14961_ (.A1(_07250_),
    .A2(_07253_),
    .B(_07718_),
    .Y(_07949_));
 OA211x2_ASAP7_75t_R _14962_ (.A1(_07671_),
    .A2(_07948_),
    .B(_07949_),
    .C(_07079_),
    .Y(_07950_));
 NAND2x1_ASAP7_75t_R _14963_ (.A(_07727_),
    .B(_07590_),
    .Y(_07951_));
 OA31x2_ASAP7_75t_R _14964_ (.A1(_07538_),
    .A2(_07947_),
    .A3(_07950_),
    .B1(_07951_),
    .Y(_07952_));
 AO21x1_ASAP7_75t_R _14965_ (.A1(_07648_),
    .A2(_07952_),
    .B(_06867_),
    .Y(_07953_));
 AO21x1_ASAP7_75t_R _14966_ (.A1(_07517_),
    .A2(_07943_),
    .B(_07953_),
    .Y(_07954_));
 AND2x2_ASAP7_75t_R _14967_ (.A(_09955_),
    .B(_06964_),
    .Y(_07955_));
 NOR2x2_ASAP7_75t_R _14968_ (.A(_07712_),
    .B(_07955_),
    .Y(_07956_));
 NOR2x2_ASAP7_75t_R _14969_ (.A(_07312_),
    .B(_07956_),
    .Y(_07957_));
 AO21x1_ASAP7_75t_R _14970_ (.A1(_07853_),
    .A2(_07558_),
    .B(_07957_),
    .Y(_07958_));
 OA21x2_ASAP7_75t_R _14971_ (.A1(_07893_),
    .A2(_07958_),
    .B(_07933_),
    .Y(_07959_));
 OA21x2_ASAP7_75t_R _14972_ (.A1(_07354_),
    .A2(_07919_),
    .B(_07366_),
    .Y(_07960_));
 OAI21x1_ASAP7_75t_R _14973_ (.A1(_00864_),
    .A2(_07960_),
    .B(_00863_),
    .Y(_07961_));
 OA21x2_ASAP7_75t_R _14974_ (.A1(_07830_),
    .A2(_07961_),
    .B(_07688_),
    .Y(_07962_));
 AND3x1_ASAP7_75t_R _14975_ (.A(_00830_),
    .B(_07642_),
    .C(_07961_),
    .Y(_07963_));
 INVx1_ASAP7_75t_R _14976_ (.A(_07963_),
    .Y(_07964_));
 NAND2x1_ASAP7_75t_R _14977_ (.A(_01202_),
    .B(_07777_),
    .Y(_07965_));
 OA21x2_ASAP7_75t_R _14978_ (.A1(_01201_),
    .A2(_07684_),
    .B(_07965_),
    .Y(_07966_));
 OA21x2_ASAP7_75t_R _14979_ (.A1(_07594_),
    .A2(_07966_),
    .B(_07591_),
    .Y(_07967_));
 OA211x2_ASAP7_75t_R _14980_ (.A1(_00830_),
    .A2(_07962_),
    .B(_07964_),
    .C(_07967_),
    .Y(_07968_));
 AOI21x1_ASAP7_75t_R _14981_ (.A1(_07954_),
    .A2(_07959_),
    .B(_07968_),
    .Y(net62));
 INVx1_ASAP7_75t_R _14982_ (.A(_00797_),
    .Y(_07969_));
 OA211x2_ASAP7_75t_R _14983_ (.A1(_07346_),
    .A2(_07355_),
    .B(_07358_),
    .C(_07368_),
    .Y(_07970_));
 XNOR2x1_ASAP7_75t_R _14984_ (.B(_07970_),
    .Y(_07971_),
    .A(_07969_));
 INVx1_ASAP7_75t_R _14985_ (.A(_00796_),
    .Y(_07972_));
 AO22x1_ASAP7_75t_R _14986_ (.A1(_01200_),
    .A2(_07595_),
    .B1(_07409_),
    .B2(_07972_),
    .Y(_07973_));
 AO222x2_ASAP7_75t_R _14987_ (.A1(_07969_),
    .A2(_07639_),
    .B1(_07386_),
    .B2(_07971_),
    .C1(_07973_),
    .C2(_07634_),
    .Y(_07974_));
 AOI211x1_ASAP7_75t_R _14988_ (.A1(_07657_),
    .A2(_07670_),
    .B(_07678_),
    .C(_07727_),
    .Y(_07975_));
 NOR2x1_ASAP7_75t_R _14989_ (.A(_07559_),
    .B(_07700_),
    .Y(_07976_));
 OA211x2_ASAP7_75t_R _14990_ (.A1(_10057_),
    .A2(_07530_),
    .B(_07571_),
    .C(_03579_),
    .Y(_07977_));
 AND3x1_ASAP7_75t_R _14991_ (.A(_07545_),
    .B(_07574_),
    .C(_07944_),
    .Y(_07978_));
 OR3x1_ASAP7_75t_R _14992_ (.A(_07438_),
    .B(_07867_),
    .C(_07868_),
    .Y(_07979_));
 OA31x2_ASAP7_75t_R _14993_ (.A1(_07079_),
    .A2(_07977_),
    .A3(_07978_),
    .B1(_07979_),
    .Y(_07980_));
 AND2x2_ASAP7_75t_R _14994_ (.A(_06964_),
    .B(_07652_),
    .Y(_07981_));
 AO211x2_ASAP7_75t_R _14995_ (.A1(_07489_),
    .A2(_07980_),
    .B(_07981_),
    .C(_07276_),
    .Y(_07982_));
 OA31x2_ASAP7_75t_R _14996_ (.A1(_07647_),
    .A2(_07975_),
    .A3(_07976_),
    .B1(_07982_),
    .Y(_07983_));
 AOI211x1_ASAP7_75t_R _14997_ (.A1(_07559_),
    .A2(_07710_),
    .B(_07955_),
    .C(_07310_),
    .Y(_07984_));
 AO31x2_ASAP7_75t_R _14998_ (.A1(_07310_),
    .A2(_07853_),
    .A3(_07721_),
    .B(_07984_),
    .Y(_07985_));
 AO222x2_ASAP7_75t_R _14999_ (.A1(_07591_),
    .A2(_07974_),
    .B1(_07983_),
    .B2(_07682_),
    .C1(_07985_),
    .C2(_07890_),
    .Y(net63));
 INVx1_ASAP7_75t_R _15000_ (.A(_01067_),
    .Y(_07986_));
 INVx1_ASAP7_75t_R _15001_ (.A(_07961_),
    .Y(_07987_));
 OA21x2_ASAP7_75t_R _15002_ (.A1(_00830_),
    .A2(_07987_),
    .B(_01201_),
    .Y(_07988_));
 OA21x2_ASAP7_75t_R _15003_ (.A1(_00797_),
    .A2(_07988_),
    .B(_00796_),
    .Y(_07989_));
 AO21x1_ASAP7_75t_R _15004_ (.A1(_07827_),
    .A2(_07989_),
    .B(_07828_),
    .Y(_07990_));
 INVx1_ASAP7_75t_R _15005_ (.A(_07989_),
    .Y(_07991_));
 INVx1_ASAP7_75t_R _15006_ (.A(_01215_),
    .Y(_07992_));
 AO22x1_ASAP7_75t_R _15007_ (.A1(_01216_),
    .A2(_07777_),
    .B1(_07635_),
    .B2(_07992_),
    .Y(_07993_));
 AO32x1_ASAP7_75t_R _15008_ (.A1(_01067_),
    .A2(_07827_),
    .A3(_07991_),
    .B1(_07993_),
    .B2(_07634_),
    .Y(_07994_));
 AO21x1_ASAP7_75t_R _15009_ (.A1(_07986_),
    .A2(_07990_),
    .B(_07994_),
    .Y(_07995_));
 OA211x2_ASAP7_75t_R _15010_ (.A1(_07578_),
    .A2(_07769_),
    .B(_07772_),
    .C(_07727_),
    .Y(_07996_));
 AOI21x1_ASAP7_75t_R _15011_ (.A1(_07853_),
    .A2(_07737_),
    .B(_07996_),
    .Y(_07997_));
 OA21x2_ASAP7_75t_R _15012_ (.A1(_07895_),
    .A2(_07896_),
    .B(_07080_),
    .Y(_07998_));
 AO21x1_ASAP7_75t_R _15013_ (.A1(_10102_),
    .A2(_07550_),
    .B(_07739_),
    .Y(_07999_));
 AND2x2_ASAP7_75t_R _15014_ (.A(_10069_),
    .B(_07530_),
    .Y(_08000_));
 AO221x1_ASAP7_75t_R _15015_ (.A1(_03576_),
    .A2(_03577_),
    .B1(_10059_),
    .B2(_07580_),
    .C(_08000_),
    .Y(_08001_));
 OA211x2_ASAP7_75t_R _15016_ (.A1(_07579_),
    .A2(_07999_),
    .B(_08001_),
    .C(_07539_),
    .Y(_08002_));
 NAND3x1_ASAP7_75t_R _15017_ (.A(_06964_),
    .B(_07534_),
    .C(_07752_),
    .Y(_08003_));
 OA31x2_ASAP7_75t_R _15018_ (.A1(_06965_),
    .A2(_07998_),
    .A3(_08002_),
    .B1(_08003_),
    .Y(_08004_));
 NAND2x1_ASAP7_75t_R _15019_ (.A(_07648_),
    .B(_08004_),
    .Y(_08005_));
 OA211x2_ASAP7_75t_R _15020_ (.A1(_07649_),
    .A2(_07997_),
    .B(_08005_),
    .C(_07893_),
    .Y(_08006_));
 AOI21x1_ASAP7_75t_R _15021_ (.A1(_07186_),
    .A2(_07712_),
    .B(_07290_),
    .Y(_08007_));
 AO32x1_ASAP7_75t_R _15022_ (.A1(_07541_),
    .A2(_09959_),
    .A3(_07580_),
    .B1(_08007_),
    .B2(_09953_),
    .Y(_08008_));
 INVx1_ASAP7_75t_R _15023_ (.A(_08008_),
    .Y(_08009_));
 OA211x2_ASAP7_75t_R _15024_ (.A1(_07657_),
    .A2(_08009_),
    .B(_07761_),
    .C(_07559_),
    .Y(_08010_));
 NOR2x1_ASAP7_75t_R _15025_ (.A(_07957_),
    .B(_08010_),
    .Y(_08011_));
 AO21x1_ASAP7_75t_R _15026_ (.A1(_06867_),
    .A2(_08011_),
    .B(_07591_),
    .Y(_08012_));
 OA22x2_ASAP7_75t_R _15027_ (.A1(_07933_),
    .A2(_07995_),
    .B1(_08006_),
    .B2(_08012_),
    .Y(net33));
 OR2x2_ASAP7_75t_R _15028_ (.A(_00796_),
    .B(_01067_),
    .Y(_08013_));
 OA211x2_ASAP7_75t_R _15029_ (.A1(_07351_),
    .A2(_07970_),
    .B(_08013_),
    .C(_01215_),
    .Y(_08014_));
 XNOR2x1_ASAP7_75t_R _15030_ (.B(_08014_),
    .Y(_08015_),
    .A(_00731_));
 NAND2x1_ASAP7_75t_R _15031_ (.A(_01199_),
    .B(_07596_),
    .Y(_08016_));
 OA21x2_ASAP7_75t_R _15032_ (.A1(_01198_),
    .A2(_07684_),
    .B(_08016_),
    .Y(_08017_));
 OA222x2_ASAP7_75t_R _15033_ (.A1(_00731_),
    .A2(_07688_),
    .B1(_07687_),
    .B2(_08015_),
    .C1(_08017_),
    .C2(_07594_),
    .Y(_08018_));
 AO221x1_ASAP7_75t_R _15034_ (.A1(_07521_),
    .A2(_07802_),
    .B1(_07803_),
    .B2(_07250_),
    .C(_07079_),
    .Y(_08019_));
 NAND2x1_ASAP7_75t_R _15035_ (.A(_06964_),
    .B(_07243_),
    .Y(_08020_));
 OR2x2_ASAP7_75t_R _15036_ (.A(_06431_),
    .B(_07549_),
    .Y(_08021_));
 AO21x1_ASAP7_75t_R _15037_ (.A1(_07730_),
    .A2(_08021_),
    .B(_07078_),
    .Y(_08022_));
 OA211x2_ASAP7_75t_R _15038_ (.A1(_07533_),
    .A2(_07257_),
    .B(_08022_),
    .C(_03580_),
    .Y(_08023_));
 OR2x2_ASAP7_75t_R _15039_ (.A(_07438_),
    .B(_07265_),
    .Y(_08024_));
 OA211x2_ASAP7_75t_R _15040_ (.A1(_07079_),
    .A2(_07999_),
    .B(_08024_),
    .C(_07521_),
    .Y(_08025_));
 OR3x1_ASAP7_75t_R _15041_ (.A(_07244_),
    .B(_08023_),
    .C(_08025_),
    .Y(_08026_));
 OAI21x1_ASAP7_75t_R _15042_ (.A1(_08019_),
    .A2(_08020_),
    .B(_08026_),
    .Y(_08027_));
 OA21x2_ASAP7_75t_R _15043_ (.A1(_07853_),
    .A2(_07811_),
    .B(_07517_),
    .Y(_08028_));
 OA21x2_ASAP7_75t_R _15044_ (.A1(_06966_),
    .A2(_07794_),
    .B(_08028_),
    .Y(_08029_));
 OAI21x1_ASAP7_75t_R _15045_ (.A1(_08027_),
    .A2(_08029_),
    .B(_07682_),
    .Y(_08030_));
 AND3x1_ASAP7_75t_R _15046_ (.A(_09953_),
    .B(_07080_),
    .C(_07290_),
    .Y(_08031_));
 OAI21x1_ASAP7_75t_R _15047_ (.A1(_07814_),
    .A2(_08031_),
    .B(_07312_),
    .Y(_08032_));
 OA21x2_ASAP7_75t_R _15048_ (.A1(_06965_),
    .A2(_07081_),
    .B(_09953_),
    .Y(_08033_));
 AO21x1_ASAP7_75t_R _15049_ (.A1(_07666_),
    .A2(_07814_),
    .B(_08033_),
    .Y(_08034_));
 NAND2x1_ASAP7_75t_R _15050_ (.A(_07277_),
    .B(_08034_),
    .Y(_08035_));
 AO21x1_ASAP7_75t_R _15051_ (.A1(_08032_),
    .A2(_08035_),
    .B(_07775_),
    .Y(_08036_));
 OA211x2_ASAP7_75t_R _15052_ (.A1(_07933_),
    .A2(_08018_),
    .B(_08030_),
    .C(_08036_),
    .Y(_08037_));
 INVx1_ASAP7_75t_R _15053_ (.A(_08037_),
    .Y(net34));
 AND3x1_ASAP7_75t_R _15054_ (.A(_07666_),
    .B(_07535_),
    .C(_07556_),
    .Y(_08038_));
 OA211x2_ASAP7_75t_R _15055_ (.A1(_06966_),
    .A2(_07081_),
    .B(_09953_),
    .C(_04169_),
    .Y(_08039_));
 OAI21x1_ASAP7_75t_R _15056_ (.A1(_08038_),
    .A2(_08039_),
    .B(_07517_),
    .Y(_08040_));
 NAND2x1_ASAP7_75t_R _15057_ (.A(_01197_),
    .B(_07596_),
    .Y(_08041_));
 OA21x2_ASAP7_75t_R _15058_ (.A1(_01196_),
    .A2(_07684_),
    .B(_08041_),
    .Y(_08042_));
 NAND2x2_ASAP7_75t_R _15059_ (.A(_07361_),
    .B(_07603_),
    .Y(_08043_));
 NAND2x1_ASAP7_75t_R _15060_ (.A(_00698_),
    .B(_08043_),
    .Y(_08044_));
 OA21x2_ASAP7_75t_R _15061_ (.A1(_07687_),
    .A2(_08043_),
    .B(_07688_),
    .Y(_08045_));
 OA222x2_ASAP7_75t_R _15062_ (.A1(_07594_),
    .A2(_08042_),
    .B1(_08044_),
    .B2(_07687_),
    .C1(_08045_),
    .C2(_00698_),
    .Y(_08046_));
 AO21x1_ASAP7_75t_R _15063_ (.A1(_10102_),
    .A2(_07552_),
    .B(_07528_),
    .Y(_08047_));
 AND3x1_ASAP7_75t_R _15064_ (.A(_07548_),
    .B(_07730_),
    .C(_08021_),
    .Y(_08048_));
 AO21x2_ASAP7_75t_R _15065_ (.A1(_07541_),
    .A2(_08047_),
    .B(_08048_),
    .Y(_08049_));
 NOR2x1_ASAP7_75t_R _15066_ (.A(_07534_),
    .B(_07946_),
    .Y(_08050_));
 AO21x1_ASAP7_75t_R _15067_ (.A1(_07540_),
    .A2(_08049_),
    .B(_08050_),
    .Y(_08051_));
 OA21x2_ASAP7_75t_R _15068_ (.A1(_07517_),
    .A2(_08051_),
    .B(_07856_),
    .Y(_08052_));
 OA21x2_ASAP7_75t_R _15069_ (.A1(_07535_),
    .A2(_07547_),
    .B(_07837_),
    .Y(_08053_));
 OA21x2_ASAP7_75t_R _15070_ (.A1(_07516_),
    .A2(_07850_),
    .B(_07728_),
    .Y(_08054_));
 OAI21x1_ASAP7_75t_R _15071_ (.A1(_07649_),
    .A2(_08053_),
    .B(_08054_),
    .Y(_08055_));
 OA211x2_ASAP7_75t_R _15072_ (.A1(_06966_),
    .A2(_08052_),
    .B(_08055_),
    .C(_07682_),
    .Y(_08056_));
 AO221x2_ASAP7_75t_R _15073_ (.A1(_07692_),
    .A2(_08040_),
    .B1(_08046_),
    .B2(_07592_),
    .C(_08056_),
    .Y(_08057_));
 INVx1_ASAP7_75t_R _15074_ (.A(_08057_),
    .Y(net35));
 AO21x1_ASAP7_75t_R _15075_ (.A1(_09953_),
    .A2(_07885_),
    .B(_06963_),
    .Y(_08058_));
 AO21x1_ASAP7_75t_R _15076_ (.A1(_07702_),
    .A2(_07719_),
    .B(_08058_),
    .Y(_08059_));
 AOI22x1_ASAP7_75t_R _15077_ (.A1(_07312_),
    .A2(_07884_),
    .B1(_07956_),
    .B2(_08059_),
    .Y(_08060_));
 OR3x1_ASAP7_75t_R _15078_ (.A(_07538_),
    .B(_07875_),
    .C(_07876_),
    .Y(_08061_));
 OA21x2_ASAP7_75t_R _15079_ (.A1(_07666_),
    .A2(_07881_),
    .B(_08061_),
    .Y(_08062_));
 OA21x2_ASAP7_75t_R _15080_ (.A1(_07977_),
    .A2(_07978_),
    .B(_07677_),
    .Y(_08063_));
 NAND2x1_ASAP7_75t_R _15081_ (.A(_10042_),
    .B(_07550_),
    .Y(_08064_));
 AND3x1_ASAP7_75t_R _15082_ (.A(_03580_),
    .B(_07523_),
    .C(_08064_),
    .Y(_08065_));
 AOI211x1_ASAP7_75t_R _15083_ (.A1(_07570_),
    .A2(_08047_),
    .B(_08065_),
    .C(_07677_),
    .Y(_08066_));
 OR2x2_ASAP7_75t_R _15084_ (.A(_07559_),
    .B(_07871_),
    .Y(_08067_));
 OA31x2_ASAP7_75t_R _15085_ (.A1(_07538_),
    .A2(_08063_),
    .A3(_08066_),
    .B1(_08067_),
    .Y(_08068_));
 NAND2x1_ASAP7_75t_R _15086_ (.A(_07649_),
    .B(_08068_),
    .Y(_08069_));
 OA211x2_ASAP7_75t_R _15087_ (.A1(_07649_),
    .A2(_08062_),
    .B(_08069_),
    .C(_07893_),
    .Y(_08070_));
 AO21x2_ASAP7_75t_R _15088_ (.A1(_06867_),
    .A2(_08060_),
    .B(_08070_),
    .Y(_08071_));
 OR2x2_ASAP7_75t_R _15089_ (.A(_00698_),
    .B(_00731_),
    .Y(_08072_));
 OA21x2_ASAP7_75t_R _15090_ (.A1(_00698_),
    .A2(_01198_),
    .B(_01196_),
    .Y(_08073_));
 OA21x2_ASAP7_75t_R _15091_ (.A1(_08014_),
    .A2(_08072_),
    .B(_08073_),
    .Y(_08074_));
 XNOR2x1_ASAP7_75t_R _15092_ (.B(_08074_),
    .Y(_08075_),
    .A(_00665_));
 OR2x2_ASAP7_75t_R _15093_ (.A(_07687_),
    .B(_08075_),
    .Y(_08076_));
 NAND2x1_ASAP7_75t_R _15094_ (.A(_01195_),
    .B(_07777_),
    .Y(_08077_));
 OA21x2_ASAP7_75t_R _15095_ (.A1(_01194_),
    .A2(_07684_),
    .B(_08077_),
    .Y(_08078_));
 OA22x2_ASAP7_75t_R _15096_ (.A1(_00665_),
    .A2(_07688_),
    .B1(_08078_),
    .B2(_07594_),
    .Y(_08079_));
 AO21x1_ASAP7_75t_R _15097_ (.A1(_08076_),
    .A2(_08079_),
    .B(_07933_),
    .Y(_08080_));
 OAI21x1_ASAP7_75t_R _15098_ (.A1(_07592_),
    .A2(_08071_),
    .B(_08080_),
    .Y(net36));
 OA211x2_ASAP7_75t_R _15099_ (.A1(_07570_),
    .A2(_07999_),
    .B(_08001_),
    .C(_07677_),
    .Y(_08081_));
 AND2x2_ASAP7_75t_R _15100_ (.A(_07523_),
    .B(_08064_),
    .Y(_08082_));
 OR3x1_ASAP7_75t_R _15101_ (.A(_07548_),
    .B(_07675_),
    .C(_07667_),
    .Y(_08083_));
 OA211x2_ASAP7_75t_R _15102_ (.A1(_07729_),
    .A2(_08082_),
    .B(_08083_),
    .C(_07702_),
    .Y(_08084_));
 OR3x1_ASAP7_75t_R _15103_ (.A(_07727_),
    .B(_08081_),
    .C(_08084_),
    .Y(_08085_));
 AO21x1_ASAP7_75t_R _15104_ (.A1(_07894_),
    .A2(_07897_),
    .B(_07665_),
    .Y(_08086_));
 AND3x1_ASAP7_75t_R _15105_ (.A(_07648_),
    .B(_08085_),
    .C(_08086_),
    .Y(_08087_));
 OAI21x1_ASAP7_75t_R _15106_ (.A1(_07535_),
    .A2(_07905_),
    .B(_07906_),
    .Y(_08088_));
 AND3x1_ASAP7_75t_R _15107_ (.A(_07728_),
    .B(_07516_),
    .C(_08088_),
    .Y(_08089_));
 AND3x1_ASAP7_75t_R _15108_ (.A(_07853_),
    .B(_07516_),
    .C(_07903_),
    .Y(_08090_));
 OR4x2_ASAP7_75t_R _15109_ (.A(_07786_),
    .B(_08087_),
    .C(_08089_),
    .D(_08090_),
    .Y(_08091_));
 AOI21x1_ASAP7_75t_R _15110_ (.A1(_07956_),
    .A2(_08058_),
    .B(_07908_),
    .Y(_08092_));
 OR3x4_ASAP7_75t_R _15111_ (.A(_07775_),
    .B(_07957_),
    .C(_08092_),
    .Y(_08093_));
 INVx1_ASAP7_75t_R _15112_ (.A(_08043_),
    .Y(_08094_));
 OA21x2_ASAP7_75t_R _15113_ (.A1(_00698_),
    .A2(_08094_),
    .B(_01196_),
    .Y(_08095_));
 OA21x2_ASAP7_75t_R _15114_ (.A1(_00665_),
    .A2(_08095_),
    .B(_01194_),
    .Y(_08096_));
 NAND2x1_ASAP7_75t_R _15115_ (.A(_07827_),
    .B(_08096_),
    .Y(_08097_));
 AO21x1_ASAP7_75t_R _15116_ (.A1(_07688_),
    .A2(_08097_),
    .B(_00632_),
    .Y(_08098_));
 INVx1_ASAP7_75t_R _15117_ (.A(_01192_),
    .Y(_08099_));
 AO22x1_ASAP7_75t_R _15118_ (.A1(_01193_),
    .A2(_07777_),
    .B1(_07635_),
    .B2(_08099_),
    .Y(_08100_));
 NOR2x1_ASAP7_75t_R _15119_ (.A(_07830_),
    .B(_08096_),
    .Y(_08101_));
 AOI22x1_ASAP7_75t_R _15120_ (.A1(_07634_),
    .A2(_08100_),
    .B1(_08101_),
    .B2(_00632_),
    .Y(_08102_));
 AO21x1_ASAP7_75t_R _15121_ (.A1(_08098_),
    .A2(_08102_),
    .B(_07933_),
    .Y(_08103_));
 NAND3x2_ASAP7_75t_R _15122_ (.B(_08093_),
    .C(_08103_),
    .Y(net37),
    .A(_08091_));
 OA21x2_ASAP7_75t_R _15123_ (.A1(_09953_),
    .A2(_07506_),
    .B(_07277_),
    .Y(_08104_));
 AO21x1_ASAP7_75t_R _15124_ (.A1(_07506_),
    .A2(_07311_),
    .B(_08104_),
    .Y(_08105_));
 OA21x2_ASAP7_75t_R _15125_ (.A1(_06867_),
    .A2(_07569_),
    .B(_08105_),
    .Y(_08106_));
 OR3x1_ASAP7_75t_R _15126_ (.A(_07545_),
    .B(_07449_),
    .C(_07527_),
    .Y(_08107_));
 NOR2x1_ASAP7_75t_R _15127_ (.A(_10042_),
    .B(_07518_),
    .Y(_08108_));
 AO221x1_ASAP7_75t_R _15128_ (.A1(_03576_),
    .A2(_03577_),
    .B1(_10034_),
    .B2(_07550_),
    .C(_08108_),
    .Y(_08109_));
 AND3x1_ASAP7_75t_R _15129_ (.A(_07702_),
    .B(_08107_),
    .C(_08109_),
    .Y(_08110_));
 AOI211x1_ASAP7_75t_R _15130_ (.A1(_07578_),
    .A2(_08049_),
    .B(_08110_),
    .C(_07727_),
    .Y(_08111_));
 NOR3x1_ASAP7_75t_R _15131_ (.A(_07559_),
    .B(_07947_),
    .C(_07950_),
    .Y(_08112_));
 OA21x2_ASAP7_75t_R _15132_ (.A1(_08111_),
    .A2(_08112_),
    .B(_07506_),
    .Y(_08113_));
 AND3x1_ASAP7_75t_R _15133_ (.A(_06866_),
    .B(_07665_),
    .C(_07590_),
    .Y(_08114_));
 OA211x2_ASAP7_75t_R _15134_ (.A1(_08113_),
    .A2(_08114_),
    .B(_07643_),
    .C(_07648_),
    .Y(_08115_));
 AO21x1_ASAP7_75t_R _15135_ (.A1(_07363_),
    .A2(_07605_),
    .B(_00599_),
    .Y(_08116_));
 AND2x2_ASAP7_75t_R _15136_ (.A(_00598_),
    .B(_08116_),
    .Y(_08117_));
 XNOR2x1_ASAP7_75t_R _15137_ (.B(_08117_),
    .Y(_08118_),
    .A(_00565_));
 NAND2x1_ASAP7_75t_R _15138_ (.A(_01190_),
    .B(_07595_),
    .Y(_08119_));
 OA21x2_ASAP7_75t_R _15139_ (.A1(_01189_),
    .A2(_07424_),
    .B(_08119_),
    .Y(_08120_));
 OA222x2_ASAP7_75t_R _15140_ (.A1(_00565_),
    .A2(_07688_),
    .B1(_07430_),
    .B2(_08118_),
    .C1(_08120_),
    .C2(_07423_),
    .Y(_08121_));
 NOR2x1_ASAP7_75t_R _15141_ (.A(_07643_),
    .B(_08121_),
    .Y(_08122_));
 OR3x4_ASAP7_75t_R _15142_ (.A(_08106_),
    .B(_08115_),
    .C(_08122_),
    .Y(net39));
 OR2x2_ASAP7_75t_R _15143_ (.A(_00565_),
    .B(_00599_),
    .Y(_08123_));
 OA21x2_ASAP7_75t_R _15144_ (.A1(_08123_),
    .A2(_07419_),
    .B(_07394_),
    .Y(_08124_));
 XNOR2x1_ASAP7_75t_R _15145_ (.B(_08124_),
    .Y(_08125_),
    .A(_00532_));
 NAND2x1_ASAP7_75t_R _15146_ (.A(_01188_),
    .B(_07777_),
    .Y(_08126_));
 OA21x2_ASAP7_75t_R _15147_ (.A1(_01187_),
    .A2(_07684_),
    .B(_08126_),
    .Y(_08127_));
 OA222x2_ASAP7_75t_R _15148_ (.A1(_00532_),
    .A2(_07688_),
    .B1(_07687_),
    .B2(_08125_),
    .C1(_08127_),
    .C2(_07594_),
    .Y(_08128_));
 AND2x2_ASAP7_75t_R _15149_ (.A(_06965_),
    .B(_07647_),
    .Y(_08129_));
 AO21x2_ASAP7_75t_R _15150_ (.A1(_10034_),
    .A2(_07186_),
    .B(_07562_),
    .Y(_08130_));
 OA21x2_ASAP7_75t_R _15151_ (.A1(_07449_),
    .A2(_07527_),
    .B(_07521_),
    .Y(_08131_));
 AOI21x1_ASAP7_75t_R _15152_ (.A1(_07729_),
    .A2(_08130_),
    .B(_08131_),
    .Y(_08132_));
 AOI211x1_ASAP7_75t_R _15153_ (.A1(_07570_),
    .A2(_08047_),
    .B(_08065_),
    .C(_07539_),
    .Y(_08133_));
 AO21x1_ASAP7_75t_R _15154_ (.A1(_07534_),
    .A2(_08132_),
    .B(_08133_),
    .Y(_08134_));
 AOI22x1_ASAP7_75t_R _15155_ (.A1(_07980_),
    .A2(_08129_),
    .B1(_08134_),
    .B2(_07749_),
    .Y(_08135_));
 AO21x1_ASAP7_75t_R _15156_ (.A1(_07724_),
    .A2(_08135_),
    .B(_06867_),
    .Y(_08136_));
 AOI21x1_ASAP7_75t_R _15157_ (.A1(_07749_),
    .A2(_07652_),
    .B(_08104_),
    .Y(_08137_));
 AO21x1_ASAP7_75t_R _15158_ (.A1(_07893_),
    .A2(_07713_),
    .B(_08137_),
    .Y(_08138_));
 AO21x1_ASAP7_75t_R _15159_ (.A1(_08136_),
    .A2(_08138_),
    .B(_07592_),
    .Y(_08139_));
 OAI21x1_ASAP7_75t_R _15160_ (.A1(_07933_),
    .A2(_08128_),
    .B(_08139_),
    .Y(net40));
 OR4x1_ASAP7_75t_R _15161_ (.A(_04169_),
    .B(_06866_),
    .C(_07648_),
    .D(_07762_),
    .Y(_08140_));
 AO21x1_ASAP7_75t_R _15162_ (.A1(_09955_),
    .A2(_06866_),
    .B(_07712_),
    .Y(_08141_));
 AO21x1_ASAP7_75t_R _15163_ (.A1(_07715_),
    .A2(_07762_),
    .B(_08141_),
    .Y(_08142_));
 AO21x1_ASAP7_75t_R _15164_ (.A1(_08140_),
    .A2(_08142_),
    .B(_07773_),
    .Y(_08143_));
 AND2x4_ASAP7_75t_R _15165_ (.A(_07692_),
    .B(_08141_),
    .Y(_08144_));
 NAND2x1_ASAP7_75t_R _15166_ (.A(_07753_),
    .B(_08144_),
    .Y(_08145_));
 OA21x2_ASAP7_75t_R _15167_ (.A1(_07674_),
    .A2(_07694_),
    .B(_07729_),
    .Y(_08146_));
 AO21x1_ASAP7_75t_R _15168_ (.A1(_07579_),
    .A2(_08130_),
    .B(_08146_),
    .Y(_08147_));
 OA211x2_ASAP7_75t_R _15169_ (.A1(_03581_),
    .A2(_08082_),
    .B(_08083_),
    .C(_07080_),
    .Y(_08148_));
 AO21x2_ASAP7_75t_R _15170_ (.A1(_07540_),
    .A2(_08147_),
    .B(_08148_),
    .Y(_08149_));
 OR3x1_ASAP7_75t_R _15171_ (.A(_07665_),
    .B(_07998_),
    .C(_08002_),
    .Y(_08150_));
 OAI21x1_ASAP7_75t_R _15172_ (.A1(_07728_),
    .A2(_08149_),
    .B(_08150_),
    .Y(_08151_));
 AO21x1_ASAP7_75t_R _15173_ (.A1(_07649_),
    .A2(_08151_),
    .B(_07786_),
    .Y(_08152_));
 NAND2x1_ASAP7_75t_R _15174_ (.A(_08145_),
    .B(_08152_),
    .Y(_08153_));
 OA21x2_ASAP7_75t_R _15175_ (.A1(_00565_),
    .A2(_07608_),
    .B(_01189_),
    .Y(_08154_));
 OA21x2_ASAP7_75t_R _15176_ (.A1(_00532_),
    .A2(_08154_),
    .B(_01187_),
    .Y(_08155_));
 OA21x2_ASAP7_75t_R _15177_ (.A1(_07347_),
    .A2(_07605_),
    .B(_08155_),
    .Y(_08156_));
 AOI21x1_ASAP7_75t_R _15178_ (.A1(_07642_),
    .A2(_08156_),
    .B(_07828_),
    .Y(_08157_));
 INVx1_ASAP7_75t_R _15179_ (.A(_00499_),
    .Y(_08158_));
 OR3x1_ASAP7_75t_R _15180_ (.A(_08158_),
    .B(_07430_),
    .C(_08156_),
    .Y(_08159_));
 NAND2x1_ASAP7_75t_R _15181_ (.A(_01186_),
    .B(_07595_),
    .Y(_08160_));
 OA21x2_ASAP7_75t_R _15182_ (.A1(_01185_),
    .A2(_07424_),
    .B(_08160_),
    .Y(_08161_));
 OA21x2_ASAP7_75t_R _15183_ (.A1(_07423_),
    .A2(_08161_),
    .B(_07336_),
    .Y(_08162_));
 OA211x2_ASAP7_75t_R _15184_ (.A1(_00499_),
    .A2(_08157_),
    .B(_08159_),
    .C(_08162_),
    .Y(_08163_));
 AO21x2_ASAP7_75t_R _15185_ (.A1(_08143_),
    .A2(_08153_),
    .B(_08163_),
    .Y(_08164_));
 INVx1_ASAP7_75t_R _15186_ (.A(_08164_),
    .Y(net41));
 OA21x2_ASAP7_75t_R _15187_ (.A1(_07348_),
    .A2(_07419_),
    .B(_07396_),
    .Y(_08165_));
 AND2x2_ASAP7_75t_R _15188_ (.A(_07827_),
    .B(_08165_),
    .Y(_08166_));
 OR3x1_ASAP7_75t_R _15189_ (.A(_00466_),
    .B(_07828_),
    .C(_08166_),
    .Y(_08167_));
 OAI21x1_ASAP7_75t_R _15190_ (.A1(_07687_),
    .A2(_08165_),
    .B(_00466_),
    .Y(_08168_));
 INVx1_ASAP7_75t_R _15191_ (.A(_01183_),
    .Y(_08169_));
 AO22x1_ASAP7_75t_R _15192_ (.A1(_01184_),
    .A2(_07596_),
    .B1(_07635_),
    .B2(_08169_),
    .Y(_08170_));
 AO21x1_ASAP7_75t_R _15193_ (.A1(_07634_),
    .A2(_08170_),
    .B(_07643_),
    .Y(_08171_));
 AO21x1_ASAP7_75t_R _15194_ (.A1(_08167_),
    .A2(_08168_),
    .B(_08171_),
    .Y(_08172_));
 OR3x1_ASAP7_75t_R _15195_ (.A(_07438_),
    .B(_07675_),
    .C(_07667_),
    .Y(_08173_));
 OR3x1_ASAP7_75t_R _15196_ (.A(_07078_),
    .B(_07674_),
    .C(_07694_),
    .Y(_08174_));
 AND3x1_ASAP7_75t_R _15197_ (.A(_07671_),
    .B(_08173_),
    .C(_08174_),
    .Y(_08175_));
 AO21x1_ASAP7_75t_R _15198_ (.A1(_10034_),
    .A2(_07550_),
    .B(_08108_),
    .Y(_08176_));
 OR3x1_ASAP7_75t_R _15199_ (.A(_07078_),
    .B(_07765_),
    .C(_07790_),
    .Y(_08177_));
 OA211x2_ASAP7_75t_R _15200_ (.A1(_07533_),
    .A2(_08176_),
    .B(_08177_),
    .C(_07541_),
    .Y(_08178_));
 OR3x1_ASAP7_75t_R _15201_ (.A(_07538_),
    .B(_08175_),
    .C(_08178_),
    .Y(_08179_));
 OR3x1_ASAP7_75t_R _15202_ (.A(_07853_),
    .B(_08023_),
    .C(_08025_),
    .Y(_08180_));
 NAND2x1_ASAP7_75t_R _15203_ (.A(_08179_),
    .B(_08180_),
    .Y(_08181_));
 AO21x1_ASAP7_75t_R _15204_ (.A1(_07649_),
    .A2(_08181_),
    .B(_07818_),
    .Y(_08182_));
 OR3x1_ASAP7_75t_R _15205_ (.A(_07775_),
    .B(_07805_),
    .C(_08104_),
    .Y(_08183_));
 OA21x2_ASAP7_75t_R _15206_ (.A1(_07786_),
    .A2(_08182_),
    .B(_08183_),
    .Y(_08184_));
 AND2x4_ASAP7_75t_R _15207_ (.A(_08172_),
    .B(_08184_),
    .Y(net42));
 AO21x1_ASAP7_75t_R _15208_ (.A1(_10009_),
    .A2(_07580_),
    .B(_07448_),
    .Y(_08185_));
 OR3x1_ASAP7_75t_R _15209_ (.A(_07729_),
    .B(_07765_),
    .C(_07790_),
    .Y(_08186_));
 OA21x2_ASAP7_75t_R _15210_ (.A1(_07579_),
    .A2(_08185_),
    .B(_08186_),
    .Y(_08187_));
 AO21x1_ASAP7_75t_R _15211_ (.A1(_08107_),
    .A2(_08109_),
    .B(_07657_),
    .Y(_08188_));
 OAI21x1_ASAP7_75t_R _15212_ (.A1(_07081_),
    .A2(_08187_),
    .B(_08188_),
    .Y(_08189_));
 NAND2x1_ASAP7_75t_R _15213_ (.A(_07728_),
    .B(_08051_),
    .Y(_08190_));
 OA21x2_ASAP7_75t_R _15214_ (.A1(_06966_),
    .A2(_08189_),
    .B(_08190_),
    .Y(_08191_));
 AND2x2_ASAP7_75t_R _15215_ (.A(_07893_),
    .B(_07648_),
    .Y(_08192_));
 AO21x1_ASAP7_75t_R _15216_ (.A1(_07749_),
    .A2(_07850_),
    .B(_08104_),
    .Y(_08193_));
 OA21x2_ASAP7_75t_R _15217_ (.A1(_06867_),
    .A2(_07843_),
    .B(_08193_),
    .Y(_08194_));
 AO221x2_ASAP7_75t_R _15218_ (.A1(_07893_),
    .A2(_07840_),
    .B1(_08191_),
    .B2(_08192_),
    .C(_08194_),
    .Y(_08195_));
 INVx1_ASAP7_75t_R _15219_ (.A(_00433_),
    .Y(_08196_));
 OA21x2_ASAP7_75t_R _15220_ (.A1(_00499_),
    .A2(_08156_),
    .B(_01185_),
    .Y(_08197_));
 OA21x2_ASAP7_75t_R _15221_ (.A1(_00466_),
    .A2(_08197_),
    .B(_01183_),
    .Y(_08198_));
 AO21x1_ASAP7_75t_R _15222_ (.A1(_07827_),
    .A2(_08198_),
    .B(_07828_),
    .Y(_08199_));
 INVx1_ASAP7_75t_R _15223_ (.A(_08198_),
    .Y(_08200_));
 INVx1_ASAP7_75t_R _15224_ (.A(_01181_),
    .Y(_08201_));
 AO22x1_ASAP7_75t_R _15225_ (.A1(_01182_),
    .A2(_07777_),
    .B1(_07635_),
    .B2(_08201_),
    .Y(_08202_));
 AO32x1_ASAP7_75t_R _15226_ (.A1(_00433_),
    .A2(_07642_),
    .A3(_08200_),
    .B1(_08202_),
    .B2(_07634_),
    .Y(_08203_));
 AO21x1_ASAP7_75t_R _15227_ (.A1(_08196_),
    .A2(_08199_),
    .B(_08203_),
    .Y(_08204_));
 OR2x2_ASAP7_75t_R _15228_ (.A(_07933_),
    .B(_08204_),
    .Y(_08205_));
 OA21x2_ASAP7_75t_R _15229_ (.A1(_07592_),
    .A2(_08195_),
    .B(_08205_),
    .Y(net44));
 OA21x2_ASAP7_75t_R _15230_ (.A1(_08063_),
    .A2(_08066_),
    .B(_07647_),
    .Y(_08206_));
 AO21x1_ASAP7_75t_R _15231_ (.A1(_07311_),
    .A2(_07884_),
    .B(_08206_),
    .Y(_08207_));
 NAND2x1_ASAP7_75t_R _15232_ (.A(_10004_),
    .B(_07518_),
    .Y(_08208_));
 OA211x2_ASAP7_75t_R _15233_ (.A1(_10014_),
    .A2(_07580_),
    .B(_08208_),
    .C(_07718_),
    .Y(_08209_));
 AOI21x1_ASAP7_75t_R _15234_ (.A1(_07570_),
    .A2(_08185_),
    .B(_08209_),
    .Y(_08210_));
 AOI211x1_ASAP7_75t_R _15235_ (.A1(_03581_),
    .A2(_08130_),
    .B(_08131_),
    .C(_07534_),
    .Y(_08211_));
 AO21x1_ASAP7_75t_R _15236_ (.A1(_07540_),
    .A2(_08210_),
    .B(_08211_),
    .Y(_08212_));
 NOR2x1_ASAP7_75t_R _15237_ (.A(_07722_),
    .B(_07881_),
    .Y(_08213_));
 AO221x1_ASAP7_75t_R _15238_ (.A1(_07728_),
    .A2(_08207_),
    .B1(_08212_),
    .B2(_07749_),
    .C(_08213_),
    .Y(_08214_));
 OA211x2_ASAP7_75t_R _15239_ (.A1(_07346_),
    .A2(_07357_),
    .B(_07398_),
    .C(_07370_),
    .Y(_08215_));
 XNOR2x1_ASAP7_75t_R _15240_ (.B(_08215_),
    .Y(_08216_),
    .A(_00400_));
 NAND2x1_ASAP7_75t_R _15241_ (.A(_01179_),
    .B(_07595_),
    .Y(_08217_));
 OA21x2_ASAP7_75t_R _15242_ (.A1(_01180_),
    .A2(_07424_),
    .B(_08217_),
    .Y(_08218_));
 OA222x2_ASAP7_75t_R _15243_ (.A1(_00400_),
    .A2(_07688_),
    .B1(_07830_),
    .B2(_08216_),
    .C1(_08218_),
    .C2(_07423_),
    .Y(_08219_));
 AND2x2_ASAP7_75t_R _15244_ (.A(_07665_),
    .B(_07881_),
    .Y(_08220_));
 AO21x1_ASAP7_75t_R _15245_ (.A1(_06965_),
    .A2(_07886_),
    .B(_07712_),
    .Y(_08221_));
 OA21x2_ASAP7_75t_R _15246_ (.A1(_08220_),
    .A2(_08221_),
    .B(_07893_),
    .Y(_08222_));
 AO21x1_ASAP7_75t_R _15247_ (.A1(_07872_),
    .A2(_08141_),
    .B(_07336_),
    .Y(_08223_));
 OAI22x1_ASAP7_75t_R _15248_ (.A1(_07643_),
    .A2(_08219_),
    .B1(_08222_),
    .B2(_08223_),
    .Y(_08224_));
 AO21x2_ASAP7_75t_R _15249_ (.A1(_07682_),
    .A2(_08214_),
    .B(_08224_),
    .Y(net45));
 NAND2x1_ASAP7_75t_R _15250_ (.A(_01177_),
    .B(_07777_),
    .Y(_08225_));
 OA21x2_ASAP7_75t_R _15251_ (.A1(_01178_),
    .A2(_07684_),
    .B(_08225_),
    .Y(_08226_));
 OA21x2_ASAP7_75t_R _15252_ (.A1(_07423_),
    .A2(_08226_),
    .B(_07591_),
    .Y(_08227_));
 INVx1_ASAP7_75t_R _15253_ (.A(_00367_),
    .Y(_08228_));
 OR3x1_ASAP7_75t_R _15254_ (.A(_00466_),
    .B(_07610_),
    .C(_07612_),
    .Y(_08229_));
 AO21x1_ASAP7_75t_R _15255_ (.A1(_01183_),
    .A2(_08229_),
    .B(_00433_),
    .Y(_08230_));
 OA211x2_ASAP7_75t_R _15256_ (.A1(_07349_),
    .A2(_07605_),
    .B(_08230_),
    .C(_01181_),
    .Y(_08231_));
 OA21x2_ASAP7_75t_R _15257_ (.A1(_00400_),
    .A2(_08231_),
    .B(_01180_),
    .Y(_08232_));
 AO21x1_ASAP7_75t_R _15258_ (.A1(_07642_),
    .A2(_08232_),
    .B(_07639_),
    .Y(_08233_));
 NAND2x1_ASAP7_75t_R _15259_ (.A(_08228_),
    .B(_08233_),
    .Y(_08234_));
 OR3x1_ASAP7_75t_R _15260_ (.A(_08228_),
    .B(_07830_),
    .C(_08232_),
    .Y(_08235_));
 AO21x1_ASAP7_75t_R _15261_ (.A1(_07894_),
    .A2(_07897_),
    .B(_07244_),
    .Y(_08236_));
 AO32x2_ASAP7_75t_R _15262_ (.A1(_08227_),
    .A2(_08234_),
    .A3(_08235_),
    .B1(_08236_),
    .B2(_08144_),
    .Y(_08237_));
 INVx1_ASAP7_75t_R _15263_ (.A(_08237_),
    .Y(_08238_));
 NAND2x1_ASAP7_75t_R _15264_ (.A(_09999_),
    .B(_07580_),
    .Y(_08239_));
 AND2x2_ASAP7_75t_R _15265_ (.A(_08239_),
    .B(_07767_),
    .Y(_08240_));
 OA211x2_ASAP7_75t_R _15266_ (.A1(_10014_),
    .A2(_07580_),
    .B(_08208_),
    .C(_07671_),
    .Y(_08241_));
 AOI21x1_ASAP7_75t_R _15267_ (.A1(_03581_),
    .A2(_08240_),
    .B(_08241_),
    .Y(_08242_));
 NAND2x1_ASAP7_75t_R _15268_ (.A(_07535_),
    .B(_08242_),
    .Y(_08243_));
 OA21x2_ASAP7_75t_R _15269_ (.A1(_07535_),
    .A2(_08147_),
    .B(_08243_),
    .Y(_08244_));
 OA21x2_ASAP7_75t_R _15270_ (.A1(_08081_),
    .A2(_08084_),
    .B(_07728_),
    .Y(_08245_));
 AOI211x1_ASAP7_75t_R _15271_ (.A1(_07666_),
    .A2(_08244_),
    .B(_08245_),
    .C(_07517_),
    .Y(_08246_));
 AO21x1_ASAP7_75t_R _15272_ (.A1(_07913_),
    .A2(_08104_),
    .B(_07786_),
    .Y(_08247_));
 OR3x4_ASAP7_75t_R _15273_ (.A(_07910_),
    .B(_08246_),
    .C(_08247_),
    .Y(_08248_));
 AND2x4_ASAP7_75t_R _15274_ (.A(_08238_),
    .B(_08248_),
    .Y(net46));
 AND4x2_ASAP7_75t_R _15275_ (.A(_07666_),
    .B(_07517_),
    .C(_07558_),
    .D(_07682_),
    .Y(_08249_));
 NAND2x1_ASAP7_75t_R _15276_ (.A(_01175_),
    .B(_07595_),
    .Y(_08250_));
 OA21x2_ASAP7_75t_R _15277_ (.A1(_01174_),
    .A2(_07684_),
    .B(_08250_),
    .Y(_08251_));
 OA21x2_ASAP7_75t_R _15278_ (.A1(_07423_),
    .A2(_08251_),
    .B(_07336_),
    .Y(_08252_));
 INVx1_ASAP7_75t_R _15279_ (.A(_00300_),
    .Y(_08253_));
 OA21x2_ASAP7_75t_R _15280_ (.A1(_00367_),
    .A2(_08232_),
    .B(_01178_),
    .Y(_08254_));
 OA21x2_ASAP7_75t_R _15281_ (.A1(_00334_),
    .A2(_08254_),
    .B(_00333_),
    .Y(_08255_));
 AO21x1_ASAP7_75t_R _15282_ (.A1(_07642_),
    .A2(_08255_),
    .B(_07639_),
    .Y(_08256_));
 NAND2x1_ASAP7_75t_R _15283_ (.A(_08253_),
    .B(_08256_),
    .Y(_08257_));
 OR3x1_ASAP7_75t_R _15284_ (.A(_08253_),
    .B(_07830_),
    .C(_08255_),
    .Y(_08258_));
 AO21x1_ASAP7_75t_R _15285_ (.A1(_07681_),
    .A2(_07957_),
    .B(_08144_),
    .Y(_08259_));
 AO32x2_ASAP7_75t_R _15286_ (.A1(_08252_),
    .A2(_08257_),
    .A3(_08258_),
    .B1(_08259_),
    .B2(_07517_),
    .Y(_08260_));
 AOI21x1_ASAP7_75t_R _15287_ (.A1(_07081_),
    .A2(_08049_),
    .B(_08110_),
    .Y(_08261_));
 OA211x2_ASAP7_75t_R _15288_ (.A1(_09999_),
    .A2(_07550_),
    .B(_07320_),
    .C(_07673_),
    .Y(_08262_));
 AO31x2_ASAP7_75t_R _15289_ (.A1(_07570_),
    .A2(_07319_),
    .A3(_07446_),
    .B(_08262_),
    .Y(_08263_));
 NOR2x1_ASAP7_75t_R _15290_ (.A(_07578_),
    .B(_08263_),
    .Y(_08264_));
 AOI211x1_ASAP7_75t_R _15291_ (.A1(_07081_),
    .A2(_08187_),
    .B(_08264_),
    .C(_07538_),
    .Y(_08265_));
 AOI21x1_ASAP7_75t_R _15292_ (.A1(_07728_),
    .A2(_08261_),
    .B(_08265_),
    .Y(_08266_));
 AO32x2_ASAP7_75t_R _15293_ (.A1(_07682_),
    .A2(_07958_),
    .A3(_08266_),
    .B1(_08144_),
    .B2(_07952_),
    .Y(_08267_));
 NOR3x2_ASAP7_75t_R _15294_ (.B(_08260_),
    .C(_08267_),
    .Y(net48),
    .A(_08249_));
 NAND2x1_ASAP7_75t_R _15295_ (.A(_07665_),
    .B(_07710_),
    .Y(_08268_));
 OAI21x1_ASAP7_75t_R _15296_ (.A1(_07506_),
    .A2(_07278_),
    .B(_07412_),
    .Y(_08269_));
 AO221x1_ASAP7_75t_R _15297_ (.A1(_07509_),
    .A2(_07721_),
    .B1(_08268_),
    .B2(_07330_),
    .C(_08269_),
    .Y(_08270_));
 AO21x2_ASAP7_75t_R _15298_ (.A1(_04809_),
    .A2(_04847_),
    .B(_07500_),
    .Y(_08271_));
 NAND2x2_ASAP7_75t_R _15299_ (.A(_09994_),
    .B(_07185_),
    .Y(_08272_));
 OA211x2_ASAP7_75t_R _15300_ (.A1(_09999_),
    .A2(_07549_),
    .B(_07320_),
    .C(_07235_),
    .Y(_08273_));
 AO31x2_ASAP7_75t_R _15301_ (.A1(_07673_),
    .A2(_08271_),
    .A3(_08272_),
    .B(_08273_),
    .Y(_08274_));
 OR2x2_ASAP7_75t_R _15302_ (.A(_07079_),
    .B(_08274_),
    .Y(_08275_));
 OA211x2_ASAP7_75t_R _15303_ (.A1(_07534_),
    .A2(_08210_),
    .B(_08275_),
    .C(_07489_),
    .Y(_08276_));
 AO21x1_ASAP7_75t_R _15304_ (.A1(_06965_),
    .A2(_08134_),
    .B(_08276_),
    .Y(_08277_));
 AO21x1_ASAP7_75t_R _15305_ (.A1(_07559_),
    .A2(_07980_),
    .B(_07981_),
    .Y(_08278_));
 OA21x2_ASAP7_75t_R _15306_ (.A1(_07506_),
    .A2(_08278_),
    .B(_07647_),
    .Y(_08279_));
 OA21x2_ASAP7_75t_R _15307_ (.A1(_06866_),
    .A2(_08277_),
    .B(_08279_),
    .Y(_08280_));
 OA21x2_ASAP7_75t_R _15308_ (.A1(_07346_),
    .A2(_07357_),
    .B(_07370_),
    .Y(_08281_));
 OA21x2_ASAP7_75t_R _15309_ (.A1(_08281_),
    .A2(_07388_),
    .B(_07400_),
    .Y(_08282_));
 OA21x2_ASAP7_75t_R _15310_ (.A1(_08282_),
    .A2(_07470_),
    .B(_07474_),
    .Y(_08283_));
 INVx1_ASAP7_75t_R _15311_ (.A(_01173_),
    .Y(_08284_));
 AO22x1_ASAP7_75t_R _15312_ (.A1(_01172_),
    .A2(_07383_),
    .B1(_07409_),
    .B2(_08284_),
    .Y(_08285_));
 NAND2x1_ASAP7_75t_R _15313_ (.A(_07408_),
    .B(_08285_),
    .Y(_08286_));
 AND3x1_ASAP7_75t_R _15314_ (.A(_00267_),
    .B(_07336_),
    .C(_08286_),
    .Y(_08287_));
 OAI21x1_ASAP7_75t_R _15315_ (.A1(_07830_),
    .A2(_08283_),
    .B(_08287_),
    .Y(_08288_));
 INVx1_ASAP7_75t_R _15316_ (.A(_08286_),
    .Y(_08289_));
 OR4x1_ASAP7_75t_R _15317_ (.A(_00267_),
    .B(_07412_),
    .C(_07639_),
    .D(_08289_),
    .Y(_08290_));
 AO21x1_ASAP7_75t_R _15318_ (.A1(_07642_),
    .A2(_08283_),
    .B(_08290_),
    .Y(_08291_));
 OA211x2_ASAP7_75t_R _15319_ (.A1(_08270_),
    .A2(_08280_),
    .B(_08288_),
    .C(_08291_),
    .Y(_08292_));
 BUFx6f_ASAP7_75t_R _15320_ (.A(_08292_),
    .Y(net49));
 OA21x2_ASAP7_75t_R _15321_ (.A1(_07957_),
    .A2(_08010_),
    .B(_07681_),
    .Y(_08293_));
 OA21x2_ASAP7_75t_R _15322_ (.A1(_08144_),
    .A2(_08293_),
    .B(_07517_),
    .Y(_08294_));
 NOR2x1_ASAP7_75t_R _15323_ (.A(_07540_),
    .B(_08242_),
    .Y(_08295_));
 NAND2x1_ASAP7_75t_R _15324_ (.A(_07729_),
    .B(_07497_),
    .Y(_08296_));
 NAND3x2_ASAP7_75t_R _15325_ (.B(_08271_),
    .C(_08272_),
    .Y(_08297_),
    .A(_07579_));
 AND3x1_ASAP7_75t_R _15326_ (.A(_07657_),
    .B(_08296_),
    .C(_08297_),
    .Y(_08298_));
 OR3x1_ASAP7_75t_R _15327_ (.A(_07538_),
    .B(_08295_),
    .C(_08298_),
    .Y(_08299_));
 OA211x2_ASAP7_75t_R _15328_ (.A1(_07666_),
    .A2(_08149_),
    .B(_08293_),
    .C(_08299_),
    .Y(_08300_));
 NAND2x1_ASAP7_75t_R _15329_ (.A(_01170_),
    .B(_07595_),
    .Y(_08301_));
 OA21x2_ASAP7_75t_R _15330_ (.A1(_01171_),
    .A2(_07684_),
    .B(_08301_),
    .Y(_08302_));
 OA21x2_ASAP7_75t_R _15331_ (.A1(_07423_),
    .A2(_08302_),
    .B(_07336_),
    .Y(_08303_));
 INVx1_ASAP7_75t_R _15332_ (.A(_00234_),
    .Y(_08304_));
 OA21x2_ASAP7_75t_R _15333_ (.A1(_07616_),
    .A2(_07617_),
    .B(_01174_),
    .Y(_08305_));
 OA21x2_ASAP7_75t_R _15334_ (.A1(_00267_),
    .A2(_08305_),
    .B(_01173_),
    .Y(_08306_));
 AO21x1_ASAP7_75t_R _15335_ (.A1(_07642_),
    .A2(_08306_),
    .B(_07639_),
    .Y(_08307_));
 NAND2x1_ASAP7_75t_R _15336_ (.A(_08304_),
    .B(_08307_),
    .Y(_08308_));
 OR3x1_ASAP7_75t_R _15337_ (.A(_08304_),
    .B(_07830_),
    .C(_08306_),
    .Y(_08309_));
 AO32x1_ASAP7_75t_R _15338_ (.A1(_08303_),
    .A2(_08308_),
    .A3(_08309_),
    .B1(_08144_),
    .B2(_08004_),
    .Y(_08310_));
 OR3x4_ASAP7_75t_R _15339_ (.A(_08294_),
    .B(_08300_),
    .C(_08310_),
    .Y(_08311_));
 INVx1_ASAP7_75t_R _15340_ (.A(_08311_),
    .Y(net50));
 OR3x1_ASAP7_75t_R _15341_ (.A(_06965_),
    .B(_07814_),
    .C(_07815_),
    .Y(_08312_));
 AOI21x1_ASAP7_75t_R _15342_ (.A1(_07330_),
    .A2(_08312_),
    .B(_08269_),
    .Y(_08313_));
 AND3x1_ASAP7_75t_R _15343_ (.A(_07079_),
    .B(_07319_),
    .C(_07446_),
    .Y(_08314_));
 AOI211x1_ASAP7_75t_R _15344_ (.A1(_07702_),
    .A2(_07495_),
    .B(_08314_),
    .C(_07570_),
    .Y(_08315_));
 AO21x1_ASAP7_75t_R _15345_ (.A1(_09989_),
    .A2(_07552_),
    .B(_07704_),
    .Y(_08316_));
 AO32x1_ASAP7_75t_R _15346_ (.A1(_07314_),
    .A2(_08239_),
    .A3(_07767_),
    .B1(_07263_),
    .B2(_08316_),
    .Y(_08317_));
 OA33x2_ASAP7_75t_R _15347_ (.A1(_08020_),
    .A2(_08175_),
    .A3(_08178_),
    .B1(_08315_),
    .B2(_08317_),
    .B3(_07244_),
    .Y(_08318_));
 OA21x2_ASAP7_75t_R _15348_ (.A1(_08019_),
    .A2(_08020_),
    .B(_06866_),
    .Y(_08319_));
 AO32x1_ASAP7_75t_R _15349_ (.A1(_07506_),
    .A2(_08032_),
    .A3(_08318_),
    .B1(_08319_),
    .B2(_08026_),
    .Y(_08320_));
 OR2x2_ASAP7_75t_R _15350_ (.A(_07388_),
    .B(_07471_),
    .Y(_08321_));
 OA21x2_ASAP7_75t_R _15351_ (.A1(_07400_),
    .A2(_07471_),
    .B(_07476_),
    .Y(_08322_));
 OA21x2_ASAP7_75t_R _15352_ (.A1(_08281_),
    .A2(_08321_),
    .B(_08322_),
    .Y(_08323_));
 INVx1_ASAP7_75t_R _15353_ (.A(_00200_),
    .Y(_08324_));
 AO22x1_ASAP7_75t_R _15354_ (.A1(_01169_),
    .A2(_07383_),
    .B1(_07409_),
    .B2(_08324_),
    .Y(_08325_));
 NAND2x1_ASAP7_75t_R _15355_ (.A(_07408_),
    .B(_08325_),
    .Y(_08326_));
 AND3x1_ASAP7_75t_R _15356_ (.A(_00201_),
    .B(_07336_),
    .C(_08326_),
    .Y(_08327_));
 OA21x2_ASAP7_75t_R _15357_ (.A1(_07830_),
    .A2(_08323_),
    .B(_08327_),
    .Y(_08328_));
 INVx1_ASAP7_75t_R _15358_ (.A(_08326_),
    .Y(_08329_));
 OR4x1_ASAP7_75t_R _15359_ (.A(_00201_),
    .B(_07412_),
    .C(_07639_),
    .D(_08329_),
    .Y(_08330_));
 AOI21x1_ASAP7_75t_R _15360_ (.A1(_07827_),
    .A2(_08323_),
    .B(_08330_),
    .Y(_08331_));
 AOI211x1_ASAP7_75t_R _15361_ (.A1(_08313_),
    .A2(_08320_),
    .B(_08328_),
    .C(_08331_),
    .Y(net51));
 OA21x2_ASAP7_75t_R _15362_ (.A1(_07728_),
    .A2(_07841_),
    .B(_07330_),
    .Y(_08332_));
 NOR2x1_ASAP7_75t_R _15363_ (.A(_08269_),
    .B(_08332_),
    .Y(_08333_));
 NOR2x1_ASAP7_75t_R _15364_ (.A(_07665_),
    .B(_07850_),
    .Y(_08334_));
 AO21x1_ASAP7_75t_R _15365_ (.A1(_07853_),
    .A2(_08051_),
    .B(_08334_),
    .Y(_08335_));
 NAND2x1_ASAP7_75t_R _15366_ (.A(_09977_),
    .B(_07552_),
    .Y(_08336_));
 AO21x1_ASAP7_75t_R _15367_ (.A1(_08336_),
    .A2(_07554_),
    .B(_07570_),
    .Y(_08337_));
 OR3x1_ASAP7_75t_R _15368_ (.A(_07541_),
    .B(_07313_),
    .C(_07494_),
    .Y(_08338_));
 AO32x1_ASAP7_75t_R _15369_ (.A1(_07243_),
    .A2(_08337_),
    .A3(_08338_),
    .B1(_07311_),
    .B2(_07556_),
    .Y(_08339_));
 AND3x1_ASAP7_75t_R _15370_ (.A(_07578_),
    .B(_07647_),
    .C(_08263_),
    .Y(_08340_));
 AO21x1_ASAP7_75t_R _15371_ (.A1(_07540_),
    .A2(_08339_),
    .B(_08340_),
    .Y(_08341_));
 AOI22x1_ASAP7_75t_R _15372_ (.A1(_08129_),
    .A2(_08189_),
    .B1(_08341_),
    .B2(_07853_),
    .Y(_08342_));
 OA22x2_ASAP7_75t_R _15373_ (.A1(_07487_),
    .A2(_08335_),
    .B1(_08342_),
    .B2(_06867_),
    .Y(_08343_));
 OR3x1_ASAP7_75t_R _15374_ (.A(_00201_),
    .B(_07619_),
    .C(_07621_),
    .Y(_08344_));
 AND2x2_ASAP7_75t_R _15375_ (.A(_00200_),
    .B(_08344_),
    .Y(_08345_));
 AOI21x1_ASAP7_75t_R _15376_ (.A1(_07827_),
    .A2(_08345_),
    .B(_07828_),
    .Y(_08346_));
 INVx1_ASAP7_75t_R _15377_ (.A(_00167_),
    .Y(_08347_));
 OR3x1_ASAP7_75t_R _15378_ (.A(_08347_),
    .B(_07430_),
    .C(_08345_),
    .Y(_08348_));
 NAND2x1_ASAP7_75t_R _15379_ (.A(_01167_),
    .B(_07595_),
    .Y(_08349_));
 OA21x2_ASAP7_75t_R _15380_ (.A1(_01168_),
    .A2(_07424_),
    .B(_08349_),
    .Y(_08350_));
 OA21x2_ASAP7_75t_R _15381_ (.A1(_07423_),
    .A2(_08350_),
    .B(_07336_),
    .Y(_08351_));
 OA211x2_ASAP7_75t_R _15382_ (.A1(_00167_),
    .A2(_08346_),
    .B(_08348_),
    .C(_08351_),
    .Y(_08352_));
 AOI21x1_ASAP7_75t_R _15383_ (.A1(_08333_),
    .A2(_08343_),
    .B(_08352_),
    .Y(net52));
 AND3x1_ASAP7_75t_R _15384_ (.A(_00200_),
    .B(_01168_),
    .C(_07386_),
    .Y(_08353_));
 OA21x2_ASAP7_75t_R _15385_ (.A1(_00201_),
    .A2(_08323_),
    .B(_08353_),
    .Y(_08354_));
 AND3x1_ASAP7_75t_R _15386_ (.A(_00167_),
    .B(_01168_),
    .C(_07642_),
    .Y(_08355_));
 INVx1_ASAP7_75t_R _15387_ (.A(_00134_),
    .Y(_08356_));
 OA31x2_ASAP7_75t_R _15388_ (.A1(_07828_),
    .A2(_08354_),
    .A3(_08355_),
    .B1(_08356_),
    .Y(_08357_));
 INVx1_ASAP7_75t_R _15389_ (.A(_00133_),
    .Y(_08358_));
 AO22x1_ASAP7_75t_R _15390_ (.A1(_01166_),
    .A2(_07596_),
    .B1(_07635_),
    .B2(_08358_),
    .Y(_08359_));
 AO21x1_ASAP7_75t_R _15391_ (.A1(_07634_),
    .A2(_08359_),
    .B(_07643_),
    .Y(_08360_));
 OA211x2_ASAP7_75t_R _15392_ (.A1(_00201_),
    .A2(_08323_),
    .B(_01168_),
    .C(_00200_),
    .Y(_08361_));
 AO21x1_ASAP7_75t_R _15393_ (.A1(_00167_),
    .A2(_01168_),
    .B(_07830_),
    .Y(_08362_));
 NOR3x1_ASAP7_75t_R _15394_ (.A(_08356_),
    .B(_08361_),
    .C(_08362_),
    .Y(_08363_));
 OAI21x1_ASAP7_75t_R _15395_ (.A1(_09962_),
    .A2(_07186_),
    .B(_07542_),
    .Y(_08364_));
 AO21x1_ASAP7_75t_R _15396_ (.A1(_08336_),
    .A2(_07554_),
    .B(_07541_),
    .Y(_08365_));
 OA211x2_ASAP7_75t_R _15397_ (.A1(_07579_),
    .A2(_08364_),
    .B(_08365_),
    .C(_07539_),
    .Y(_08366_));
 AO21x1_ASAP7_75t_R _15398_ (.A1(_07578_),
    .A2(_08274_),
    .B(_08366_),
    .Y(_08367_));
 AO221x1_ASAP7_75t_R _15399_ (.A1(_07509_),
    .A2(_07884_),
    .B1(_08059_),
    .B2(_07330_),
    .C(_08269_),
    .Y(_08368_));
 AO221x1_ASAP7_75t_R _15400_ (.A1(_07443_),
    .A2(_08212_),
    .B1(_08367_),
    .B2(_07507_),
    .C(_08368_),
    .Y(_08369_));
 AO21x1_ASAP7_75t_R _15401_ (.A1(_07488_),
    .A2(_08068_),
    .B(_08369_),
    .Y(_08370_));
 OA31x2_ASAP7_75t_R _15402_ (.A1(_08357_),
    .A2(_08360_),
    .A3(_08363_),
    .B1(_08370_),
    .Y(net53));
 AND2x2_ASAP7_75t_R _15403_ (.A(_08296_),
    .B(_08297_),
    .Y(_08371_));
 AO21x1_ASAP7_75t_R _15404_ (.A1(_07503_),
    .A2(_07504_),
    .B(_07570_),
    .Y(_08372_));
 OA211x2_ASAP7_75t_R _15405_ (.A1(_03581_),
    .A2(_08364_),
    .B(_08372_),
    .C(_07534_),
    .Y(_08373_));
 INVx1_ASAP7_75t_R _15406_ (.A(_08373_),
    .Y(_08374_));
 OA211x2_ASAP7_75t_R _15407_ (.A1(_07535_),
    .A2(_08371_),
    .B(_08374_),
    .C(_07853_),
    .Y(_08375_));
 AO21x1_ASAP7_75t_R _15408_ (.A1(_06966_),
    .A2(_08244_),
    .B(_08375_),
    .Y(_08376_));
 AO21x1_ASAP7_75t_R _15409_ (.A1(_08085_),
    .A2(_08086_),
    .B(_07893_),
    .Y(_08377_));
 AO21x1_ASAP7_75t_R _15410_ (.A1(_07509_),
    .A2(_07908_),
    .B(_07330_),
    .Y(_08378_));
 OA21x2_ASAP7_75t_R _15411_ (.A1(_07908_),
    .A2(_08058_),
    .B(_08378_),
    .Y(_08379_));
 NOR2x1_ASAP7_75t_R _15412_ (.A(_08269_),
    .B(_08379_),
    .Y(_08380_));
 OA211x2_ASAP7_75t_R _15413_ (.A1(_06867_),
    .A2(_08376_),
    .B(_08377_),
    .C(_08380_),
    .Y(_08381_));
 NAND2x1_ASAP7_75t_R _15414_ (.A(_01165_),
    .B(_07596_),
    .Y(_08382_));
 OR3x1_ASAP7_75t_R _15415_ (.A(_00099_),
    .B(_07596_),
    .C(_07828_),
    .Y(_08383_));
 AO21x1_ASAP7_75t_R _15416_ (.A1(_08382_),
    .A2(_08383_),
    .B(_07594_),
    .Y(_08384_));
 AO21x1_ASAP7_75t_R _15417_ (.A1(_00133_),
    .A2(_07625_),
    .B(_07687_),
    .Y(_08385_));
 AOI211x1_ASAP7_75t_R _15418_ (.A1(_07827_),
    .A2(_07626_),
    .B(_00100_),
    .C(_07828_),
    .Y(_08386_));
 AO21x1_ASAP7_75t_R _15419_ (.A1(_00100_),
    .A2(_08385_),
    .B(_08386_),
    .Y(_08387_));
 AO32x2_ASAP7_75t_R _15420_ (.A1(_07592_),
    .A2(_08384_),
    .A3(_08387_),
    .B1(_08380_),
    .B2(_07517_),
    .Y(_08388_));
 NOR2x2_ASAP7_75t_R _15421_ (.A(_08381_),
    .B(_08388_),
    .Y(net55));
 CKINVDCx20_ASAP7_75t_R _15422_ (.A(net31),
    .Y(_01219_));
 INVx1_ASAP7_75t_R _15423_ (.A(net26),
    .Y(_08389_));
 OA21x2_ASAP7_75t_R _15424_ (.A1(_04072_),
    .A2(_08389_),
    .B(_03566_),
    .Y(_08390_));
 AO21x1_ASAP7_75t_R _15425_ (.A1(_04849_),
    .A2(_08390_),
    .B(_05346_),
    .Y(_08391_));
 BUFx6f_ASAP7_75t_R _15426_ (.A(_08391_),
    .Y(_08392_));
 BUFx4f_ASAP7_75t_R _15427_ (.A(_08392_),
    .Y(_08393_));
 NAND2x2_ASAP7_75t_R _15428_ (.A(_04165_),
    .B(_08390_),
    .Y(_08394_));
 AND2x6_ASAP7_75t_R _15429_ (.A(_04174_),
    .B(_08394_),
    .Y(_08395_));
 AND3x1_ASAP7_75t_R _15430_ (.A(_03602_),
    .B(_03770_),
    .C(_08395_),
    .Y(_08396_));
 AO21x1_ASAP7_75t_R _15431_ (.A1(net65),
    .A2(_08393_),
    .B(_08396_),
    .Y(_10105_));
 AND3x1_ASAP7_75t_R _15432_ (.A(_07190_),
    .B(_07233_),
    .C(_08395_),
    .Y(_08397_));
 AO21x2_ASAP7_75t_R _15433_ (.A1(net76),
    .A2(_08393_),
    .B(_08397_),
    .Y(_09944_));
 BUFx4f_ASAP7_75t_R _15434_ (.A(_08392_),
    .Y(_08398_));
 BUFx6f_ASAP7_75t_R _15435_ (.A(_08392_),
    .Y(_08399_));
 NAND2x1_ASAP7_75t_R _15436_ (.A(_10109_),
    .B(_08399_),
    .Y(_08400_));
 OA21x2_ASAP7_75t_R _15437_ (.A1(_10092_),
    .A2(_08398_),
    .B(_08400_),
    .Y(_10107_));
 NAND2x1_ASAP7_75t_R _15438_ (.A(_10110_),
    .B(_08399_),
    .Y(_08401_));
 OA21x2_ASAP7_75t_R _15439_ (.A1(_10087_),
    .A2(_08398_),
    .B(_08401_),
    .Y(_10113_));
 NAND2x1_ASAP7_75t_R _15440_ (.A(_10084_),
    .B(_08395_),
    .Y(_08402_));
 OA21x2_ASAP7_75t_R _15441_ (.A1(net91),
    .A2(_08395_),
    .B(_08402_),
    .Y(_10115_));
 NAND2x1_ASAP7_75t_R _15442_ (.A(_01080_),
    .B(_08399_),
    .Y(_08403_));
 OA21x2_ASAP7_75t_R _15443_ (.A1(_10077_),
    .A2(_08398_),
    .B(_08403_),
    .Y(_10117_));
 BUFx6f_ASAP7_75t_R _15444_ (.A(_08392_),
    .Y(_08404_));
 NAND2x1_ASAP7_75t_R _15445_ (.A(_03479_),
    .B(_08404_),
    .Y(_08405_));
 OA21x2_ASAP7_75t_R _15446_ (.A1(_10072_),
    .A2(_08398_),
    .B(_08405_),
    .Y(_10119_));
 NAND2x1_ASAP7_75t_R _15447_ (.A(_01086_),
    .B(_08404_),
    .Y(_08406_));
 OA21x2_ASAP7_75t_R _15448_ (.A1(_10067_),
    .A2(_08398_),
    .B(_08406_),
    .Y(_10121_));
 BUFx6f_ASAP7_75t_R _15449_ (.A(_08392_),
    .Y(_08407_));
 NOR2x1_ASAP7_75t_R _15450_ (.A(_10064_),
    .B(_08407_),
    .Y(_08408_));
 AO21x1_ASAP7_75t_R _15451_ (.A1(net95),
    .A2(_08399_),
    .B(_08408_),
    .Y(_10123_));
 NOR2x1_ASAP7_75t_R _15452_ (.A(_10059_),
    .B(_08407_),
    .Y(_08409_));
 AO21x1_ASAP7_75t_R _15453_ (.A1(net96),
    .A2(_08399_),
    .B(_08409_),
    .Y(_10125_));
 NOR2x1_ASAP7_75t_R _15454_ (.A(_10102_),
    .B(_08407_),
    .Y(_08410_));
 AO21x1_ASAP7_75t_R _15455_ (.A1(net66),
    .A2(_08399_),
    .B(_08410_),
    .Y(_10127_));
 NOR2x1_ASAP7_75t_R _15456_ (.A(_10054_),
    .B(_08407_),
    .Y(_08411_));
 AO21x1_ASAP7_75t_R _15457_ (.A1(net67),
    .A2(_08399_),
    .B(_08411_),
    .Y(_10129_));
 NAND2x1_ASAP7_75t_R _15458_ (.A(_01101_),
    .B(_08404_),
    .Y(_08412_));
 OA21x2_ASAP7_75t_R _15459_ (.A1(_10047_),
    .A2(_08398_),
    .B(_08412_),
    .Y(_10131_));
 NAND2x1_ASAP7_75t_R _15460_ (.A(_01104_),
    .B(_08404_),
    .Y(_08413_));
 OA21x2_ASAP7_75t_R _15461_ (.A1(_10042_),
    .A2(_08398_),
    .B(_08413_),
    .Y(_10133_));
 NAND2x1_ASAP7_75t_R _15462_ (.A(_01107_),
    .B(_08404_),
    .Y(_08414_));
 OA21x2_ASAP7_75t_R _15463_ (.A1(_10037_),
    .A2(_08398_),
    .B(_08414_),
    .Y(_10135_));
 NOR2x1_ASAP7_75t_R _15464_ (.A(_10034_),
    .B(_08407_),
    .Y(_08415_));
 AO21x1_ASAP7_75t_R _15465_ (.A1(net71),
    .A2(_08399_),
    .B(_08415_),
    .Y(_10137_));
 NAND2x1_ASAP7_75t_R _15466_ (.A(_01113_),
    .B(_08404_),
    .Y(_08416_));
 OA21x2_ASAP7_75t_R _15467_ (.A1(_10027_),
    .A2(_08398_),
    .B(_08416_),
    .Y(_10139_));
 NAND2x1_ASAP7_75t_R _15468_ (.A(_10024_),
    .B(_08395_),
    .Y(_08417_));
 OA21x2_ASAP7_75t_R _15469_ (.A1(net73),
    .A2(_08395_),
    .B(_08417_),
    .Y(_10141_));
 NOR2x1_ASAP7_75t_R _15470_ (.A(_10019_),
    .B(_08392_),
    .Y(_08418_));
 AO21x1_ASAP7_75t_R _15471_ (.A1(net74),
    .A2(_08399_),
    .B(_08418_),
    .Y(_10143_));
 NAND2x1_ASAP7_75t_R _15472_ (.A(_01122_),
    .B(_08404_),
    .Y(_08419_));
 OA21x2_ASAP7_75t_R _15473_ (.A1(_10012_),
    .A2(_08398_),
    .B(_08419_),
    .Y(_10145_));
 AND2x2_ASAP7_75t_R _15474_ (.A(net77),
    .B(_08392_),
    .Y(_08420_));
 AO21x1_ASAP7_75t_R _15475_ (.A1(_10007_),
    .A2(_08395_),
    .B(_08420_),
    .Y(_10147_));
 NAND2x1_ASAP7_75t_R _15476_ (.A(_01128_),
    .B(_08404_),
    .Y(_08421_));
 OA21x2_ASAP7_75t_R _15477_ (.A1(_10004_),
    .A2(_08393_),
    .B(_08421_),
    .Y(_10149_));
 NAND2x1_ASAP7_75t_R _15478_ (.A(_01131_),
    .B(_08404_),
    .Y(_08422_));
 OA21x2_ASAP7_75t_R _15479_ (.A1(_09999_),
    .A2(_08393_),
    .B(_08422_),
    .Y(_10151_));
 NAND2x1_ASAP7_75t_R _15480_ (.A(_01134_),
    .B(_08404_),
    .Y(_08423_));
 OA21x2_ASAP7_75t_R _15481_ (.A1(_09992_),
    .A2(_08393_),
    .B(_08423_),
    .Y(_10153_));
 NAND2x1_ASAP7_75t_R _15482_ (.A(_01137_),
    .B(_08407_),
    .Y(_08424_));
 OA21x2_ASAP7_75t_R _15483_ (.A1(_09987_),
    .A2(_08393_),
    .B(_08424_),
    .Y(_10155_));
 AND3x1_ASAP7_75t_R _15484_ (.A(_04809_),
    .B(_04847_),
    .C(_08395_),
    .Y(_08425_));
 AO21x1_ASAP7_75t_R _15485_ (.A1(net82),
    .A2(_08399_),
    .B(_08425_),
    .Y(_10157_));
 NAND2x1_ASAP7_75t_R _15486_ (.A(_01143_),
    .B(_08407_),
    .Y(_08426_));
 OA21x2_ASAP7_75t_R _15487_ (.A1(_09979_),
    .A2(_08393_),
    .B(_08426_),
    .Y(_10159_));
 AND2x2_ASAP7_75t_R _15488_ (.A(net84),
    .B(_08392_),
    .Y(_08427_));
 AO21x1_ASAP7_75t_R _15489_ (.A1(_09974_),
    .A2(_08395_),
    .B(_08427_),
    .Y(_10161_));
 NAND2x1_ASAP7_75t_R _15490_ (.A(_01149_),
    .B(_08407_),
    .Y(_08428_));
 OA21x2_ASAP7_75t_R _15491_ (.A1(_09969_),
    .A2(_08393_),
    .B(_08428_),
    .Y(_10163_));
 NAND2x1_ASAP7_75t_R _15492_ (.A(_01152_),
    .B(_08407_),
    .Y(_08429_));
 OA21x2_ASAP7_75t_R _15493_ (.A1(_09964_),
    .A2(_08393_),
    .B(_08429_),
    .Y(_10165_));
 NAND2x1_ASAP7_75t_R _15494_ (.A(_01155_),
    .B(_08407_),
    .Y(_08430_));
 OA21x2_ASAP7_75t_R _15495_ (.A1(_09959_),
    .A2(_08393_),
    .B(_08430_),
    .Y(_10167_));
 AND2x2_ASAP7_75t_R _15496_ (.A(_04253_),
    .B(_05301_),
    .Y(_10148_));
 AND3x2_ASAP7_75t_R _15497_ (.A(_03497_),
    .B(_03503_),
    .C(_05853_),
    .Y(_08431_));
 XNOR2x2_ASAP7_75t_R _15498_ (.A(_04056_),
    .B(_08431_),
    .Y(_08432_));
 XNOR2x2_ASAP7_75t_R _15499_ (.A(_09955_),
    .B(_08431_),
    .Y(_08433_));
 NAND2x1_ASAP7_75t_R _15500_ (.A(_08432_),
    .B(_08433_),
    .Y(_08434_));
 OAI21x1_ASAP7_75t_R _15501_ (.A1(_04123_),
    .A2(_04160_),
    .B(_03447_),
    .Y(_08435_));
 AO221x1_ASAP7_75t_R _15502_ (.A1(_04453_),
    .A2(_04469_),
    .B1(_04484_),
    .B2(_04500_),
    .C(_04431_),
    .Y(_08436_));
 MAJx2_ASAP7_75t_R _15503_ (.A(_04320_),
    .B(_09964_),
    .C(_08436_),
    .Y(_08437_));
 MAJx2_ASAP7_75t_R _15504_ (.A(_08435_),
    .B(_09959_),
    .C(_08437_),
    .Y(_08438_));
 AO32x1_ASAP7_75t_R _15505_ (.A1(_04784_),
    .A2(_04809_),
    .A3(_04847_),
    .B1(_04895_),
    .B2(_09987_),
    .Y(_08439_));
 AO21x1_ASAP7_75t_R _15506_ (.A1(_04809_),
    .A2(_04847_),
    .B(_04784_),
    .Y(_08440_));
 OAI21x1_ASAP7_75t_R _15507_ (.A1(_04655_),
    .A2(_04682_),
    .B(_03447_),
    .Y(_08441_));
 AND2x2_ASAP7_75t_R _15508_ (.A(_08441_),
    .B(_09979_),
    .Y(_08442_));
 AO221x1_ASAP7_75t_R _15509_ (.A1(_04566_),
    .A2(_09974_),
    .B1(_08439_),
    .B2(_08440_),
    .C(_08442_),
    .Y(_08443_));
 NAND2x1_ASAP7_75t_R _15510_ (.A(_04683_),
    .B(_09977_),
    .Y(_08444_));
 MAJx2_ASAP7_75t_R _15511_ (.A(_04566_),
    .B(_09974_),
    .C(_08444_),
    .Y(_08445_));
 AND4x1_ASAP7_75t_R _15512_ (.A(_08434_),
    .B(_08438_),
    .C(_08443_),
    .D(_08445_),
    .Y(_08446_));
 AO21x1_ASAP7_75t_R _15513_ (.A1(_04431_),
    .A2(_09969_),
    .B(_09964_),
    .Y(_08447_));
 AND3x1_ASAP7_75t_R _15514_ (.A(_09964_),
    .B(_04431_),
    .C(_09969_),
    .Y(_08448_));
 AO221x1_ASAP7_75t_R _15515_ (.A1(_08435_),
    .A2(_09959_),
    .B1(_04320_),
    .B2(_08447_),
    .C(_08448_),
    .Y(_08449_));
 AOI22x1_ASAP7_75t_R _15516_ (.A1(_04161_),
    .A2(_09957_),
    .B1(_08432_),
    .B2(_08433_),
    .Y(_08450_));
 NOR2x1_ASAP7_75t_R _15517_ (.A(_08432_),
    .B(_08433_),
    .Y(_08451_));
 AO21x1_ASAP7_75t_R _15518_ (.A1(_08449_),
    .A2(_08450_),
    .B(_08451_),
    .Y(_08452_));
 AOI211x1_ASAP7_75t_R _15519_ (.A1(_05014_),
    .A2(_09992_),
    .B(_08446_),
    .C(_08452_),
    .Y(_08453_));
 INVx1_ASAP7_75t_R _15520_ (.A(_05209_),
    .Y(_08454_));
 AOI22x1_ASAP7_75t_R _15521_ (.A1(_05104_),
    .A2(_09999_),
    .B1(_08454_),
    .B2(_10004_),
    .Y(_08455_));
 AO22x1_ASAP7_75t_R _15522_ (.A1(_05209_),
    .A2(_10002_),
    .B1(_05300_),
    .B2(_10009_),
    .Y(_08456_));
 OAI22x1_ASAP7_75t_R _15523_ (.A1(_05014_),
    .A2(_09992_),
    .B1(_05104_),
    .B2(_09999_),
    .Y(_08457_));
 AO21x1_ASAP7_75t_R _15524_ (.A1(_08455_),
    .A2(_08456_),
    .B(_08457_),
    .Y(_08458_));
 NAND2x1_ASAP7_75t_R _15525_ (.A(_05694_),
    .B(_10027_),
    .Y(_08459_));
 MAJx2_ASAP7_75t_R _15526_ (.A(_05596_),
    .B(_10024_),
    .C(_08459_),
    .Y(_08460_));
 OR3x1_ASAP7_75t_R _15527_ (.A(_05494_),
    .B(_05529_),
    .C(_05545_),
    .Y(_08461_));
 OA211x2_ASAP7_75t_R _15528_ (.A1(_05396_),
    .A2(_10014_),
    .B(_08460_),
    .C(_08461_),
    .Y(_08462_));
 OA21x2_ASAP7_75t_R _15529_ (.A1(_05529_),
    .A2(_05545_),
    .B(_05494_),
    .Y(_08463_));
 MAJx2_ASAP7_75t_R _15530_ (.A(_05396_),
    .B(_10014_),
    .C(_08463_),
    .Y(_08464_));
 OR4x1_ASAP7_75t_R _15531_ (.A(_10002_),
    .B(_05300_),
    .C(_05342_),
    .D(_05345_),
    .Y(_08465_));
 OR4x1_ASAP7_75t_R _15532_ (.A(_05209_),
    .B(_05300_),
    .C(_05342_),
    .D(_05345_),
    .Y(_08466_));
 AO31x2_ASAP7_75t_R _15533_ (.A1(_08465_),
    .A2(_08466_),
    .A3(_08455_),
    .B(_08457_),
    .Y(_08467_));
 OA31x2_ASAP7_75t_R _15534_ (.A1(_08458_),
    .A2(_08462_),
    .A3(_08464_),
    .B1(_08467_),
    .Y(_08468_));
 AND2x2_ASAP7_75t_R _15535_ (.A(_08453_),
    .B(_08468_),
    .Y(_08469_));
 OA211x2_ASAP7_75t_R _15536_ (.A1(_04895_),
    .A2(_09987_),
    .B(_04809_),
    .C(_04847_),
    .Y(_08470_));
 OA21x2_ASAP7_75t_R _15537_ (.A1(_04895_),
    .A2(_09987_),
    .B(_04784_),
    .Y(_08471_));
 AO32x1_ASAP7_75t_R _15538_ (.A1(_04784_),
    .A2(_04809_),
    .A3(_04847_),
    .B1(_09979_),
    .B2(_08441_),
    .Y(_08472_));
 OA31x2_ASAP7_75t_R _15539_ (.A1(_08470_),
    .A2(_08471_),
    .A3(_08472_),
    .B1(_08444_),
    .Y(_08473_));
 MAJx2_ASAP7_75t_R _15540_ (.A(_04566_),
    .B(_09974_),
    .C(_08473_),
    .Y(_08474_));
 AO21x1_ASAP7_75t_R _15541_ (.A1(_08434_),
    .A2(_08438_),
    .B(_08451_),
    .Y(_08475_));
 OAI21x1_ASAP7_75t_R _15542_ (.A1(_08452_),
    .A2(_08474_),
    .B(_08475_),
    .Y(_08476_));
 AOI221x1_ASAP7_75t_R _15543_ (.A1(_05715_),
    .A2(_05725_),
    .B1(_05741_),
    .B2(_05753_),
    .C(_05694_),
    .Y(_08477_));
 MAJx2_ASAP7_75t_R _15544_ (.A(_05596_),
    .B(_10024_),
    .C(_08477_),
    .Y(_08478_));
 OA211x2_ASAP7_75t_R _15545_ (.A1(_05396_),
    .A2(_10014_),
    .B(_08461_),
    .C(_08478_),
    .Y(_08479_));
 OA21x2_ASAP7_75t_R _15546_ (.A1(_08464_),
    .A2(_08479_),
    .B(_08467_),
    .Y(_08480_));
 NAND2x1_ASAP7_75t_R _15547_ (.A(_05014_),
    .B(_09992_),
    .Y(_08481_));
 OA21x2_ASAP7_75t_R _15548_ (.A1(_08458_),
    .A2(_08480_),
    .B(_08481_),
    .Y(_08482_));
 NOR2x1_ASAP7_75t_R _15549_ (.A(_08476_),
    .B(_08482_),
    .Y(_08483_));
 OA21x2_ASAP7_75t_R _15550_ (.A1(net128),
    .A2(_10069_),
    .B(_10074_),
    .Y(_08484_));
 NAND3x1_ASAP7_75t_R _15551_ (.A(_06863_),
    .B(_06878_),
    .C(_06888_),
    .Y(_08485_));
 NAND3x1_ASAP7_75t_R _15552_ (.A(_06863_),
    .B(_06898_),
    .C(_06908_),
    .Y(_08486_));
 AO31x2_ASAP7_75t_R _15553_ (.A1(_10079_),
    .A2(_08485_),
    .A3(_08486_),
    .B(net126),
    .Y(_08487_));
 OR3x1_ASAP7_75t_R _15554_ (.A(_10079_),
    .B(net125),
    .C(_10084_),
    .Y(_08488_));
 MAJx2_ASAP7_75t_R _15555_ (.A(net128),
    .B(_10069_),
    .C(net127),
    .Y(_08489_));
 AO31x2_ASAP7_75t_R _15556_ (.A1(_08484_),
    .A2(_08487_),
    .A3(_08488_),
    .B(_08489_),
    .Y(_08490_));
 AO221x1_ASAP7_75t_R _15557_ (.A1(net128),
    .A2(_10069_),
    .B1(_08487_),
    .B2(_08488_),
    .C(_10074_),
    .Y(_08491_));
 NAND2x1_ASAP7_75t_R _15558_ (.A(_08490_),
    .B(_08491_),
    .Y(_08492_));
 OR2x2_ASAP7_75t_R _15559_ (.A(_06961_),
    .B(_10087_),
    .Y(_08493_));
 AND2x2_ASAP7_75t_R _15560_ (.A(_07179_),
    .B(_07190_),
    .Y(_08494_));
 AO221x2_ASAP7_75t_R _15561_ (.A1(_07200_),
    .A2(_07215_),
    .B1(_07232_),
    .B2(_07190_),
    .C(_07179_),
    .Y(_08495_));
 AO21x1_ASAP7_75t_R _15562_ (.A1(_03602_),
    .A2(_03770_),
    .B(_03478_),
    .Y(_08496_));
 AO21x1_ASAP7_75t_R _15563_ (.A1(_07075_),
    .A2(_10092_),
    .B(_10087_),
    .Y(_08497_));
 AO21x1_ASAP7_75t_R _15564_ (.A1(_07075_),
    .A2(_10092_),
    .B(_06961_),
    .Y(_08498_));
 AO222x2_ASAP7_75t_R _15565_ (.A1(_07233_),
    .A2(_08494_),
    .B1(_08495_),
    .B2(_08496_),
    .C1(_08497_),
    .C2(_08498_),
    .Y(_08499_));
 AND2x2_ASAP7_75t_R _15566_ (.A(_07092_),
    .B(_07099_),
    .Y(_08500_));
 AO211x2_ASAP7_75t_R _15567_ (.A1(_08500_),
    .A2(_07104_),
    .B(_07127_),
    .C(_07075_),
    .Y(_08501_));
 AO21x1_ASAP7_75t_R _15568_ (.A1(_06961_),
    .A2(_10087_),
    .B(_08501_),
    .Y(_08502_));
 AND3x1_ASAP7_75t_R _15569_ (.A(_08493_),
    .B(_08499_),
    .C(_08502_),
    .Y(_08503_));
 NAND2x1_ASAP7_75t_R _15570_ (.A(net128),
    .B(_10069_),
    .Y(_08504_));
 AO221x1_ASAP7_75t_R _15571_ (.A1(_06878_),
    .A2(_06888_),
    .B1(_06898_),
    .B2(_06908_),
    .C(_06863_),
    .Y(_08505_));
 MAJx2_ASAP7_75t_R _15572_ (.A(_06761_),
    .B(_10077_),
    .C(_08505_),
    .Y(_08506_));
 AO211x2_ASAP7_75t_R _15573_ (.A1(_06572_),
    .A2(_10067_),
    .B(_06669_),
    .C(_10072_),
    .Y(_08507_));
 MAJx2_ASAP7_75t_R _15574_ (.A(_06572_),
    .B(_10067_),
    .C(_06669_),
    .Y(_08508_));
 AO21x1_ASAP7_75t_R _15575_ (.A1(_06572_),
    .A2(_10067_),
    .B(_10072_),
    .Y(_08509_));
 AO32x1_ASAP7_75t_R _15576_ (.A1(_08504_),
    .A2(_08506_),
    .A3(_08507_),
    .B1(_08508_),
    .B2(_08509_),
    .Y(_08510_));
 OA21x2_ASAP7_75t_R _15577_ (.A1(_08492_),
    .A2(_08503_),
    .B(_08510_),
    .Y(_08511_));
 AND5x1_ASAP7_75t_R _15578_ (.A(_03478_),
    .B(_03602_),
    .C(_03770_),
    .D(_10092_),
    .E(_08495_),
    .Y(_08512_));
 AND5x1_ASAP7_75t_R _15579_ (.A(_03478_),
    .B(_03602_),
    .C(_03770_),
    .D(_07075_),
    .E(_08495_),
    .Y(_08513_));
 OA211x2_ASAP7_75t_R _15580_ (.A1(_07075_),
    .A2(_10092_),
    .B(_07233_),
    .C(_08494_),
    .Y(_08514_));
 AO22x1_ASAP7_75t_R _15581_ (.A1(_06961_),
    .A2(_10087_),
    .B1(_07075_),
    .B2(_10092_),
    .Y(_08515_));
 OR4x1_ASAP7_75t_R _15582_ (.A(_08512_),
    .B(_08513_),
    .C(_08514_),
    .D(_08515_),
    .Y(_08516_));
 NAND3x1_ASAP7_75t_R _15583_ (.A(_08516_),
    .B(_08510_),
    .C(_08493_),
    .Y(_08517_));
 OA31x2_ASAP7_75t_R _15584_ (.A1(_10059_),
    .A2(_06472_),
    .A3(_10064_),
    .B1(_06377_),
    .Y(_08518_));
 OA21x2_ASAP7_75t_R _15585_ (.A1(_06472_),
    .A2(_10064_),
    .B(_10059_),
    .Y(_08519_));
 OR3x1_ASAP7_75t_R _15586_ (.A(_06284_),
    .B(_08518_),
    .C(_08519_),
    .Y(_08520_));
 OA33x2_ASAP7_75t_R _15587_ (.A1(_06186_),
    .A2(_06207_),
    .A3(_06238_),
    .B1(_06284_),
    .B2(_06290_),
    .B3(_06331_),
    .Y(_08521_));
 OA31x2_ASAP7_75t_R _15588_ (.A1(_10102_),
    .A2(_08518_),
    .A3(_08519_),
    .B1(_08521_),
    .Y(_08522_));
 AND2x2_ASAP7_75t_R _15589_ (.A(_06186_),
    .B(_10054_),
    .Y(_08523_));
 AO21x1_ASAP7_75t_R _15590_ (.A1(_08520_),
    .A2(_08522_),
    .B(_08523_),
    .Y(_08524_));
 XOR2x1_ASAP7_75t_R _15591_ (.A(_05900_),
    .Y(_08525_),
    .B(_10037_));
 XNOR2x1_ASAP7_75t_R _15592_ (.B(_10034_),
    .Y(_08526_),
    .A(_05803_));
 OR2x2_ASAP7_75t_R _15593_ (.A(_06081_),
    .B(_10047_),
    .Y(_08527_));
 MAJx2_ASAP7_75t_R _15594_ (.A(_05995_),
    .B(_10042_),
    .C(_08527_),
    .Y(_08528_));
 OA21x2_ASAP7_75t_R _15595_ (.A1(_05971_),
    .A2(_05994_),
    .B(_03447_),
    .Y(_08529_));
 NAND2x1_ASAP7_75t_R _15596_ (.A(_06081_),
    .B(_10047_),
    .Y(_08530_));
 MAJx2_ASAP7_75t_R _15597_ (.A(_08529_),
    .B(_10044_),
    .C(_08530_),
    .Y(_08531_));
 AND4x1_ASAP7_75t_R _15598_ (.A(_08525_),
    .B(_08526_),
    .C(_08528_),
    .D(_08531_),
    .Y(_08532_));
 AND2x2_ASAP7_75t_R _15599_ (.A(_08490_),
    .B(_08491_),
    .Y(_08533_));
 INVx1_ASAP7_75t_R _15600_ (.A(_06186_),
    .Y(_08534_));
 NOR2x1_ASAP7_75t_R _15601_ (.A(_06377_),
    .B(_10059_),
    .Y(_08535_));
 AOI21x1_ASAP7_75t_R _15602_ (.A1(_07301_),
    .A2(_07302_),
    .B(_06284_),
    .Y(_08536_));
 AOI22x1_ASAP7_75t_R _15603_ (.A1(_06377_),
    .A2(_10059_),
    .B1(_06472_),
    .B2(_10064_),
    .Y(_08537_));
 OAI21x1_ASAP7_75t_R _15604_ (.A1(_06290_),
    .A2(_06331_),
    .B(_06284_),
    .Y(_08538_));
 OA31x2_ASAP7_75t_R _15605_ (.A1(_08535_),
    .A2(_08536_),
    .A3(_08537_),
    .B1(_08538_),
    .Y(_08539_));
 MAJx2_ASAP7_75t_R _15606_ (.A(_08534_),
    .B(_10052_),
    .C(_08539_),
    .Y(_08540_));
 AND5x1_ASAP7_75t_R _15607_ (.A(_08517_),
    .B(_08524_),
    .C(_08532_),
    .D(_08533_),
    .E(_08540_),
    .Y(_08541_));
 AND2x2_ASAP7_75t_R _15608_ (.A(_08511_),
    .B(_08541_),
    .Y(_08542_));
 OR3x1_ASAP7_75t_R _15609_ (.A(_03528_),
    .B(_03483_),
    .C(_05945_),
    .Y(_08543_));
 AO31x2_ASAP7_75t_R _15610_ (.A1(_08469_),
    .A2(_08483_),
    .A3(_08542_),
    .B(_08543_),
    .Y(_08544_));
 NAND2x2_ASAP7_75t_R _15611_ (.A(_08453_),
    .B(_08468_),
    .Y(_08545_));
 NAND2x1_ASAP7_75t_R _15612_ (.A(_08511_),
    .B(_08541_),
    .Y(_08546_));
 OR3x1_ASAP7_75t_R _15613_ (.A(_03528_),
    .B(_03483_),
    .C(_03534_),
    .Y(_08547_));
 AND2x2_ASAP7_75t_R _15614_ (.A(_03382_),
    .B(_08547_),
    .Y(_08548_));
 OR5x1_ASAP7_75t_R _15615_ (.A(_08545_),
    .B(_08476_),
    .C(_08482_),
    .D(_08546_),
    .E(_08548_),
    .Y(_08549_));
 AO21x2_ASAP7_75t_R _15616_ (.A1(_08544_),
    .A2(_08549_),
    .B(_03504_),
    .Y(_08550_));
 AOI21x1_ASAP7_75t_R _15617_ (.A1(_08520_),
    .A2(_08522_),
    .B(_08523_),
    .Y(_08551_));
 AND2x2_ASAP7_75t_R _15618_ (.A(_05803_),
    .B(_10032_),
    .Y(_08552_));
 AND2x2_ASAP7_75t_R _15619_ (.A(_06081_),
    .B(_10047_),
    .Y(_08553_));
 MAJx2_ASAP7_75t_R _15620_ (.A(_05995_),
    .B(_10042_),
    .C(_08553_),
    .Y(_08554_));
 MAJx2_ASAP7_75t_R _15621_ (.A(_05900_),
    .B(_10037_),
    .C(_08554_),
    .Y(_08555_));
 OR3x1_ASAP7_75t_R _15622_ (.A(_08551_),
    .B(_08552_),
    .C(_08555_),
    .Y(_08556_));
 OR3x1_ASAP7_75t_R _15623_ (.A(_08552_),
    .B(_08540_),
    .C(_08555_),
    .Y(_08557_));
 MAJx2_ASAP7_75t_R _15624_ (.A(_05900_),
    .B(_10037_),
    .C(_08528_),
    .Y(_08558_));
 MAJx2_ASAP7_75t_R _15625_ (.A(_05803_),
    .B(_10032_),
    .C(_08558_),
    .Y(_08559_));
 OA211x2_ASAP7_75t_R _15626_ (.A1(_08511_),
    .A2(_08556_),
    .B(_08557_),
    .C(_08559_),
    .Y(_08560_));
 OR2x2_ASAP7_75t_R _15627_ (.A(_08458_),
    .B(_08480_),
    .Y(_08561_));
 AOI21x1_ASAP7_75t_R _15628_ (.A1(_08453_),
    .A2(_08561_),
    .B(_08476_),
    .Y(_08562_));
 OAI21x1_ASAP7_75t_R _15629_ (.A1(_08545_),
    .A2(_08560_),
    .B(_08562_),
    .Y(_08563_));
 OR3x1_ASAP7_75t_R _15630_ (.A(_03534_),
    .B(_03504_),
    .C(_07239_),
    .Y(_08564_));
 INVx1_ASAP7_75t_R _15631_ (.A(_08564_),
    .Y(_08565_));
 AND3x1_ASAP7_75t_R _15632_ (.A(_03534_),
    .B(_06139_),
    .C(_05755_),
    .Y(_08566_));
 OA211x2_ASAP7_75t_R _15633_ (.A1(_08545_),
    .A2(_08560_),
    .B(_08562_),
    .C(_08566_),
    .Y(_08567_));
 NAND2x1_ASAP7_75t_R _15634_ (.A(_03502_),
    .B(_03678_),
    .Y(_08568_));
 AOI21x1_ASAP7_75t_R _15635_ (.A1(_03570_),
    .A2(_03571_),
    .B(_08568_),
    .Y(_08569_));
 BUFx6f_ASAP7_75t_R _15636_ (.A(_08569_),
    .Y(_08570_));
 AOI211x1_ASAP7_75t_R _15637_ (.A1(_08563_),
    .A2(_08565_),
    .B(_08567_),
    .C(_08570_),
    .Y(_08571_));
 NAND2x2_ASAP7_75t_R _15638_ (.A(_08550_),
    .B(_08571_),
    .Y(_08572_));
 BUFx6f_ASAP7_75t_R _15639_ (.A(_08572_),
    .Y(_08573_));
 BUFx4f_ASAP7_75t_R _15640_ (.A(_08550_),
    .Y(_08574_));
 BUFx4f_ASAP7_75t_R _15641_ (.A(_08571_),
    .Y(_08575_));
 INVx1_ASAP7_75t_R _15642_ (.A(_01069_),
    .Y(_08576_));
 AO21x1_ASAP7_75t_R _15643_ (.A1(_08574_),
    .A2(_08575_),
    .B(_08576_),
    .Y(_08577_));
 OA21x2_ASAP7_75t_R _15644_ (.A1(net65),
    .A2(_08573_),
    .B(_08577_),
    .Y(_01220_));
 INVx1_ASAP7_75t_R _15645_ (.A(_01072_),
    .Y(_08578_));
 AO21x1_ASAP7_75t_R _15646_ (.A1(_08574_),
    .A2(_08575_),
    .B(_08578_),
    .Y(_08579_));
 OA21x2_ASAP7_75t_R _15647_ (.A1(net76),
    .A2(_08573_),
    .B(_08579_),
    .Y(_01221_));
 INVx1_ASAP7_75t_R _15648_ (.A(_00732_),
    .Y(_01223_));
 INVx1_ASAP7_75t_R _15649_ (.A(_00699_),
    .Y(_01224_));
 INVx1_ASAP7_75t_R _15650_ (.A(_00666_),
    .Y(_01225_));
 INVx1_ASAP7_75t_R _15651_ (.A(_00633_),
    .Y(_01226_));
 INVx1_ASAP7_75t_R _15652_ (.A(_00600_),
    .Y(_01227_));
 INVx1_ASAP7_75t_R _15653_ (.A(_00566_),
    .Y(_01228_));
 INVx1_ASAP7_75t_R _15654_ (.A(_00500_),
    .Y(_01230_));
 INVx1_ASAP7_75t_R _15655_ (.A(_00467_),
    .Y(_01231_));
 INVx1_ASAP7_75t_R _15656_ (.A(_00434_),
    .Y(_01232_));
 INVx1_ASAP7_75t_R _15657_ (.A(_01031_),
    .Y(_01233_));
 INVx1_ASAP7_75t_R _15658_ (.A(_00401_),
    .Y(_01234_));
 INVx1_ASAP7_75t_R _15659_ (.A(_00368_),
    .Y(_01235_));
 INVx1_ASAP7_75t_R _15660_ (.A(_00335_),
    .Y(_01236_));
 INVx1_ASAP7_75t_R _15661_ (.A(_00301_),
    .Y(_01237_));
 INVx1_ASAP7_75t_R _15662_ (.A(_00268_),
    .Y(_01238_));
 INVx1_ASAP7_75t_R _15663_ (.A(_00235_),
    .Y(_01239_));
 INVx1_ASAP7_75t_R _15664_ (.A(_00202_),
    .Y(_01240_));
 INVx1_ASAP7_75t_R _15665_ (.A(_00168_),
    .Y(_01241_));
 INVx1_ASAP7_75t_R _15666_ (.A(_00135_),
    .Y(_01242_));
 INVx1_ASAP7_75t_R _15667_ (.A(_00101_),
    .Y(_01243_));
 INVx1_ASAP7_75t_R _15668_ (.A(_00998_),
    .Y(_01244_));
 INVx1_ASAP7_75t_R _15669_ (.A(_00067_),
    .Y(_01245_));
 INVx1_ASAP7_75t_R _15670_ (.A(_00035_),
    .Y(_01246_));
 INVx1_ASAP7_75t_R _15671_ (.A(_00965_),
    .Y(_01247_));
 INVx1_ASAP7_75t_R _15672_ (.A(_00932_),
    .Y(_01248_));
 INVx1_ASAP7_75t_R _15673_ (.A(_00898_),
    .Y(_01249_));
 INVx1_ASAP7_75t_R _15674_ (.A(_00865_),
    .Y(_01250_));
 INVx1_ASAP7_75t_R _15675_ (.A(_00831_),
    .Y(_01251_));
 INVx1_ASAP7_75t_R _15676_ (.A(_00798_),
    .Y(_01252_));
 INVx1_ASAP7_75t_R _15677_ (.A(_00764_),
    .Y(_01253_));
 NOR2x2_ASAP7_75t_R _15678_ (.A(_03559_),
    .B(_03560_),
    .Y(_08580_));
 AO21x1_ASAP7_75t_R _15679_ (.A1(_07646_),
    .A2(_07593_),
    .B(_08580_),
    .Y(_08581_));
 OR2x4_ASAP7_75t_R _15680_ (.A(_07589_),
    .B(_08581_),
    .Y(_08582_));
 BUFx6f_ASAP7_75t_R _15681_ (.A(_03574_),
    .Y(_08583_));
 AND2x2_ASAP7_75t_R _15682_ (.A(_08583_),
    .B(_08394_),
    .Y(_08584_));
 BUFx6f_ASAP7_75t_R _15683_ (.A(_07514_),
    .Y(_08585_));
 AND3x1_ASAP7_75t_R _15684_ (.A(\dmem.inter_dmem1[0] ),
    .B(net47),
    .C(_08585_),
    .Y(_08586_));
 BUFx4f_ASAP7_75t_R _15685_ (.A(_03562_),
    .Y(_08587_));
 AO21x1_ASAP7_75t_R _15686_ (.A1(\dmem.inter_dmem0[0] ),
    .A2(\dmem.ce_mem[3] ),
    .B(_08587_),
    .Y(_08588_));
 BUFx4f_ASAP7_75t_R _15687_ (.A(_07514_),
    .Y(_08589_));
 AND4x1_ASAP7_75t_R _15688_ (.A(\dmem.inter_dmem2[0] ),
    .B(_07416_),
    .C(net38),
    .D(_08589_),
    .Y(_08590_));
 BUFx4f_ASAP7_75t_R _15689_ (.A(_07465_),
    .Y(_08591_));
 AND4x1_ASAP7_75t_R _15690_ (.A(\dmem.inter_dmem3[0] ),
    .B(_07416_),
    .C(_08591_),
    .D(_08589_),
    .Y(_08592_));
 OR4x1_ASAP7_75t_R _15691_ (.A(_08586_),
    .B(_08588_),
    .C(_08590_),
    .D(_08592_),
    .Y(_08593_));
 BUFx6f_ASAP7_75t_R _15692_ (.A(_08570_),
    .Y(_08594_));
 AO32x1_ASAP7_75t_R _15693_ (.A1(_08576_),
    .A2(_04849_),
    .A3(_08390_),
    .B1(_08594_),
    .B2(net65),
    .Y(_08595_));
 AO31x2_ASAP7_75t_R _15694_ (.A1(_08582_),
    .A2(_08584_),
    .A3(_08593_),
    .B(_08595_),
    .Y(_08596_));
 BUFx4f_ASAP7_75t_R _15695_ (.A(_08596_),
    .Y(_08597_));
 OA21x2_ASAP7_75t_R _15696_ (.A1(_04072_),
    .A2(_07130_),
    .B(_03566_),
    .Y(_08598_));
 AND2x2_ASAP7_75t_R _15697_ (.A(_03568_),
    .B(_03566_),
    .Y(_08599_));
 AO32x2_ASAP7_75t_R _15698_ (.A1(_03530_),
    .A2(_03557_),
    .A3(_03562_),
    .B1(_08599_),
    .B2(_07372_),
    .Y(_08600_));
 AO21x2_ASAP7_75t_R _15699_ (.A1(_03574_),
    .A2(_08600_),
    .B(_06140_),
    .Y(_08601_));
 NOR2x2_ASAP7_75t_R _15700_ (.A(_08598_),
    .B(_08601_),
    .Y(_08602_));
 NAND2x2_ASAP7_75t_R _15701_ (.A(_03566_),
    .B(_07020_),
    .Y(_08603_));
 INVx1_ASAP7_75t_R _15702_ (.A(net2),
    .Y(_08604_));
 OR3x2_ASAP7_75t_R _15703_ (.A(_04072_),
    .B(net3),
    .C(_08604_),
    .Y(_08605_));
 NOR2x2_ASAP7_75t_R _15704_ (.A(_08603_),
    .B(_08605_),
    .Y(_08606_));
 BUFx12_ASAP7_75t_R _15705_ (.A(_08606_),
    .Y(_08607_));
 NAND2x2_ASAP7_75t_R _15706_ (.A(_08602_),
    .B(_08607_),
    .Y(_08608_));
 BUFx6f_ASAP7_75t_R _15707_ (.A(_08608_),
    .Y(_08609_));
 BUFx12_ASAP7_75t_R _15708_ (.A(_08608_),
    .Y(_08610_));
 NAND2x1_ASAP7_75t_R _15709_ (.A(_00010_),
    .B(_08610_),
    .Y(_08611_));
 OA21x2_ASAP7_75t_R _15710_ (.A1(_08597_),
    .A2(_08609_),
    .B(_08611_),
    .Y(_01254_));
 OR3x1_ASAP7_75t_R _15711_ (.A(_03562_),
    .B(_05853_),
    .C(_05946_),
    .Y(_08612_));
 AND2x2_ASAP7_75t_R _15712_ (.A(_08580_),
    .B(_08612_),
    .Y(_08613_));
 AND3x4_ASAP7_75t_R _15713_ (.A(_07416_),
    .B(net38),
    .C(_07514_),
    .Y(_08614_));
 BUFx6f_ASAP7_75t_R _15714_ (.A(_08614_),
    .Y(\dmem.ce_mem[1] ));
 AND3x1_ASAP7_75t_R _15715_ (.A(\dmem.inter_dmem1[10] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_08615_));
 AOI21x1_ASAP7_75t_R _15716_ (.A1(_07280_),
    .A2(_07327_),
    .B(_07337_),
    .Y(_08616_));
 BUFx3_ASAP7_75t_R _15717_ (.A(_08616_),
    .Y(_08617_));
 BUFx3_ASAP7_75t_R _15718_ (.A(_08617_),
    .Y(_08618_));
 NOR2x2_ASAP7_75t_R _15719_ (.A(_07407_),
    .B(_07413_),
    .Y(_08619_));
 BUFx3_ASAP7_75t_R _15720_ (.A(_08619_),
    .Y(_08620_));
 BUFx6f_ASAP7_75t_R _15721_ (.A(_08620_),
    .Y(_08621_));
 OA211x2_ASAP7_75t_R _15722_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08591_),
    .C(\dmem.inter_dmem3[10] ),
    .Y(_08622_));
 OA21x2_ASAP7_75t_R _15723_ (.A1(_08615_),
    .A2(_08622_),
    .B(_08585_),
    .Y(_08623_));
 AO221x1_ASAP7_75t_R _15724_ (.A1(\dmem.inter_dmem0[10] ),
    .A2(\dmem.ce_mem[3] ),
    .B1(\dmem.ce_mem[1] ),
    .B2(\dmem.inter_dmem2[10] ),
    .C(_08623_),
    .Y(_08624_));
 OA211x2_ASAP7_75t_R _15725_ (.A1(_07420_),
    .A2(_07433_),
    .B(\dmem.inter_dmem2[7] ),
    .C(_07464_),
    .Y(_08625_));
 AO221x1_ASAP7_75t_R _15726_ (.A1(_07339_),
    .A2(_07415_),
    .B1(_07465_),
    .B2(\dmem.inter_dmem3[7] ),
    .C(_08625_),
    .Y(_08626_));
 OA211x2_ASAP7_75t_R _15727_ (.A1(\dmem.inter_dmem1[7] ),
    .A2(_07416_),
    .B(_07514_),
    .C(_08626_),
    .Y(_08627_));
 BUFx4f_ASAP7_75t_R _15728_ (.A(_07515_),
    .Y(_08628_));
 AND2x2_ASAP7_75t_R _15729_ (.A(\dmem.inter_dmem0[7] ),
    .B(_08628_),
    .Y(_08629_));
 OR4x1_ASAP7_75t_R _15730_ (.A(_03528_),
    .B(_03534_),
    .C(_03559_),
    .D(_07239_),
    .Y(_08630_));
 AND3x2_ASAP7_75t_R _15731_ (.A(_08580_),
    .B(_05852_),
    .C(_05945_),
    .Y(_08631_));
 OA211x2_ASAP7_75t_R _15732_ (.A1(_08627_),
    .A2(_08629_),
    .B(_08630_),
    .C(_08631_),
    .Y(_08632_));
 AND3x4_ASAP7_75t_R _15733_ (.A(_03562_),
    .B(_03574_),
    .C(_08394_),
    .Y(_08633_));
 BUFx10_ASAP7_75t_R _15734_ (.A(_08633_),
    .Y(_08634_));
 OA21x2_ASAP7_75t_R _15735_ (.A1(_01073_),
    .A2(_01160_),
    .B(_01076_),
    .Y(_08635_));
 OA21x2_ASAP7_75t_R _15736_ (.A1(_01075_),
    .A2(_08635_),
    .B(_01079_),
    .Y(_08636_));
 OA21x2_ASAP7_75t_R _15737_ (.A1(_01078_),
    .A2(_08636_),
    .B(_01082_),
    .Y(_08637_));
 OA21x2_ASAP7_75t_R _15738_ (.A1(_01088_),
    .A2(_01087_),
    .B(_01091_),
    .Y(_08638_));
 OA21x2_ASAP7_75t_R _15739_ (.A1(_01090_),
    .A2(_08638_),
    .B(_01094_),
    .Y(_08639_));
 AND3x1_ASAP7_75t_R _15740_ (.A(_01085_),
    .B(_01097_),
    .C(_08639_),
    .Y(_08640_));
 OA21x2_ASAP7_75t_R _15741_ (.A1(_01081_),
    .A2(_08637_),
    .B(_08640_),
    .Y(_08641_));
 OR3x1_ASAP7_75t_R _15742_ (.A(_01084_),
    .B(_01087_),
    .C(_01090_),
    .Y(_08642_));
 AND3x1_ASAP7_75t_R _15743_ (.A(_01097_),
    .B(_08639_),
    .C(_08642_),
    .Y(_08643_));
 AO21x1_ASAP7_75t_R _15744_ (.A1(_01093_),
    .A2(_01097_),
    .B(_08643_),
    .Y(_08644_));
 OR2x2_ASAP7_75t_R _15745_ (.A(_08641_),
    .B(_08644_),
    .Y(_08645_));
 XOR2x1_ASAP7_75t_R _15746_ (.A(_01096_),
    .Y(_08646_),
    .B(_08645_));
 AND2x4_ASAP7_75t_R _15747_ (.A(_04165_),
    .B(_08390_),
    .Y(_08647_));
 BUFx6f_ASAP7_75t_R _15748_ (.A(_08647_),
    .Y(_08648_));
 OR3x2_ASAP7_75t_R _15749_ (.A(_01077_),
    .B(_01080_),
    .C(_01218_),
    .Y(_08649_));
 OR5x2_ASAP7_75t_R _15750_ (.A(_03479_),
    .B(_01086_),
    .C(_01089_),
    .D(_01092_),
    .E(_08649_),
    .Y(_08650_));
 BUFx4f_ASAP7_75t_R _15751_ (.A(_08650_),
    .Y(_08651_));
 XNOR2x1_ASAP7_75t_R _15752_ (.B(_08651_),
    .Y(_08652_),
    .A(net66));
 AO222x2_ASAP7_75t_R _15753_ (.A1(net33),
    .A2(_08634_),
    .B1(_08646_),
    .B2(_08648_),
    .C1(_08652_),
    .C2(_08570_),
    .Y(_08653_));
 AO211x2_ASAP7_75t_R _15754_ (.A1(_08613_),
    .A2(_08624_),
    .B(_08632_),
    .C(_08653_),
    .Y(_08654_));
 NAND2x1_ASAP7_75t_R _15755_ (.A(_00742_),
    .B(_08610_),
    .Y(_08655_));
 OA21x2_ASAP7_75t_R _15756_ (.A1(_08609_),
    .A2(_08654_),
    .B(_08655_),
    .Y(_01255_));
 OA211x2_ASAP7_75t_R _15757_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08591_),
    .C(\dmem.inter_dmem3[11] ),
    .Y(_08656_));
 AO21x1_ASAP7_75t_R _15758_ (.A1(\dmem.inter_dmem1[11] ),
    .A2(net47),
    .B(_08656_),
    .Y(_08657_));
 BUFx6f_ASAP7_75t_R _15759_ (.A(_08589_),
    .Y(_08658_));
 AND2x2_ASAP7_75t_R _15760_ (.A(\dmem.inter_dmem0[11] ),
    .B(\dmem.ce_mem[3] ),
    .Y(_08659_));
 AO221x1_ASAP7_75t_R _15761_ (.A1(\dmem.inter_dmem2[11] ),
    .A2(\dmem.ce_mem[1] ),
    .B1(_08657_),
    .B2(_08658_),
    .C(_08659_),
    .Y(_08660_));
 OR3x4_ASAP7_75t_R _15762_ (.A(_08580_),
    .B(_08569_),
    .C(_08647_),
    .Y(_08661_));
 BUFx6f_ASAP7_75t_R _15763_ (.A(_08661_),
    .Y(_08662_));
 OA21x2_ASAP7_75t_R _15764_ (.A1(_01071_),
    .A2(_09946_),
    .B(_01074_),
    .Y(_08663_));
 OA21x2_ASAP7_75t_R _15765_ (.A1(_01073_),
    .A2(_08663_),
    .B(_01076_),
    .Y(_08664_));
 AND3x1_ASAP7_75t_R _15766_ (.A(_01079_),
    .B(_01082_),
    .C(_01085_),
    .Y(_08665_));
 OA21x2_ASAP7_75t_R _15767_ (.A1(_01075_),
    .A2(_08664_),
    .B(_08665_),
    .Y(_08666_));
 AO21x1_ASAP7_75t_R _15768_ (.A1(_01078_),
    .A2(_01082_),
    .B(_01081_),
    .Y(_08667_));
 AND2x2_ASAP7_75t_R _15769_ (.A(_01085_),
    .B(_08667_),
    .Y(_08668_));
 OR5x2_ASAP7_75t_R _15770_ (.A(_01093_),
    .B(_01096_),
    .C(_08642_),
    .D(_08666_),
    .E(_08668_),
    .Y(_08669_));
 OA21x2_ASAP7_75t_R _15771_ (.A1(_01093_),
    .A2(_08639_),
    .B(_01097_),
    .Y(_08670_));
 OA21x2_ASAP7_75t_R _15772_ (.A1(_01096_),
    .A2(_08670_),
    .B(_01100_),
    .Y(_08671_));
 AND2x2_ASAP7_75t_R _15773_ (.A(_08669_),
    .B(_08671_),
    .Y(_08672_));
 XOR2x2_ASAP7_75t_R _15774_ (.A(_01099_),
    .B(_08672_),
    .Y(_08673_));
 OR3x2_ASAP7_75t_R _15775_ (.A(_10109_),
    .B(_10110_),
    .C(_01077_),
    .Y(_08674_));
 OR2x2_ASAP7_75t_R _15776_ (.A(_01080_),
    .B(_08674_),
    .Y(_08675_));
 OR4x2_ASAP7_75t_R _15777_ (.A(_03479_),
    .B(_01086_),
    .C(_01089_),
    .D(_08675_),
    .Y(_08676_));
 OR3x1_ASAP7_75t_R _15778_ (.A(_01092_),
    .B(_01095_),
    .C(_08676_),
    .Y(_08677_));
 XNOR2x1_ASAP7_75t_R _15779_ (.B(_08677_),
    .Y(_08678_),
    .A(net67));
 AOI22x1_ASAP7_75t_R _15780_ (.A1(_08648_),
    .A2(_08673_),
    .B1(_08678_),
    .B2(_08594_),
    .Y(_08679_));
 OAI21x1_ASAP7_75t_R _15781_ (.A1(_08037_),
    .A2(_08662_),
    .B(_08679_),
    .Y(_08680_));
 AO211x2_ASAP7_75t_R _15782_ (.A1(_08613_),
    .A2(_08660_),
    .B(_08680_),
    .C(_08632_),
    .Y(_08681_));
 NAND2x1_ASAP7_75t_R _15783_ (.A(_00709_),
    .B(_08610_),
    .Y(_08682_));
 OA21x2_ASAP7_75t_R _15784_ (.A1(_08609_),
    .A2(_08681_),
    .B(_08682_),
    .Y(_01256_));
 AND3x1_ASAP7_75t_R _15785_ (.A(\dmem.inter_dmem1[12] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_08683_));
 OA211x2_ASAP7_75t_R _15786_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08591_),
    .C(\dmem.inter_dmem3[12] ),
    .Y(_08684_));
 OA21x2_ASAP7_75t_R _15787_ (.A1(_08683_),
    .A2(_08684_),
    .B(_08585_),
    .Y(_08685_));
 AO221x1_ASAP7_75t_R _15788_ (.A1(\dmem.inter_dmem0[12] ),
    .A2(\dmem.ce_mem[3] ),
    .B1(\dmem.ce_mem[1] ),
    .B2(\dmem.inter_dmem2[12] ),
    .C(_08685_),
    .Y(_08686_));
 BUFx10_ASAP7_75t_R _15789_ (.A(_08647_),
    .Y(_08687_));
 OR3x1_ASAP7_75t_R _15790_ (.A(_01096_),
    .B(_08641_),
    .C(_08644_),
    .Y(_08688_));
 AO21x1_ASAP7_75t_R _15791_ (.A1(_01100_),
    .A2(_08688_),
    .B(_01099_),
    .Y(_08689_));
 AND2x2_ASAP7_75t_R _15792_ (.A(_01103_),
    .B(_08689_),
    .Y(_08690_));
 XNOR2x1_ASAP7_75t_R _15793_ (.B(_08690_),
    .Y(_08691_),
    .A(_01102_));
 OR3x1_ASAP7_75t_R _15794_ (.A(_01095_),
    .B(_01098_),
    .C(_08651_),
    .Y(_08692_));
 XNOR2x1_ASAP7_75t_R _15795_ (.B(_08692_),
    .Y(_08693_),
    .A(net68));
 INVx1_ASAP7_75t_R _15796_ (.A(_08693_),
    .Y(_08694_));
 AO221x1_ASAP7_75t_R _15797_ (.A1(_08687_),
    .A2(_08691_),
    .B1(_08694_),
    .B2(_08570_),
    .C(_08580_),
    .Y(_08695_));
 AOI21x1_ASAP7_75t_R _15798_ (.A1(_08057_),
    .A2(_08584_),
    .B(_08695_),
    .Y(_08696_));
 AO211x2_ASAP7_75t_R _15799_ (.A1(_08613_),
    .A2(_08686_),
    .B(_08696_),
    .C(_08632_),
    .Y(_08697_));
 NAND2x1_ASAP7_75t_R _15800_ (.A(_00676_),
    .B(_08610_),
    .Y(_08698_));
 OA21x2_ASAP7_75t_R _15801_ (.A1(_08609_),
    .A2(_08697_),
    .B(_08698_),
    .Y(_01257_));
 AND2x6_ASAP7_75t_R _15802_ (.A(_08602_),
    .B(_08607_),
    .Y(_08699_));
 BUFx10_ASAP7_75t_R _15803_ (.A(_08699_),
    .Y(_08700_));
 AND2x2_ASAP7_75t_R _15804_ (.A(_07643_),
    .B(_08633_),
    .Y(_08701_));
 INVx2_ASAP7_75t_R _15805_ (.A(\dmem.inter_dmem2[13] ),
    .Y(_08702_));
 BUFx3_ASAP7_75t_R _15806_ (.A(_07465_),
    .Y(_08703_));
 OR4x1_ASAP7_75t_R _15807_ (.A(_08702_),
    .B(_07417_),
    .C(_08703_),
    .D(_07515_),
    .Y(_08704_));
 NAND2x1_ASAP7_75t_R _15808_ (.A(\dmem.inter_dmem0[13] ),
    .B(_07515_),
    .Y(_08705_));
 AND3x1_ASAP7_75t_R _15809_ (.A(\dmem.inter_dmem1[13] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_08706_));
 OA211x2_ASAP7_75t_R _15810_ (.A1(_08617_),
    .A2(_08620_),
    .B(_07465_),
    .C(\dmem.inter_dmem3[13] ),
    .Y(_08707_));
 OAI21x1_ASAP7_75t_R _15811_ (.A1(_08706_),
    .A2(_08707_),
    .B(_08589_),
    .Y(_08708_));
 AO33x2_ASAP7_75t_R _15812_ (.A1(_08580_),
    .A2(_05852_),
    .A3(_05945_),
    .B1(_08704_),
    .B2(_08705_),
    .B3(_08708_),
    .Y(_08709_));
 OR4x1_ASAP7_75t_R _15813_ (.A(_03528_),
    .B(_03534_),
    .C(_03559_),
    .D(_07239_),
    .Y(_08710_));
 AND2x2_ASAP7_75t_R _15814_ (.A(_08631_),
    .B(_08710_),
    .Y(_08711_));
 AO21x1_ASAP7_75t_R _15815_ (.A1(\dmem.inter_dmem0[7] ),
    .A2(_07515_),
    .B(_03562_),
    .Y(_08712_));
 OAI22x1_ASAP7_75t_R _15816_ (.A1(_03562_),
    .A2(_08711_),
    .B1(_08712_),
    .B2(_08627_),
    .Y(_08713_));
 OR2x2_ASAP7_75t_R _15817_ (.A(_01092_),
    .B(_08676_),
    .Y(_08714_));
 BUFx4f_ASAP7_75t_R _15818_ (.A(_08714_),
    .Y(_08715_));
 OR4x1_ASAP7_75t_R _15819_ (.A(_01095_),
    .B(_01098_),
    .C(_01101_),
    .D(_08715_),
    .Y(_08716_));
 XNOR2x1_ASAP7_75t_R _15820_ (.B(_08716_),
    .Y(_08717_),
    .A(_01104_));
 AND3x1_ASAP7_75t_R _15821_ (.A(_07591_),
    .B(_08079_),
    .C(_08633_),
    .Y(_08718_));
 OA21x2_ASAP7_75t_R _15822_ (.A1(_01099_),
    .A2(_08672_),
    .B(_01103_),
    .Y(_08719_));
 OA21x2_ASAP7_75t_R _15823_ (.A1(_01102_),
    .A2(_08719_),
    .B(_01106_),
    .Y(_08720_));
 XNOR2x2_ASAP7_75t_R _15824_ (.A(_01105_),
    .B(_08720_),
    .Y(_08721_));
 AO222x2_ASAP7_75t_R _15825_ (.A1(_08570_),
    .A2(_08717_),
    .B1(_08718_),
    .B2(_08076_),
    .C1(_08687_),
    .C2(_08721_),
    .Y(_08722_));
 AO221x1_ASAP7_75t_R _15826_ (.A1(_08071_),
    .A2(_08701_),
    .B1(_08709_),
    .B2(_08713_),
    .C(_08722_),
    .Y(_08723_));
 BUFx6f_ASAP7_75t_R _15827_ (.A(_08723_),
    .Y(_08724_));
 BUFx6f_ASAP7_75t_R _15828_ (.A(_08724_),
    .Y(_08725_));
 BUFx12_ASAP7_75t_R _15829_ (.A(_08608_),
    .Y(_08726_));
 AND2x2_ASAP7_75t_R _15830_ (.A(_00643_),
    .B(_08726_),
    .Y(_08727_));
 AOI21x1_ASAP7_75t_R _15831_ (.A1(_08700_),
    .A2(_08725_),
    .B(_08727_),
    .Y(_01258_));
 AND3x1_ASAP7_75t_R _15832_ (.A(\dmem.inter_dmem1[14] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_08728_));
 OA211x2_ASAP7_75t_R _15833_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08591_),
    .C(\dmem.inter_dmem3[14] ),
    .Y(_08729_));
 OA21x2_ASAP7_75t_R _15834_ (.A1(_08728_),
    .A2(_08729_),
    .B(_08585_),
    .Y(_08730_));
 AO221x1_ASAP7_75t_R _15835_ (.A1(\dmem.inter_dmem0[14] ),
    .A2(\dmem.ce_mem[3] ),
    .B1(\dmem.ce_mem[1] ),
    .B2(\dmem.inter_dmem2[14] ),
    .C(_08730_),
    .Y(_08731_));
 NAND2x1_ASAP7_75t_R _15836_ (.A(_08583_),
    .B(_08394_),
    .Y(_08732_));
 OR5x2_ASAP7_75t_R _15837_ (.A(_01095_),
    .B(_01098_),
    .C(_01101_),
    .D(_01104_),
    .E(_08651_),
    .Y(_08733_));
 XNOR2x1_ASAP7_75t_R _15838_ (.B(_08733_),
    .Y(_08734_),
    .A(net70));
 OR3x2_ASAP7_75t_R _15839_ (.A(_01099_),
    .B(_01102_),
    .C(_01105_),
    .Y(_08735_));
 OA21x2_ASAP7_75t_R _15840_ (.A1(_01100_),
    .A2(_01099_),
    .B(_01103_),
    .Y(_08736_));
 OA21x2_ASAP7_75t_R _15841_ (.A1(_01102_),
    .A2(_08736_),
    .B(_01106_),
    .Y(_08737_));
 OA21x2_ASAP7_75t_R _15842_ (.A1(_01105_),
    .A2(_08737_),
    .B(_01109_),
    .Y(_08738_));
 OA21x2_ASAP7_75t_R _15843_ (.A1(_08688_),
    .A2(_08735_),
    .B(_08738_),
    .Y(_08739_));
 XNOR2x2_ASAP7_75t_R _15844_ (.A(_01108_),
    .B(_08739_),
    .Y(_08740_));
 NAND2x1_ASAP7_75t_R _15845_ (.A(_08647_),
    .B(_08740_),
    .Y(_08741_));
 OA211x2_ASAP7_75t_R _15846_ (.A1(_08583_),
    .A2(_08734_),
    .B(_08741_),
    .C(_08587_),
    .Y(_08742_));
 OA21x2_ASAP7_75t_R _15847_ (.A1(net37),
    .A2(_08732_),
    .B(_08742_),
    .Y(_08743_));
 AO211x2_ASAP7_75t_R _15848_ (.A1(_08613_),
    .A2(_08731_),
    .B(_08743_),
    .C(_08632_),
    .Y(_08744_));
 NAND2x1_ASAP7_75t_R _15849_ (.A(_00610_),
    .B(_08610_),
    .Y(_08745_));
 OA21x2_ASAP7_75t_R _15850_ (.A1(_08609_),
    .A2(_08744_),
    .B(_08745_),
    .Y(_01259_));
 OA22x2_ASAP7_75t_R _15851_ (.A1(_03562_),
    .A2(_08711_),
    .B1(_08712_),
    .B2(_08627_),
    .Y(_08746_));
 BUFx6f_ASAP7_75t_R _15852_ (.A(_08746_),
    .Y(_08747_));
 BUFx12f_ASAP7_75t_R _15853_ (.A(_08747_),
    .Y(_08748_));
 AND2x2_ASAP7_75t_R _15854_ (.A(\dmem.inter_dmem0[15] ),
    .B(_07515_),
    .Y(_08749_));
 OA211x2_ASAP7_75t_R _15855_ (.A1(_08616_),
    .A2(_08619_),
    .B(net38),
    .C(\dmem.inter_dmem2[15] ),
    .Y(_08750_));
 AND3x1_ASAP7_75t_R _15856_ (.A(\dmem.inter_dmem1[15] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_08751_));
 OA21x2_ASAP7_75t_R _15857_ (.A1(_08750_),
    .A2(_08751_),
    .B(_07514_),
    .Y(_08752_));
 AND4x2_ASAP7_75t_R _15858_ (.A(\dmem.inter_dmem3[15] ),
    .B(_07416_),
    .C(_07465_),
    .D(_07514_),
    .Y(_08753_));
 OA33x2_ASAP7_75t_R _15859_ (.A1(_08587_),
    .A2(_05853_),
    .A3(_05946_),
    .B1(_08749_),
    .B2(_08752_),
    .B3(_08753_),
    .Y(_08754_));
 OR5x2_ASAP7_75t_R _15860_ (.A(_01095_),
    .B(_01098_),
    .C(_01101_),
    .D(_01104_),
    .E(_01107_),
    .Y(_08755_));
 NOR2x1_ASAP7_75t_R _15861_ (.A(_08715_),
    .B(_08755_),
    .Y(_08756_));
 XNOR2x1_ASAP7_75t_R _15862_ (.B(_08756_),
    .Y(_08757_),
    .A(net71));
 OA21x2_ASAP7_75t_R _15863_ (.A1(_01103_),
    .A2(_01102_),
    .B(_01106_),
    .Y(_08758_));
 OA21x2_ASAP7_75t_R _15864_ (.A1(_01105_),
    .A2(_08758_),
    .B(_01109_),
    .Y(_08759_));
 OA21x2_ASAP7_75t_R _15865_ (.A1(_08672_),
    .A2(_08735_),
    .B(_08759_),
    .Y(_08760_));
 OA21x2_ASAP7_75t_R _15866_ (.A1(_01108_),
    .A2(_08760_),
    .B(_01112_),
    .Y(_08761_));
 XOR2x1_ASAP7_75t_R _15867_ (.A(_01111_),
    .Y(_08762_),
    .B(_08761_));
 NOR2x1_ASAP7_75t_R _15868_ (.A(_08394_),
    .B(_08762_),
    .Y(_08763_));
 AOI221x1_ASAP7_75t_R _15869_ (.A1(_08591_),
    .A2(_08634_),
    .B1(_08757_),
    .B2(_08594_),
    .C(_08763_),
    .Y(_08764_));
 OAI21x1_ASAP7_75t_R _15870_ (.A1(_08748_),
    .A2(_08754_),
    .B(_08764_),
    .Y(_08765_));
 BUFx10_ASAP7_75t_R _15871_ (.A(_08765_),
    .Y(_08766_));
 AND2x2_ASAP7_75t_R _15872_ (.A(_00576_),
    .B(_08726_),
    .Y(_08767_));
 AOI21x1_ASAP7_75t_R _15873_ (.A1(_08700_),
    .A2(_08766_),
    .B(_08767_),
    .Y(_01260_));
 OR3x1_ASAP7_75t_R _15874_ (.A(_04072_),
    .B(_03562_),
    .C(_07241_),
    .Y(_08768_));
 BUFx4f_ASAP7_75t_R _15875_ (.A(_08768_),
    .Y(_08769_));
 BUFx6f_ASAP7_75t_R _15876_ (.A(_08769_),
    .Y(_08770_));
 BUFx3_ASAP7_75t_R _15877_ (.A(_08614_),
    .Y(_08771_));
 BUFx6f_ASAP7_75t_R _15878_ (.A(_07417_),
    .Y(_08772_));
 BUFx3_ASAP7_75t_R _15879_ (.A(_08616_),
    .Y(_08773_));
 BUFx3_ASAP7_75t_R _15880_ (.A(_08619_),
    .Y(_08774_));
 OA211x2_ASAP7_75t_R _15881_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[16] ),
    .Y(_08775_));
 AO21x1_ASAP7_75t_R _15882_ (.A1(\dmem.inter_dmem1[16] ),
    .A2(_08772_),
    .B(_08775_),
    .Y(_08776_));
 AND2x2_ASAP7_75t_R _15883_ (.A(\dmem.inter_dmem0[16] ),
    .B(_08628_),
    .Y(_08777_));
 AO221x1_ASAP7_75t_R _15884_ (.A1(\dmem.inter_dmem2[16] ),
    .A2(_08771_),
    .B1(_08776_),
    .B2(_08658_),
    .C(_08777_),
    .Y(_08778_));
 AND5x1_ASAP7_75t_R _15885_ (.A(_03382_),
    .B(_08389_),
    .C(_07332_),
    .D(_03526_),
    .E(_07274_),
    .Y(_08779_));
 OA31x2_ASAP7_75t_R _15886_ (.A1(_08749_),
    .A2(_08752_),
    .A3(_08753_),
    .B1(_08779_),
    .Y(_08780_));
 BUFx4f_ASAP7_75t_R _15887_ (.A(_08780_),
    .Y(_08781_));
 AO211x2_ASAP7_75t_R _15888_ (.A1(_08770_),
    .A2(_08778_),
    .B(_08781_),
    .C(_08748_),
    .Y(_08782_));
 BUFx10_ASAP7_75t_R _15889_ (.A(_08782_),
    .Y(_08783_));
 NAND2x2_ASAP7_75t_R _15890_ (.A(_08631_),
    .B(_08713_),
    .Y(_08784_));
 BUFx12f_ASAP7_75t_R _15891_ (.A(_08784_),
    .Y(_08785_));
 OR2x6_ASAP7_75t_R _15892_ (.A(net39),
    .B(_08661_),
    .Y(_08786_));
 OR3x1_ASAP7_75t_R _15893_ (.A(_01110_),
    .B(_08651_),
    .C(_08755_),
    .Y(_08787_));
 XNOR2x1_ASAP7_75t_R _15894_ (.B(_08787_),
    .Y(_08788_),
    .A(_01113_));
 OR5x1_ASAP7_75t_R _15895_ (.A(_01096_),
    .B(_01108_),
    .C(_08641_),
    .D(_08644_),
    .E(_08735_),
    .Y(_08789_));
 OA21x2_ASAP7_75t_R _15896_ (.A1(_01108_),
    .A2(_08738_),
    .B(_01112_),
    .Y(_08790_));
 AO21x1_ASAP7_75t_R _15897_ (.A1(_08789_),
    .A2(_08790_),
    .B(_01111_),
    .Y(_08791_));
 AND2x2_ASAP7_75t_R _15898_ (.A(_01115_),
    .B(_08791_),
    .Y(_08792_));
 XNOR2x1_ASAP7_75t_R _15899_ (.B(_08792_),
    .Y(_08793_),
    .A(_01114_));
 AOI22x1_ASAP7_75t_R _15900_ (.A1(_08594_),
    .A2(_08788_),
    .B1(_08793_),
    .B2(_08648_),
    .Y(_08794_));
 AND3x1_ASAP7_75t_R _15901_ (.A(_08700_),
    .B(_08786_),
    .C(_08794_),
    .Y(_08795_));
 BUFx6f_ASAP7_75t_R _15902_ (.A(_08608_),
    .Y(_08796_));
 INVx1_ASAP7_75t_R _15903_ (.A(_00543_),
    .Y(_08797_));
 AO32x1_ASAP7_75t_R _15904_ (.A1(_08783_),
    .A2(_08785_),
    .A3(_08795_),
    .B1(_08796_),
    .B2(_08797_),
    .Y(_01261_));
 BUFx6f_ASAP7_75t_R _15905_ (.A(_08784_),
    .Y(_08798_));
 BUFx4f_ASAP7_75t_R _15906_ (.A(_08798_),
    .Y(_08799_));
 OA211x2_ASAP7_75t_R _15907_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[17] ),
    .Y(_08800_));
 AO21x1_ASAP7_75t_R _15908_ (.A1(\dmem.inter_dmem1[17] ),
    .A2(_08772_),
    .B(_08800_),
    .Y(_08801_));
 AND2x2_ASAP7_75t_R _15909_ (.A(\dmem.inter_dmem0[17] ),
    .B(_08628_),
    .Y(_08802_));
 AO221x1_ASAP7_75t_R _15910_ (.A1(\dmem.inter_dmem2[17] ),
    .A2(_08771_),
    .B1(_08801_),
    .B2(_08658_),
    .C(_08802_),
    .Y(_08803_));
 AO211x2_ASAP7_75t_R _15911_ (.A1(_08770_),
    .A2(_08803_),
    .B(_08781_),
    .C(_08748_),
    .Y(_08804_));
 BUFx4f_ASAP7_75t_R _15912_ (.A(_08804_),
    .Y(_08805_));
 BUFx4f_ASAP7_75t_R _15913_ (.A(_08699_),
    .Y(_08806_));
 AND3x2_ASAP7_75t_R _15914_ (.A(_07592_),
    .B(_08128_),
    .C(_08634_),
    .Y(_08807_));
 AND3x2_ASAP7_75t_R _15915_ (.A(_08136_),
    .B(_08138_),
    .C(_08701_),
    .Y(_08808_));
 OR3x2_ASAP7_75t_R _15916_ (.A(_01110_),
    .B(_01113_),
    .C(_08755_),
    .Y(_08809_));
 NOR2x1_ASAP7_75t_R _15917_ (.A(_08715_),
    .B(_08809_),
    .Y(_08810_));
 XNOR2x2_ASAP7_75t_R _15918_ (.A(net73),
    .B(_08810_),
    .Y(_08811_));
 OR3x1_ASAP7_75t_R _15919_ (.A(_01108_),
    .B(_01111_),
    .C(_08735_),
    .Y(_08812_));
 AO21x1_ASAP7_75t_R _15920_ (.A1(_08669_),
    .A2(_08671_),
    .B(_08812_),
    .Y(_08813_));
 OR3x1_ASAP7_75t_R _15921_ (.A(_01108_),
    .B(_01111_),
    .C(_08759_),
    .Y(_08814_));
 OA21x2_ASAP7_75t_R _15922_ (.A1(_01112_),
    .A2(_01111_),
    .B(_08814_),
    .Y(_08815_));
 AND3x1_ASAP7_75t_R _15923_ (.A(_01115_),
    .B(_08813_),
    .C(_08815_),
    .Y(_08816_));
 OA21x2_ASAP7_75t_R _15924_ (.A1(_01114_),
    .A2(_08816_),
    .B(_01118_),
    .Y(_08817_));
 XNOR2x1_ASAP7_75t_R _15925_ (.B(_08817_),
    .Y(_08818_),
    .A(_01117_));
 AOI22x1_ASAP7_75t_R _15926_ (.A1(_08569_),
    .A2(_08811_),
    .B1(_08818_),
    .B2(_08647_),
    .Y(_08819_));
 INVx2_ASAP7_75t_R _15927_ (.A(_08819_),
    .Y(_08820_));
 NOR3x2_ASAP7_75t_R _15928_ (.B(_08808_),
    .C(_08820_),
    .Y(_08821_),
    .A(_08807_));
 AND2x2_ASAP7_75t_R _15929_ (.A(_08806_),
    .B(_08821_),
    .Y(_08822_));
 INVx1_ASAP7_75t_R _15930_ (.A(_00510_),
    .Y(_08823_));
 AO32x1_ASAP7_75t_R _15931_ (.A1(_08799_),
    .A2(_08805_),
    .A3(_08822_),
    .B1(_08796_),
    .B2(_08823_),
    .Y(_01262_));
 OA211x2_ASAP7_75t_R _15932_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[18] ),
    .Y(_08824_));
 AO21x1_ASAP7_75t_R _15933_ (.A1(\dmem.inter_dmem1[18] ),
    .A2(_08772_),
    .B(_08824_),
    .Y(_08825_));
 BUFx3_ASAP7_75t_R _15934_ (.A(_08589_),
    .Y(_08826_));
 AND2x2_ASAP7_75t_R _15935_ (.A(\dmem.inter_dmem0[18] ),
    .B(_08628_),
    .Y(_08827_));
 AO221x1_ASAP7_75t_R _15936_ (.A1(\dmem.inter_dmem2[18] ),
    .A2(_08771_),
    .B1(_08825_),
    .B2(_08826_),
    .C(_08827_),
    .Y(_08828_));
 AO211x2_ASAP7_75t_R _15937_ (.A1(_08770_),
    .A2(_08828_),
    .B(_08781_),
    .C(_08748_),
    .Y(_08829_));
 BUFx4f_ASAP7_75t_R _15938_ (.A(_08829_),
    .Y(_08830_));
 INVx1_ASAP7_75t_R _15939_ (.A(_08163_),
    .Y(_08831_));
 AND3x1_ASAP7_75t_R _15940_ (.A(_08145_),
    .B(_08831_),
    .C(_08152_),
    .Y(_08832_));
 NAND2x1_ASAP7_75t_R _15941_ (.A(_08143_),
    .B(_08634_),
    .Y(_08833_));
 OR2x6_ASAP7_75t_R _15942_ (.A(_08832_),
    .B(_08833_),
    .Y(_08834_));
 OR3x1_ASAP7_75t_R _15943_ (.A(_01116_),
    .B(_08651_),
    .C(_08809_),
    .Y(_08835_));
 XNOR2x1_ASAP7_75t_R _15944_ (.B(_08835_),
    .Y(_08836_),
    .A(_01119_));
 OA21x2_ASAP7_75t_R _15945_ (.A1(_01118_),
    .A2(_01117_),
    .B(_01121_),
    .Y(_08837_));
 OR3x1_ASAP7_75t_R _15946_ (.A(_01114_),
    .B(_01117_),
    .C(_08792_),
    .Y(_08838_));
 AND2x2_ASAP7_75t_R _15947_ (.A(_08837_),
    .B(_08838_),
    .Y(_08839_));
 XNOR2x1_ASAP7_75t_R _15948_ (.B(_08839_),
    .Y(_08840_),
    .A(_01120_));
 AOI22x1_ASAP7_75t_R _15949_ (.A1(_08594_),
    .A2(_08836_),
    .B1(_08840_),
    .B2(_08648_),
    .Y(_08841_));
 AND3x1_ASAP7_75t_R _15950_ (.A(_08806_),
    .B(_08834_),
    .C(_08841_),
    .Y(_08842_));
 INVx1_ASAP7_75t_R _15951_ (.A(_00477_),
    .Y(_08843_));
 AO32x1_ASAP7_75t_R _15952_ (.A1(_08799_),
    .A2(_08830_),
    .A3(_08842_),
    .B1(_08796_),
    .B2(_08843_),
    .Y(_01263_));
 OA211x2_ASAP7_75t_R _15953_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[19] ),
    .Y(_08844_));
 AO21x1_ASAP7_75t_R _15954_ (.A1(\dmem.inter_dmem1[19] ),
    .A2(_08772_),
    .B(_08844_),
    .Y(_08845_));
 BUFx3_ASAP7_75t_R _15955_ (.A(_07515_),
    .Y(_08846_));
 AND2x2_ASAP7_75t_R _15956_ (.A(\dmem.inter_dmem0[19] ),
    .B(_08846_),
    .Y(_08847_));
 AO221x1_ASAP7_75t_R _15957_ (.A1(\dmem.inter_dmem2[19] ),
    .A2(_08771_),
    .B1(_08845_),
    .B2(_08826_),
    .C(_08847_),
    .Y(_08848_));
 AO211x2_ASAP7_75t_R _15958_ (.A1(_08770_),
    .A2(_08848_),
    .B(_08781_),
    .C(_08748_),
    .Y(_08849_));
 BUFx4f_ASAP7_75t_R _15959_ (.A(_08849_),
    .Y(_08850_));
 AO21x2_ASAP7_75t_R _15960_ (.A1(_08172_),
    .A2(_08184_),
    .B(_08662_),
    .Y(_08851_));
 OR2x2_ASAP7_75t_R _15961_ (.A(_01116_),
    .B(_08809_),
    .Y(_08852_));
 OR3x1_ASAP7_75t_R _15962_ (.A(_01119_),
    .B(_08715_),
    .C(_08852_),
    .Y(_08853_));
 XNOR2x1_ASAP7_75t_R _15963_ (.B(_08853_),
    .Y(_08854_),
    .A(_01122_));
 AND3x1_ASAP7_75t_R _15964_ (.A(_01115_),
    .B(_01124_),
    .C(_08837_),
    .Y(_08855_));
 OA211x2_ASAP7_75t_R _15965_ (.A1(_01114_),
    .A2(_01117_),
    .B(_01124_),
    .C(_08837_),
    .Y(_08856_));
 AO21x1_ASAP7_75t_R _15966_ (.A1(_01120_),
    .A2(_01124_),
    .B(_08856_),
    .Y(_08857_));
 AO31x2_ASAP7_75t_R _15967_ (.A1(_08813_),
    .A2(_08815_),
    .A3(_08855_),
    .B(_08857_),
    .Y(_08858_));
 XNOR2x1_ASAP7_75t_R _15968_ (.B(_08858_),
    .Y(_08859_),
    .A(_01123_));
 AOI22x1_ASAP7_75t_R _15969_ (.A1(_08594_),
    .A2(_08854_),
    .B1(_08859_),
    .B2(_08648_),
    .Y(_08860_));
 AND3x1_ASAP7_75t_R _15970_ (.A(_08806_),
    .B(_08851_),
    .C(_08860_),
    .Y(_08861_));
 INVx1_ASAP7_75t_R _15971_ (.A(_00444_),
    .Y(_08862_));
 AO32x1_ASAP7_75t_R _15972_ (.A1(_08799_),
    .A2(_08850_),
    .A3(_08861_),
    .B1(_08796_),
    .B2(_08862_),
    .Y(_01264_));
 OA211x2_ASAP7_75t_R _15973_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08591_),
    .C(\dmem.inter_dmem3[1] ),
    .Y(_08863_));
 AO21x1_ASAP7_75t_R _15974_ (.A1(\dmem.inter_dmem1[1] ),
    .A2(net47),
    .B(_08863_),
    .Y(_08864_));
 AND2x2_ASAP7_75t_R _15975_ (.A(\dmem.inter_dmem0[1] ),
    .B(\dmem.ce_mem[3] ),
    .Y(_08865_));
 AO221x1_ASAP7_75t_R _15976_ (.A1(\dmem.inter_dmem2[1] ),
    .A2(\dmem.ce_mem[1] ),
    .B1(_08864_),
    .B2(_08658_),
    .C(_08865_),
    .Y(_08866_));
 AOI22x1_ASAP7_75t_R _15977_ (.A1(net76),
    .A2(_08570_),
    .B1(_08687_),
    .B2(_08578_),
    .Y(_08867_));
 AND2x2_ASAP7_75t_R _15978_ (.A(_08587_),
    .B(_08867_),
    .Y(_08868_));
 AOI22x1_ASAP7_75t_R _15979_ (.A1(_08732_),
    .A2(_08867_),
    .B1(_08868_),
    .B2(_07726_),
    .Y(_08869_));
 OA21x2_ASAP7_75t_R _15980_ (.A1(_08587_),
    .A2(_08866_),
    .B(_08869_),
    .Y(_08870_));
 BUFx12f_ASAP7_75t_R _15981_ (.A(_08602_),
    .Y(_08871_));
 INVx1_ASAP7_75t_R _15982_ (.A(_01041_),
    .Y(_08872_));
 AO21x1_ASAP7_75t_R _15983_ (.A1(_08871_),
    .A2(_08607_),
    .B(_08872_),
    .Y(_08873_));
 OA21x2_ASAP7_75t_R _15984_ (.A1(_08609_),
    .A2(_08870_),
    .B(_08873_),
    .Y(_01265_));
 OA211x2_ASAP7_75t_R _15985_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[20] ),
    .Y(_08874_));
 AO21x1_ASAP7_75t_R _15986_ (.A1(\dmem.inter_dmem1[20] ),
    .A2(_08772_),
    .B(_08874_),
    .Y(_08875_));
 AND2x2_ASAP7_75t_R _15987_ (.A(\dmem.inter_dmem0[20] ),
    .B(_08846_),
    .Y(_08876_));
 AO221x1_ASAP7_75t_R _15988_ (.A1(\dmem.inter_dmem2[20] ),
    .A2(_08771_),
    .B1(_08875_),
    .B2(_08826_),
    .C(_08876_),
    .Y(_08877_));
 AO211x2_ASAP7_75t_R _15989_ (.A1(_08770_),
    .A2(_08877_),
    .B(_08781_),
    .C(_08748_),
    .Y(_08878_));
 BUFx4f_ASAP7_75t_R _15990_ (.A(_08878_),
    .Y(_08879_));
 NAND2x1_ASAP7_75t_R _15991_ (.A(_07933_),
    .B(_08634_),
    .Y(_08880_));
 OR3x1_ASAP7_75t_R _15992_ (.A(_07933_),
    .B(_08204_),
    .C(_08661_),
    .Y(_08881_));
 OR4x1_ASAP7_75t_R _15993_ (.A(_01111_),
    .B(_01114_),
    .C(_01117_),
    .D(_01120_),
    .Y(_08882_));
 AO21x1_ASAP7_75t_R _15994_ (.A1(_08789_),
    .A2(_08790_),
    .B(_08882_),
    .Y(_08883_));
 OR4x1_ASAP7_75t_R _15995_ (.A(_01115_),
    .B(_01114_),
    .C(_01117_),
    .D(_01120_),
    .Y(_08884_));
 OA21x2_ASAP7_75t_R _15996_ (.A1(_01120_),
    .A2(_08837_),
    .B(_08884_),
    .Y(_08885_));
 AND3x1_ASAP7_75t_R _15997_ (.A(_01124_),
    .B(_08883_),
    .C(_08885_),
    .Y(_08886_));
 OAI21x1_ASAP7_75t_R _15998_ (.A1(_01123_),
    .A2(_08886_),
    .B(_01127_),
    .Y(_08887_));
 XNOR2x1_ASAP7_75t_R _15999_ (.B(_08887_),
    .Y(_08888_),
    .A(_01126_));
 OR4x1_ASAP7_75t_R _16000_ (.A(_01119_),
    .B(_01122_),
    .C(_08650_),
    .D(_08852_),
    .Y(_08889_));
 XNOR2x1_ASAP7_75t_R _16001_ (.B(_08889_),
    .Y(_08890_),
    .A(net77));
 OA22x2_ASAP7_75t_R _16002_ (.A1(_08394_),
    .A2(_08888_),
    .B1(_08890_),
    .B2(_08583_),
    .Y(_08891_));
 OA211x2_ASAP7_75t_R _16003_ (.A1(_08195_),
    .A2(_08880_),
    .B(_08881_),
    .C(_08891_),
    .Y(_08892_));
 AND2x2_ASAP7_75t_R _16004_ (.A(_08806_),
    .B(_08892_),
    .Y(_08893_));
 INVx1_ASAP7_75t_R _16005_ (.A(_00411_),
    .Y(_08894_));
 AO32x1_ASAP7_75t_R _16006_ (.A1(_08799_),
    .A2(_08879_),
    .A3(_08893_),
    .B1(_08796_),
    .B2(_08894_),
    .Y(_01266_));
 BUFx3_ASAP7_75t_R _16007_ (.A(_07465_),
    .Y(_08895_));
 OA211x2_ASAP7_75t_R _16008_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[21] ),
    .Y(_08896_));
 AO21x1_ASAP7_75t_R _16009_ (.A1(\dmem.inter_dmem1[21] ),
    .A2(_08772_),
    .B(_08896_),
    .Y(_08897_));
 AND2x2_ASAP7_75t_R _16010_ (.A(\dmem.inter_dmem0[21] ),
    .B(_08846_),
    .Y(_08898_));
 AO221x1_ASAP7_75t_R _16011_ (.A1(\dmem.inter_dmem2[21] ),
    .A2(_08771_),
    .B1(_08897_),
    .B2(_08826_),
    .C(_08898_),
    .Y(_08899_));
 AO211x2_ASAP7_75t_R _16012_ (.A1(_08770_),
    .A2(_08899_),
    .B(_08781_),
    .C(_08748_),
    .Y(_08900_));
 BUFx4f_ASAP7_75t_R _16013_ (.A(_08900_),
    .Y(_08901_));
 OR2x6_ASAP7_75t_R _16014_ (.A(net45),
    .B(_08661_),
    .Y(_08902_));
 OR4x2_ASAP7_75t_R _16015_ (.A(_01119_),
    .B(_01122_),
    .C(_01125_),
    .D(_08852_),
    .Y(_08903_));
 NOR2x1_ASAP7_75t_R _16016_ (.A(_08715_),
    .B(_08903_),
    .Y(_08904_));
 XNOR2x1_ASAP7_75t_R _16017_ (.B(_08904_),
    .Y(_08905_),
    .A(net78));
 OR2x2_ASAP7_75t_R _16018_ (.A(_01123_),
    .B(_01126_),
    .Y(_08906_));
 OA21x2_ASAP7_75t_R _16019_ (.A1(_01127_),
    .A2(_01126_),
    .B(_01130_),
    .Y(_08907_));
 OA21x2_ASAP7_75t_R _16020_ (.A1(_08858_),
    .A2(_08906_),
    .B(_08907_),
    .Y(_08908_));
 XNOR2x1_ASAP7_75t_R _16021_ (.B(_08908_),
    .Y(_08909_),
    .A(_01129_));
 AOI22x1_ASAP7_75t_R _16022_ (.A1(_08594_),
    .A2(_08905_),
    .B1(_08909_),
    .B2(_08648_),
    .Y(_08910_));
 AND3x1_ASAP7_75t_R _16023_ (.A(_08806_),
    .B(_08902_),
    .C(_08910_),
    .Y(_08911_));
 INVx1_ASAP7_75t_R _16024_ (.A(_00378_),
    .Y(_08912_));
 AO32x1_ASAP7_75t_R _16025_ (.A1(_08799_),
    .A2(_08901_),
    .A3(_08911_),
    .B1(_08796_),
    .B2(_08912_),
    .Y(_01267_));
 OA211x2_ASAP7_75t_R _16026_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[22] ),
    .Y(_08913_));
 AO21x1_ASAP7_75t_R _16027_ (.A1(\dmem.inter_dmem1[22] ),
    .A2(_08772_),
    .B(_08913_),
    .Y(_08914_));
 AND2x2_ASAP7_75t_R _16028_ (.A(\dmem.inter_dmem0[22] ),
    .B(_08846_),
    .Y(_08915_));
 AO221x1_ASAP7_75t_R _16029_ (.A1(\dmem.inter_dmem2[22] ),
    .A2(_08771_),
    .B1(_08914_),
    .B2(_08826_),
    .C(_08915_),
    .Y(_08916_));
 AO211x2_ASAP7_75t_R _16030_ (.A1(_08770_),
    .A2(_08916_),
    .B(_08781_),
    .C(_08747_),
    .Y(_08917_));
 BUFx3_ASAP7_75t_R _16031_ (.A(_08917_),
    .Y(_08918_));
 AND2x2_ASAP7_75t_R _16032_ (.A(_08883_),
    .B(_08885_),
    .Y(_08919_));
 AND3x1_ASAP7_75t_R _16033_ (.A(_01124_),
    .B(_01127_),
    .C(_01130_),
    .Y(_08920_));
 AND3x1_ASAP7_75t_R _16034_ (.A(_01123_),
    .B(_01127_),
    .C(_01130_),
    .Y(_08921_));
 AO221x1_ASAP7_75t_R _16035_ (.A1(_01126_),
    .A2(_01130_),
    .B1(_08919_),
    .B2(_08920_),
    .C(_08921_),
    .Y(_08922_));
 OA21x2_ASAP7_75t_R _16036_ (.A1(_01129_),
    .A2(_08922_),
    .B(_01133_),
    .Y(_08923_));
 XNOR2x1_ASAP7_75t_R _16037_ (.B(_08923_),
    .Y(_08924_),
    .A(_01132_));
 NAND2x1_ASAP7_75t_R _16038_ (.A(_08687_),
    .B(_08924_),
    .Y(_08925_));
 OR3x1_ASAP7_75t_R _16039_ (.A(_01128_),
    .B(_08651_),
    .C(_08903_),
    .Y(_08926_));
 XNOR2x1_ASAP7_75t_R _16040_ (.B(_08926_),
    .Y(_08927_),
    .A(_01131_));
 AOI22x1_ASAP7_75t_R _16041_ (.A1(_08237_),
    .A2(_08634_),
    .B1(_08927_),
    .B2(_08569_),
    .Y(_08928_));
 OA211x2_ASAP7_75t_R _16042_ (.A1(_08248_),
    .A2(_08662_),
    .B(_08925_),
    .C(_08928_),
    .Y(_08929_));
 AND2x2_ASAP7_75t_R _16043_ (.A(_08806_),
    .B(_08929_),
    .Y(_08930_));
 INVx1_ASAP7_75t_R _16044_ (.A(_00345_),
    .Y(_08931_));
 AO32x1_ASAP7_75t_R _16045_ (.A1(_08799_),
    .A2(_08918_),
    .A3(_08930_),
    .B1(_08796_),
    .B2(_08931_),
    .Y(_01268_));
 OA211x2_ASAP7_75t_R _16046_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[23] ),
    .Y(_08932_));
 AO21x1_ASAP7_75t_R _16047_ (.A1(\dmem.inter_dmem1[23] ),
    .A2(_08772_),
    .B(_08932_),
    .Y(_08933_));
 AND2x2_ASAP7_75t_R _16048_ (.A(\dmem.inter_dmem0[23] ),
    .B(_08846_),
    .Y(_08934_));
 AO221x1_ASAP7_75t_R _16049_ (.A1(\dmem.inter_dmem2[23] ),
    .A2(_08771_),
    .B1(_08933_),
    .B2(_08826_),
    .C(_08934_),
    .Y(_08935_));
 AO211x2_ASAP7_75t_R _16050_ (.A1(_08770_),
    .A2(_08935_),
    .B(_08781_),
    .C(_08747_),
    .Y(_08936_));
 BUFx4f_ASAP7_75t_R _16051_ (.A(_08936_),
    .Y(_08937_));
 OA21x2_ASAP7_75t_R _16052_ (.A1(_01129_),
    .A2(_08908_),
    .B(_01133_),
    .Y(_08938_));
 OA21x2_ASAP7_75t_R _16053_ (.A1(_01132_),
    .A2(_08938_),
    .B(_01136_),
    .Y(_08939_));
 XOR2x1_ASAP7_75t_R _16054_ (.A(_01135_),
    .Y(_08940_),
    .B(_08939_));
 OR4x1_ASAP7_75t_R _16055_ (.A(_01128_),
    .B(_01131_),
    .C(_08715_),
    .D(_08903_),
    .Y(_08941_));
 XNOR2x1_ASAP7_75t_R _16056_ (.B(_08941_),
    .Y(_08942_),
    .A(net80));
 OA222x2_ASAP7_75t_R _16057_ (.A1(net47),
    .A2(_08662_),
    .B1(_08940_),
    .B2(_08394_),
    .C1(_08942_),
    .C2(_08583_),
    .Y(_08943_));
 AND2x2_ASAP7_75t_R _16058_ (.A(_08806_),
    .B(_08943_),
    .Y(_08944_));
 INVx1_ASAP7_75t_R _16059_ (.A(_00311_),
    .Y(_08945_));
 AO32x1_ASAP7_75t_R _16060_ (.A1(_08799_),
    .A2(_08937_),
    .A3(_08944_),
    .B1(_08796_),
    .B2(_08945_),
    .Y(_01269_));
 OA211x2_ASAP7_75t_R _16061_ (.A1(_08617_),
    .A2(_08620_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[24] ),
    .Y(_08946_));
 AO21x1_ASAP7_75t_R _16062_ (.A1(\dmem.inter_dmem1[24] ),
    .A2(_08772_),
    .B(_08946_),
    .Y(_08947_));
 AND2x2_ASAP7_75t_R _16063_ (.A(\dmem.inter_dmem0[24] ),
    .B(_08846_),
    .Y(_08948_));
 AO221x1_ASAP7_75t_R _16064_ (.A1(\dmem.inter_dmem2[24] ),
    .A2(_08771_),
    .B1(_08947_),
    .B2(_08826_),
    .C(_08948_),
    .Y(_08949_));
 AO211x2_ASAP7_75t_R _16065_ (.A1(_08770_),
    .A2(_08949_),
    .B(_08781_),
    .C(_08747_),
    .Y(_08950_));
 BUFx4f_ASAP7_75t_R _16066_ (.A(_08950_),
    .Y(_08951_));
 OR3x1_ASAP7_75t_R _16067_ (.A(_01129_),
    .B(_01132_),
    .C(_01135_),
    .Y(_08952_));
 OR2x2_ASAP7_75t_R _16068_ (.A(_01133_),
    .B(_01132_),
    .Y(_08953_));
 AO21x1_ASAP7_75t_R _16069_ (.A1(_01136_),
    .A2(_08953_),
    .B(_01135_),
    .Y(_08954_));
 OA21x2_ASAP7_75t_R _16070_ (.A1(_08922_),
    .A2(_08952_),
    .B(_08954_),
    .Y(_08955_));
 AND2x2_ASAP7_75t_R _16071_ (.A(_01139_),
    .B(_08955_),
    .Y(_08956_));
 XNOR2x2_ASAP7_75t_R _16072_ (.A(_01138_),
    .B(_08956_),
    .Y(_08957_));
 OR4x2_ASAP7_75t_R _16073_ (.A(_01128_),
    .B(_01131_),
    .C(_01134_),
    .D(_08903_),
    .Y(_08958_));
 NOR2x1_ASAP7_75t_R _16074_ (.A(_08651_),
    .B(_08958_),
    .Y(_08959_));
 XNOR2x1_ASAP7_75t_R _16075_ (.B(_08959_),
    .Y(_08960_),
    .A(net81));
 AOI22x1_ASAP7_75t_R _16076_ (.A1(_08687_),
    .A2(_08957_),
    .B1(_08960_),
    .B2(_08570_),
    .Y(_08961_));
 OA21x2_ASAP7_75t_R _16077_ (.A1(net48),
    .A2(_08662_),
    .B(_08961_),
    .Y(_08962_));
 AND2x2_ASAP7_75t_R _16078_ (.A(_08806_),
    .B(_08962_),
    .Y(_08963_));
 INVx1_ASAP7_75t_R _16079_ (.A(_00278_),
    .Y(_08964_));
 AO32x1_ASAP7_75t_R _16080_ (.A1(_08799_),
    .A2(_08951_),
    .A3(_08963_),
    .B1(_08796_),
    .B2(_08964_),
    .Y(_01270_));
 OA211x2_ASAP7_75t_R _16081_ (.A1(_08617_),
    .A2(_08620_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[25] ),
    .Y(_08965_));
 AO21x1_ASAP7_75t_R _16082_ (.A1(\dmem.inter_dmem1[25] ),
    .A2(_07417_),
    .B(_08965_),
    .Y(_08966_));
 AND2x2_ASAP7_75t_R _16083_ (.A(\dmem.inter_dmem0[25] ),
    .B(_08846_),
    .Y(_08967_));
 AO221x1_ASAP7_75t_R _16084_ (.A1(\dmem.inter_dmem2[25] ),
    .A2(_08771_),
    .B1(_08966_),
    .B2(_08826_),
    .C(_08967_),
    .Y(_08968_));
 AO211x2_ASAP7_75t_R _16085_ (.A1(_08769_),
    .A2(_08968_),
    .B(_08780_),
    .C(_08747_),
    .Y(_08969_));
 BUFx4f_ASAP7_75t_R _16086_ (.A(_08969_),
    .Y(_08970_));
 OR2x2_ASAP7_75t_R _16087_ (.A(_01135_),
    .B(_08939_),
    .Y(_08971_));
 AO21x1_ASAP7_75t_R _16088_ (.A1(_01139_),
    .A2(_08971_),
    .B(_01138_),
    .Y(_08972_));
 AND2x2_ASAP7_75t_R _16089_ (.A(_01142_),
    .B(_08972_),
    .Y(_08973_));
 XNOR2x2_ASAP7_75t_R _16090_ (.A(_01141_),
    .B(_08973_),
    .Y(_08974_));
 OR3x1_ASAP7_75t_R _16091_ (.A(_01137_),
    .B(_08715_),
    .C(_08958_),
    .Y(_08975_));
 XNOR2x1_ASAP7_75t_R _16092_ (.B(_08975_),
    .Y(_08976_),
    .A(net82));
 INVx1_ASAP7_75t_R _16093_ (.A(_08976_),
    .Y(_08977_));
 AOI22x1_ASAP7_75t_R _16094_ (.A1(_08687_),
    .A2(_08974_),
    .B1(_08977_),
    .B2(_08570_),
    .Y(_08978_));
 OA21x2_ASAP7_75t_R _16095_ (.A1(net49),
    .A2(_08662_),
    .B(_08978_),
    .Y(_08979_));
 AND2x2_ASAP7_75t_R _16096_ (.A(_08699_),
    .B(_08979_),
    .Y(_08980_));
 INVx1_ASAP7_75t_R _16097_ (.A(_00245_),
    .Y(_08981_));
 AO32x1_ASAP7_75t_R _16098_ (.A1(_08799_),
    .A2(_08970_),
    .A3(_08980_),
    .B1(_08796_),
    .B2(_08981_),
    .Y(_01271_));
 OA211x2_ASAP7_75t_R _16099_ (.A1(_08617_),
    .A2(_08620_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[26] ),
    .Y(_08982_));
 AO21x1_ASAP7_75t_R _16100_ (.A1(\dmem.inter_dmem1[26] ),
    .A2(_07417_),
    .B(_08982_),
    .Y(_08983_));
 AND2x2_ASAP7_75t_R _16101_ (.A(\dmem.inter_dmem0[26] ),
    .B(_08846_),
    .Y(_08984_));
 AO221x1_ASAP7_75t_R _16102_ (.A1(\dmem.inter_dmem2[26] ),
    .A2(_08614_),
    .B1(_08983_),
    .B2(_08826_),
    .C(_08984_),
    .Y(_08985_));
 AO211x2_ASAP7_75t_R _16103_ (.A1(_08769_),
    .A2(_08985_),
    .B(_08780_),
    .C(_08747_),
    .Y(_08986_));
 BUFx4f_ASAP7_75t_R _16104_ (.A(_08986_),
    .Y(_08987_));
 AND3x1_ASAP7_75t_R _16105_ (.A(_01139_),
    .B(_01142_),
    .C(_01145_),
    .Y(_08988_));
 AND3x1_ASAP7_75t_R _16106_ (.A(_01138_),
    .B(_01142_),
    .C(_01145_),
    .Y(_08989_));
 AO21x1_ASAP7_75t_R _16107_ (.A1(_01141_),
    .A2(_01145_),
    .B(_08989_),
    .Y(_08990_));
 AO21x1_ASAP7_75t_R _16108_ (.A1(_08955_),
    .A2(_08988_),
    .B(_08990_),
    .Y(_08991_));
 XNOR2x1_ASAP7_75t_R _16109_ (.B(_08991_),
    .Y(_08992_),
    .A(_01144_));
 OR3x2_ASAP7_75t_R _16110_ (.A(_01137_),
    .B(_01140_),
    .C(_08958_),
    .Y(_08993_));
 NOR2x1_ASAP7_75t_R _16111_ (.A(_08651_),
    .B(_08993_),
    .Y(_08994_));
 XNOR2x1_ASAP7_75t_R _16112_ (.B(_08994_),
    .Y(_08995_),
    .A(net83));
 AO222x2_ASAP7_75t_R _16113_ (.A1(_08311_),
    .A2(_08634_),
    .B1(_08992_),
    .B2(_08648_),
    .C1(_08995_),
    .C2(_08570_),
    .Y(_08996_));
 BUFx10_ASAP7_75t_R _16114_ (.A(_08996_),
    .Y(_08997_));
 NOR2x1_ASAP7_75t_R _16115_ (.A(_08726_),
    .B(_08997_),
    .Y(_08998_));
 INVx1_ASAP7_75t_R _16116_ (.A(_00212_),
    .Y(_08999_));
 AO32x1_ASAP7_75t_R _16117_ (.A1(_08799_),
    .A2(_08987_),
    .A3(_08998_),
    .B1(_08726_),
    .B2(_08999_),
    .Y(_01272_));
 INVx1_ASAP7_75t_R _16118_ (.A(_00178_),
    .Y(_09000_));
 OA211x2_ASAP7_75t_R _16119_ (.A1(_08773_),
    .A2(_08774_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[27] ),
    .Y(_09001_));
 AO21x1_ASAP7_75t_R _16120_ (.A1(\dmem.inter_dmem1[27] ),
    .A2(net47),
    .B(_09001_),
    .Y(_09002_));
 AND2x2_ASAP7_75t_R _16121_ (.A(\dmem.inter_dmem0[27] ),
    .B(_08628_),
    .Y(_09003_));
 AO221x1_ASAP7_75t_R _16122_ (.A1(\dmem.inter_dmem2[27] ),
    .A2(\dmem.ce_mem[1] ),
    .B1(_09002_),
    .B2(_08658_),
    .C(_09003_),
    .Y(_09004_));
 AO211x2_ASAP7_75t_R _16123_ (.A1(_08770_),
    .A2(_09004_),
    .B(_08781_),
    .C(_08748_),
    .Y(_09005_));
 BUFx4f_ASAP7_75t_R _16124_ (.A(_09005_),
    .Y(_09006_));
 AO21x1_ASAP7_75t_R _16125_ (.A1(\dmem.inter_dmem0[7] ),
    .A2(_08628_),
    .B(_08612_),
    .Y(_09007_));
 OR3x1_ASAP7_75t_R _16126_ (.A(_01143_),
    .B(_08715_),
    .C(_08993_),
    .Y(_09008_));
 XNOR2x1_ASAP7_75t_R _16127_ (.B(_09008_),
    .Y(_09009_),
    .A(_01146_));
 NAND2x1_ASAP7_75t_R _16128_ (.A(_08569_),
    .B(_09009_),
    .Y(_09010_));
 OA21x2_ASAP7_75t_R _16129_ (.A1(_03562_),
    .A2(_08630_),
    .B(_09010_),
    .Y(_09011_));
 OA21x2_ASAP7_75t_R _16130_ (.A1(net51),
    .A2(_08661_),
    .B(_09011_),
    .Y(_09012_));
 AO21x1_ASAP7_75t_R _16131_ (.A1(_08971_),
    .A2(_08988_),
    .B(_08990_),
    .Y(_09013_));
 OA21x2_ASAP7_75t_R _16132_ (.A1(_01144_),
    .A2(_09013_),
    .B(_01148_),
    .Y(_09014_));
 XNOR2x2_ASAP7_75t_R _16133_ (.A(_01147_),
    .B(_09014_),
    .Y(_09015_));
 NAND2x1_ASAP7_75t_R _16134_ (.A(_08687_),
    .B(_09015_),
    .Y(_09016_));
 OA211x2_ASAP7_75t_R _16135_ (.A1(_08627_),
    .A2(_09007_),
    .B(_09012_),
    .C(_09016_),
    .Y(_09017_));
 AND2x2_ASAP7_75t_R _16136_ (.A(_08700_),
    .B(_09017_),
    .Y(_09018_));
 AO22x1_ASAP7_75t_R _16137_ (.A1(_09000_),
    .A2(_08610_),
    .B1(_09006_),
    .B2(_09018_),
    .Y(_01273_));
 BUFx4f_ASAP7_75t_R _16138_ (.A(_08798_),
    .Y(_09019_));
 OA211x2_ASAP7_75t_R _16139_ (.A1(_08617_),
    .A2(_08620_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[28] ),
    .Y(_09020_));
 AO21x1_ASAP7_75t_R _16140_ (.A1(\dmem.inter_dmem1[28] ),
    .A2(_07417_),
    .B(_09020_),
    .Y(_09021_));
 AND2x2_ASAP7_75t_R _16141_ (.A(\dmem.inter_dmem0[28] ),
    .B(_08846_),
    .Y(_09022_));
 AO221x1_ASAP7_75t_R _16142_ (.A1(\dmem.inter_dmem2[28] ),
    .A2(_08614_),
    .B1(_09021_),
    .B2(_08826_),
    .C(_09022_),
    .Y(_09023_));
 AO211x2_ASAP7_75t_R _16143_ (.A1(_08769_),
    .A2(_09023_),
    .B(_08780_),
    .C(_08747_),
    .Y(_09024_));
 BUFx3_ASAP7_75t_R _16144_ (.A(_09024_),
    .Y(_09025_));
 OR2x2_ASAP7_75t_R _16145_ (.A(_01144_),
    .B(_01147_),
    .Y(_09026_));
 OA21x2_ASAP7_75t_R _16146_ (.A1(_01148_),
    .A2(_01147_),
    .B(_01151_),
    .Y(_09027_));
 OA21x2_ASAP7_75t_R _16147_ (.A1(_08991_),
    .A2(_09026_),
    .B(_09027_),
    .Y(_09028_));
 XNOR2x2_ASAP7_75t_R _16148_ (.A(_01150_),
    .B(_09028_),
    .Y(_09029_));
 NAND2x2_ASAP7_75t_R _16149_ (.A(_08687_),
    .B(_09029_),
    .Y(_09030_));
 OR2x6_ASAP7_75t_R _16150_ (.A(net52),
    .B(_08661_),
    .Y(_09031_));
 OR2x2_ASAP7_75t_R _16151_ (.A(_01143_),
    .B(_08993_),
    .Y(_09032_));
 OR3x1_ASAP7_75t_R _16152_ (.A(_01146_),
    .B(_08651_),
    .C(_09032_),
    .Y(_09033_));
 XNOR2x1_ASAP7_75t_R _16153_ (.B(_09033_),
    .Y(_09034_),
    .A(net85));
 OR2x6_ASAP7_75t_R _16154_ (.A(_08583_),
    .B(_09034_),
    .Y(_09035_));
 AND4x1_ASAP7_75t_R _16155_ (.A(_08699_),
    .B(_09030_),
    .C(_09031_),
    .D(_09035_),
    .Y(_09036_));
 INVx1_ASAP7_75t_R _16156_ (.A(_00145_),
    .Y(_09037_));
 AO32x1_ASAP7_75t_R _16157_ (.A1(_09019_),
    .A2(_09025_),
    .A3(_09036_),
    .B1(_08726_),
    .B2(_09037_),
    .Y(_01274_));
 OA211x2_ASAP7_75t_R _16158_ (.A1(_08617_),
    .A2(_08620_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[29] ),
    .Y(_09038_));
 AO21x1_ASAP7_75t_R _16159_ (.A1(\dmem.inter_dmem1[29] ),
    .A2(_07417_),
    .B(_09038_),
    .Y(_09039_));
 AND2x2_ASAP7_75t_R _16160_ (.A(\dmem.inter_dmem0[29] ),
    .B(_08846_),
    .Y(_09040_));
 AO221x1_ASAP7_75t_R _16161_ (.A1(\dmem.inter_dmem2[29] ),
    .A2(_08614_),
    .B1(_09039_),
    .B2(_08585_),
    .C(_09040_),
    .Y(_09041_));
 AO211x2_ASAP7_75t_R _16162_ (.A1(_08769_),
    .A2(_09041_),
    .B(_08780_),
    .C(_08747_),
    .Y(_09042_));
 BUFx4f_ASAP7_75t_R _16163_ (.A(_09042_),
    .Y(_09043_));
 OR3x1_ASAP7_75t_R _16164_ (.A(_01144_),
    .B(_01147_),
    .C(_01150_),
    .Y(_09044_));
 OA21x2_ASAP7_75t_R _16165_ (.A1(_01150_),
    .A2(_09027_),
    .B(_01154_),
    .Y(_09045_));
 OA21x2_ASAP7_75t_R _16166_ (.A1(_09013_),
    .A2(_09044_),
    .B(_09045_),
    .Y(_09046_));
 XNOR2x2_ASAP7_75t_R _16167_ (.A(_01153_),
    .B(_09046_),
    .Y(_09047_));
 NAND2x2_ASAP7_75t_R _16168_ (.A(_08648_),
    .B(_09047_),
    .Y(_09048_));
 OR4x2_ASAP7_75t_R _16169_ (.A(_01146_),
    .B(_01149_),
    .C(_08715_),
    .D(_09032_),
    .Y(_09049_));
 XNOR2x1_ASAP7_75t_R _16170_ (.B(_09049_),
    .Y(_09050_),
    .A(net86));
 OA22x2_ASAP7_75t_R _16171_ (.A1(net53),
    .A2(_08662_),
    .B1(_09050_),
    .B2(_08583_),
    .Y(_09051_));
 AND3x1_ASAP7_75t_R _16172_ (.A(_08806_),
    .B(_09048_),
    .C(_09051_),
    .Y(_09052_));
 INVx1_ASAP7_75t_R _16173_ (.A(_00111_),
    .Y(_09053_));
 AO32x1_ASAP7_75t_R _16174_ (.A1(_09019_),
    .A2(_09043_),
    .A3(_09052_),
    .B1(_08726_),
    .B2(_09053_),
    .Y(_01275_));
 XOR2x1_ASAP7_75t_R _16175_ (.A(_01073_),
    .Y(_09054_),
    .B(_01160_));
 AO32x1_ASAP7_75t_R _16176_ (.A1(_04849_),
    .A2(_08390_),
    .A3(_09054_),
    .B1(_08569_),
    .B2(_10109_),
    .Y(_09055_));
 AND2x2_ASAP7_75t_R _16177_ (.A(\dmem.inter_dmem0[2] ),
    .B(_07515_),
    .Y(_09056_));
 AND3x1_ASAP7_75t_R _16178_ (.A(\dmem.inter_dmem1[2] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_09057_));
 OA211x2_ASAP7_75t_R _16179_ (.A1(_08617_),
    .A2(_08620_),
    .B(_07465_),
    .C(\dmem.inter_dmem3[2] ),
    .Y(_09058_));
 OA21x2_ASAP7_75t_R _16180_ (.A1(_09057_),
    .A2(_09058_),
    .B(_08585_),
    .Y(_09059_));
 AND4x1_ASAP7_75t_R _16181_ (.A(\dmem.inter_dmem2[2] ),
    .B(_07416_),
    .C(net38),
    .D(_08589_),
    .Y(_09060_));
 OR4x1_ASAP7_75t_R _16182_ (.A(_08587_),
    .B(_09056_),
    .C(_09059_),
    .D(_09060_),
    .Y(_09061_));
 OR3x1_ASAP7_75t_R _16183_ (.A(_08580_),
    .B(net54),
    .C(_09055_),
    .Y(_09062_));
 OA211x2_ASAP7_75t_R _16184_ (.A1(_08584_),
    .A2(_09055_),
    .B(_09061_),
    .C(_09062_),
    .Y(_09063_));
 NAND2x1_ASAP7_75t_R _16185_ (.A(_01008_),
    .B(_08610_),
    .Y(_09064_));
 OA21x2_ASAP7_75t_R _16186_ (.A1(_08609_),
    .A2(_09063_),
    .B(_09064_),
    .Y(_01276_));
 OA211x2_ASAP7_75t_R _16187_ (.A1(_08617_),
    .A2(_08620_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[30] ),
    .Y(_09065_));
 AO21x1_ASAP7_75t_R _16188_ (.A1(\dmem.inter_dmem1[30] ),
    .A2(_07417_),
    .B(_09065_),
    .Y(_09066_));
 AND2x2_ASAP7_75t_R _16189_ (.A(\dmem.inter_dmem0[30] ),
    .B(_07515_),
    .Y(_09067_));
 AO221x1_ASAP7_75t_R _16190_ (.A1(\dmem.inter_dmem2[30] ),
    .A2(_08614_),
    .B1(_09066_),
    .B2(_08585_),
    .C(_09067_),
    .Y(_09068_));
 AO211x2_ASAP7_75t_R _16191_ (.A1(_08769_),
    .A2(_09068_),
    .B(_08780_),
    .C(_08747_),
    .Y(_09069_));
 BUFx4f_ASAP7_75t_R _16192_ (.A(_09069_),
    .Y(_09070_));
 OA21x2_ASAP7_75t_R _16193_ (.A1(_01150_),
    .A2(_09028_),
    .B(_01154_),
    .Y(_09071_));
 OA21x2_ASAP7_75t_R _16194_ (.A1(_01153_),
    .A2(_09071_),
    .B(_01157_),
    .Y(_09072_));
 XNOR2x2_ASAP7_75t_R _16195_ (.A(_01156_),
    .B(_09072_),
    .Y(_09073_));
 NAND2x2_ASAP7_75t_R _16196_ (.A(_08687_),
    .B(_09073_),
    .Y(_09074_));
 OR5x1_ASAP7_75t_R _16197_ (.A(_01146_),
    .B(_01149_),
    .C(_01152_),
    .D(_08651_),
    .E(_09032_),
    .Y(_09075_));
 XNOR2x1_ASAP7_75t_R _16198_ (.B(_09075_),
    .Y(_09076_),
    .A(net88));
 OR2x6_ASAP7_75t_R _16199_ (.A(_08583_),
    .B(_09076_),
    .Y(_09077_));
 OAI21x1_ASAP7_75t_R _16200_ (.A1(_08381_),
    .A2(_08388_),
    .B(_08634_),
    .Y(_09078_));
 AND4x1_ASAP7_75t_R _16201_ (.A(_08699_),
    .B(_09074_),
    .C(_09077_),
    .D(_09078_),
    .Y(_09079_));
 INVx1_ASAP7_75t_R _16202_ (.A(_00077_),
    .Y(_09080_));
 AO32x1_ASAP7_75t_R _16203_ (.A1(_09019_),
    .A2(_09070_),
    .A3(_09079_),
    .B1(_08726_),
    .B2(_09080_),
    .Y(_01277_));
 OA211x2_ASAP7_75t_R _16204_ (.A1(_08617_),
    .A2(_08620_),
    .B(_08895_),
    .C(\dmem.inter_dmem3[31] ),
    .Y(_09081_));
 AO21x1_ASAP7_75t_R _16205_ (.A1(\dmem.inter_dmem1[31] ),
    .A2(_07417_),
    .B(_09081_),
    .Y(_09082_));
 AND2x2_ASAP7_75t_R _16206_ (.A(\dmem.inter_dmem0[31] ),
    .B(_07515_),
    .Y(_09083_));
 AO221x1_ASAP7_75t_R _16207_ (.A1(\dmem.inter_dmem2[31] ),
    .A2(_08614_),
    .B1(_09082_),
    .B2(_08585_),
    .C(_09083_),
    .Y(_09084_));
 AO211x2_ASAP7_75t_R _16208_ (.A1(_08769_),
    .A2(_09084_),
    .B(_08780_),
    .C(_08747_),
    .Y(_09085_));
 BUFx3_ASAP7_75t_R _16209_ (.A(_09085_),
    .Y(_09086_));
 OR3x1_ASAP7_75t_R _16210_ (.A(_01150_),
    .B(_01153_),
    .C(_09026_),
    .Y(_09087_));
 OA21x2_ASAP7_75t_R _16211_ (.A1(_01153_),
    .A2(_09045_),
    .B(_01157_),
    .Y(_09088_));
 OA21x2_ASAP7_75t_R _16212_ (.A1(_09013_),
    .A2(_09087_),
    .B(_09088_),
    .Y(_09089_));
 OA21x2_ASAP7_75t_R _16213_ (.A1(_01156_),
    .A2(_09089_),
    .B(_01158_),
    .Y(_09090_));
 AND2x2_ASAP7_75t_R _16214_ (.A(_09955_),
    .B(_08395_),
    .Y(_09091_));
 XNOR2x1_ASAP7_75t_R _16215_ (.B(_09091_),
    .Y(_09092_),
    .A(_04062_));
 XNOR2x2_ASAP7_75t_R _16216_ (.A(_09090_),
    .B(_09092_),
    .Y(_09093_));
 OR2x6_ASAP7_75t_R _16217_ (.A(_08394_),
    .B(_09093_),
    .Y(_09094_));
 OR3x1_ASAP7_75t_R _16218_ (.A(_01152_),
    .B(_01155_),
    .C(_09049_),
    .Y(_09095_));
 XNOR2x1_ASAP7_75t_R _16219_ (.B(_09095_),
    .Y(_09096_),
    .A(_04072_));
 AOI22x1_ASAP7_75t_R _16220_ (.A1(_08658_),
    .A2(_08634_),
    .B1(_09096_),
    .B2(_08594_),
    .Y(_09097_));
 AND3x1_ASAP7_75t_R _16221_ (.A(_08806_),
    .B(_09094_),
    .C(_09097_),
    .Y(_09098_));
 INVx1_ASAP7_75t_R _16222_ (.A(_00045_),
    .Y(_09099_));
 AO32x1_ASAP7_75t_R _16223_ (.A1(_09019_),
    .A2(_09086_),
    .A3(_09098_),
    .B1(_08726_),
    .B2(_09099_),
    .Y(_01278_));
 OA211x2_ASAP7_75t_R _16224_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[3] ),
    .Y(_09100_));
 AO21x1_ASAP7_75t_R _16225_ (.A1(\dmem.inter_dmem1[3] ),
    .A2(net47),
    .B(_09100_),
    .Y(_09101_));
 AND2x2_ASAP7_75t_R _16226_ (.A(\dmem.inter_dmem0[3] ),
    .B(_08628_),
    .Y(_09102_));
 AO221x1_ASAP7_75t_R _16227_ (.A1(\dmem.inter_dmem2[3] ),
    .A2(\dmem.ce_mem[1] ),
    .B1(_09101_),
    .B2(_08658_),
    .C(_09102_),
    .Y(_09103_));
 XOR2x1_ASAP7_75t_R _16228_ (.A(_01075_),
    .Y(_09104_),
    .B(_08664_));
 INVx1_ASAP7_75t_R _16229_ (.A(_01217_),
    .Y(_09105_));
 AO32x1_ASAP7_75t_R _16230_ (.A1(_04849_),
    .A2(_08390_),
    .A3(_09104_),
    .B1(_08569_),
    .B2(_09105_),
    .Y(_09106_));
 OR2x2_ASAP7_75t_R _16231_ (.A(_08584_),
    .B(_09106_),
    .Y(_09107_));
 OR3x1_ASAP7_75t_R _16232_ (.A(_08580_),
    .B(net57),
    .C(_09106_),
    .Y(_09108_));
 OA211x2_ASAP7_75t_R _16233_ (.A1(_08587_),
    .A2(_09103_),
    .B(_09107_),
    .C(_09108_),
    .Y(_09109_));
 NAND2x1_ASAP7_75t_R _16234_ (.A(_00975_),
    .B(_08610_),
    .Y(_09110_));
 OA21x2_ASAP7_75t_R _16235_ (.A1(_08609_),
    .A2(_09109_),
    .B(_09110_),
    .Y(_01279_));
 AND2x2_ASAP7_75t_R _16236_ (.A(_07416_),
    .B(_08589_),
    .Y(_09111_));
 OR2x2_ASAP7_75t_R _16237_ (.A(\dmem.inter_dmem0[4] ),
    .B(_08589_),
    .Y(_09112_));
 AND3x1_ASAP7_75t_R _16238_ (.A(\dmem.inter_dmem1[4] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_09113_));
 OA211x2_ASAP7_75t_R _16239_ (.A1(_08773_),
    .A2(_08774_),
    .B(net38),
    .C(\dmem.inter_dmem2[4] ),
    .Y(_09114_));
 OR3x1_ASAP7_75t_R _16240_ (.A(_08628_),
    .B(_09113_),
    .C(_09114_),
    .Y(_09115_));
 AO32x1_ASAP7_75t_R _16241_ (.A1(\dmem.inter_dmem3[4] ),
    .A2(_08591_),
    .A3(_09111_),
    .B1(_09112_),
    .B2(_09115_),
    .Y(_09116_));
 XOR2x1_ASAP7_75t_R _16242_ (.A(_01078_),
    .Y(_09117_),
    .B(_08636_));
 XOR2x1_ASAP7_75t_R _16243_ (.A(_01077_),
    .Y(_09118_),
    .B(_01218_));
 AO32x1_ASAP7_75t_R _16244_ (.A1(_04848_),
    .A2(_08390_),
    .A3(_09117_),
    .B1(_09118_),
    .B2(_08569_),
    .Y(_09119_));
 OR2x2_ASAP7_75t_R _16245_ (.A(_08584_),
    .B(_09119_),
    .Y(_09120_));
 OR3x1_ASAP7_75t_R _16246_ (.A(_08580_),
    .B(net58),
    .C(_09119_),
    .Y(_09121_));
 OA211x2_ASAP7_75t_R _16247_ (.A1(_08587_),
    .A2(_09116_),
    .B(_09120_),
    .C(_09121_),
    .Y(_09122_));
 NAND2x1_ASAP7_75t_R _16248_ (.A(_00942_),
    .B(_08610_),
    .Y(_09123_));
 OA21x2_ASAP7_75t_R _16249_ (.A1(_08609_),
    .A2(_09122_),
    .B(_09123_),
    .Y(_01280_));
 OA21x2_ASAP7_75t_R _16250_ (.A1(_01075_),
    .A2(_08664_),
    .B(_01079_),
    .Y(_09124_));
 OA21x2_ASAP7_75t_R _16251_ (.A1(_01078_),
    .A2(_09124_),
    .B(_01082_),
    .Y(_09125_));
 XNOR2x1_ASAP7_75t_R _16252_ (.B(_09125_),
    .Y(_09126_),
    .A(_01081_));
 AND3x1_ASAP7_75t_R _16253_ (.A(_07416_),
    .B(_08703_),
    .C(_07514_),
    .Y(_09127_));
 BUFx6f_ASAP7_75t_R _16254_ (.A(_09127_),
    .Y(\dmem.ce_mem[0] ));
 NAND2x1_ASAP7_75t_R _16255_ (.A(\dmem.inter_dmem3[5] ),
    .B(\dmem.ce_mem[0] ),
    .Y(_09128_));
 NOR2x1_ASAP7_75t_R _16256_ (.A(\dmem.inter_dmem0[5] ),
    .B(_08585_),
    .Y(_09129_));
 OA211x2_ASAP7_75t_R _16257_ (.A1(_08618_),
    .A2(_08621_),
    .B(net38),
    .C(\dmem.inter_dmem2[5] ),
    .Y(_09130_));
 AOI211x1_ASAP7_75t_R _16258_ (.A1(\dmem.inter_dmem1[5] ),
    .A2(_08772_),
    .B(_08628_),
    .C(_09130_),
    .Y(_09131_));
 OA21x2_ASAP7_75t_R _16259_ (.A1(_09129_),
    .A2(_09131_),
    .B(_08580_),
    .Y(_09132_));
 XNOR2x1_ASAP7_75t_R _16260_ (.B(_08674_),
    .Y(_09133_),
    .A(net92));
 OAI22x1_ASAP7_75t_R _16261_ (.A1(net59),
    .A2(_08662_),
    .B1(_09133_),
    .B2(_08583_),
    .Y(_09134_));
 AO221x1_ASAP7_75t_R _16262_ (.A1(_08648_),
    .A2(_09126_),
    .B1(_09128_),
    .B2(_09132_),
    .C(_09134_),
    .Y(_09135_));
 BUFx6f_ASAP7_75t_R _16263_ (.A(_09135_),
    .Y(_09136_));
 BUFx10_ASAP7_75t_R _16264_ (.A(_09136_),
    .Y(_09137_));
 AND2x2_ASAP7_75t_R _16265_ (.A(_00908_),
    .B(_08726_),
    .Y(_09138_));
 AOI21x1_ASAP7_75t_R _16266_ (.A1(_08700_),
    .A2(_09137_),
    .B(_09138_),
    .Y(_01281_));
 OA211x2_ASAP7_75t_R _16267_ (.A1(_08618_),
    .A2(_08621_),
    .B(net38),
    .C(\dmem.inter_dmem2[6] ),
    .Y(_09139_));
 AO21x1_ASAP7_75t_R _16268_ (.A1(\dmem.inter_dmem1[6] ),
    .A2(net47),
    .B(_09139_),
    .Y(_09140_));
 AOI22x1_ASAP7_75t_R _16269_ (.A1(\dmem.inter_dmem3[6] ),
    .A2(\dmem.ce_mem[0] ),
    .B1(_09140_),
    .B2(_08658_),
    .Y(_09141_));
 AOI21x1_ASAP7_75t_R _16270_ (.A1(\dmem.inter_dmem0[6] ),
    .A2(\dmem.ce_mem[3] ),
    .B(_08587_),
    .Y(_09142_));
 OA211x2_ASAP7_75t_R _16271_ (.A1(_07592_),
    .A2(_07915_),
    .B(_07924_),
    .C(_08634_),
    .Y(_09143_));
 OA21x2_ASAP7_75t_R _16272_ (.A1(_01081_),
    .A2(_08637_),
    .B(_01085_),
    .Y(_09144_));
 XNOR2x1_ASAP7_75t_R _16273_ (.B(_09144_),
    .Y(_09145_),
    .A(_01084_));
 XNOR2x1_ASAP7_75t_R _16274_ (.B(_08649_),
    .Y(_09146_),
    .A(_03479_));
 AO32x1_ASAP7_75t_R _16275_ (.A1(_04849_),
    .A2(_08390_),
    .A3(_09145_),
    .B1(_09146_),
    .B2(_08594_),
    .Y(_09147_));
 AOI211x1_ASAP7_75t_R _16276_ (.A1(_09141_),
    .A2(_09142_),
    .B(_09143_),
    .C(_09147_),
    .Y(_09148_));
 NOR2x1_ASAP7_75t_R _16277_ (.A(_00875_),
    .B(_08700_),
    .Y(_09149_));
 AO21x1_ASAP7_75t_R _16278_ (.A1(_08700_),
    .A2(_09148_),
    .B(_09149_),
    .Y(_01282_));
 OR3x1_ASAP7_75t_R _16279_ (.A(_01084_),
    .B(_08666_),
    .C(_08668_),
    .Y(_09150_));
 AND2x2_ASAP7_75t_R _16280_ (.A(_01088_),
    .B(_09150_),
    .Y(_09151_));
 XNOR2x2_ASAP7_75t_R _16281_ (.A(_01087_),
    .B(_09151_),
    .Y(_09152_));
 NOR2x1_ASAP7_75t_R _16282_ (.A(_03479_),
    .B(_08675_),
    .Y(_09153_));
 XNOR2x1_ASAP7_75t_R _16283_ (.B(_09153_),
    .Y(_09154_),
    .A(net94));
 AOI22x1_ASAP7_75t_R _16284_ (.A1(_08648_),
    .A2(_09152_),
    .B1(_09154_),
    .B2(_08594_),
    .Y(_09155_));
 AND2x4_ASAP7_75t_R _16285_ (.A(_07417_),
    .B(_08589_),
    .Y(\dmem.ce_mem[2] ));
 AO21x1_ASAP7_75t_R _16286_ (.A1(\dmem.inter_dmem3[7] ),
    .A2(_08591_),
    .B(_08625_),
    .Y(_09156_));
 AO221x1_ASAP7_75t_R _16287_ (.A1(\dmem.inter_dmem1[7] ),
    .A2(\dmem.ce_mem[2] ),
    .B1(_09111_),
    .B2(_09156_),
    .C(_08712_),
    .Y(_09157_));
 OA211x2_ASAP7_75t_R _16288_ (.A1(net61),
    .A2(_08662_),
    .B(_09155_),
    .C(_09157_),
    .Y(_09158_));
 INVx1_ASAP7_75t_R _16289_ (.A(_00841_),
    .Y(_09159_));
 AND2x2_ASAP7_75t_R _16290_ (.A(_09159_),
    .B(_08726_),
    .Y(_09160_));
 AO21x1_ASAP7_75t_R _16291_ (.A1(_08700_),
    .A2(_09158_),
    .B(_09160_),
    .Y(_01283_));
 AND4x1_ASAP7_75t_R _16292_ (.A(\dmem.inter_dmem2[8] ),
    .B(_07416_),
    .C(net38),
    .D(_08589_),
    .Y(_09161_));
 AND2x2_ASAP7_75t_R _16293_ (.A(\dmem.inter_dmem0[8] ),
    .B(\dmem.ce_mem[3] ),
    .Y(_09162_));
 AND3x1_ASAP7_75t_R _16294_ (.A(\dmem.inter_dmem1[8] ),
    .B(_07339_),
    .C(_07415_),
    .Y(_09163_));
 OA211x2_ASAP7_75t_R _16295_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08591_),
    .C(\dmem.inter_dmem3[8] ),
    .Y(_09164_));
 OA21x2_ASAP7_75t_R _16296_ (.A1(_09163_),
    .A2(_09164_),
    .B(_08585_),
    .Y(_09165_));
 OA33x2_ASAP7_75t_R _16297_ (.A1(_08587_),
    .A2(_05853_),
    .A3(_05946_),
    .B1(_09161_),
    .B2(_09162_),
    .B3(_09165_),
    .Y(_09166_));
 OA21x2_ASAP7_75t_R _16298_ (.A1(_01084_),
    .A2(_09144_),
    .B(_01088_),
    .Y(_09167_));
 OA21x2_ASAP7_75t_R _16299_ (.A1(_01087_),
    .A2(_09167_),
    .B(_01091_),
    .Y(_09168_));
 XOR2x1_ASAP7_75t_R _16300_ (.A(_01090_),
    .Y(_09169_),
    .B(_09168_));
 OR3x1_ASAP7_75t_R _16301_ (.A(_03479_),
    .B(_01086_),
    .C(_08649_),
    .Y(_09170_));
 XNOR2x1_ASAP7_75t_R _16302_ (.B(_09170_),
    .Y(_09171_),
    .A(net95));
 OA222x2_ASAP7_75t_R _16303_ (.A1(net62),
    .A2(_08662_),
    .B1(_09169_),
    .B2(_08394_),
    .C1(_09171_),
    .C2(_08583_),
    .Y(_09172_));
 OA21x2_ASAP7_75t_R _16304_ (.A1(_08748_),
    .A2(_09166_),
    .B(_09172_),
    .Y(_09173_));
 NOR2x1_ASAP7_75t_R _16305_ (.A(_00808_),
    .B(_08700_),
    .Y(_09174_));
 AO21x1_ASAP7_75t_R _16306_ (.A1(_08700_),
    .A2(_09173_),
    .B(_09174_),
    .Y(_01284_));
 OR2x2_ASAP7_75t_R _16307_ (.A(net63),
    .B(_08661_),
    .Y(_09175_));
 XNOR2x2_ASAP7_75t_R _16308_ (.A(_01092_),
    .B(_08676_),
    .Y(_09176_));
 OA21x2_ASAP7_75t_R _16309_ (.A1(_01087_),
    .A2(_09151_),
    .B(_01091_),
    .Y(_09177_));
 OA21x2_ASAP7_75t_R _16310_ (.A1(_01090_),
    .A2(_09177_),
    .B(_01094_),
    .Y(_09178_));
 XNOR2x1_ASAP7_75t_R _16311_ (.B(_09178_),
    .Y(_09179_),
    .A(_01093_));
 AOI22x1_ASAP7_75t_R _16312_ (.A1(_08570_),
    .A2(_09176_),
    .B1(_09179_),
    .B2(_08687_),
    .Y(_09180_));
 OA211x2_ASAP7_75t_R _16313_ (.A1(_08618_),
    .A2(_08621_),
    .B(_08703_),
    .C(\dmem.inter_dmem3[9] ),
    .Y(_09181_));
 AO21x1_ASAP7_75t_R _16314_ (.A1(\dmem.inter_dmem1[9] ),
    .A2(net47),
    .B(_09181_),
    .Y(_09182_));
 AND2x2_ASAP7_75t_R _16315_ (.A(\dmem.inter_dmem0[9] ),
    .B(_08628_),
    .Y(_09183_));
 AO221x1_ASAP7_75t_R _16316_ (.A1(\dmem.inter_dmem2[9] ),
    .A2(\dmem.ce_mem[1] ),
    .B1(_09182_),
    .B2(_08658_),
    .C(_09183_),
    .Y(_09184_));
 AND3x1_ASAP7_75t_R _16317_ (.A(_08612_),
    .B(_09175_),
    .C(_09180_),
    .Y(_09185_));
 AO32x2_ASAP7_75t_R _16318_ (.A1(_08748_),
    .A2(_09175_),
    .A3(_09180_),
    .B1(_09184_),
    .B2(_09185_),
    .Y(_09186_));
 NAND2x1_ASAP7_75t_R _16319_ (.A(_00774_),
    .B(_08610_),
    .Y(_09187_));
 OA21x2_ASAP7_75t_R _16320_ (.A1(_08609_),
    .A2(_09186_),
    .B(_09187_),
    .Y(_01285_));
 INVx1_ASAP7_75t_R _16321_ (.A(_06140_),
    .Y(_09188_));
 AO21x2_ASAP7_75t_R _16322_ (.A1(_03574_),
    .A2(_08600_),
    .B(_09188_),
    .Y(_09189_));
 NOR2x2_ASAP7_75t_R _16323_ (.A(_08598_),
    .B(_09189_),
    .Y(_09190_));
 BUFx12f_ASAP7_75t_R _16324_ (.A(_09190_),
    .Y(_09191_));
 NAND2x2_ASAP7_75t_R _16325_ (.A(_08607_),
    .B(_09191_),
    .Y(_09192_));
 BUFx6f_ASAP7_75t_R _16326_ (.A(_09192_),
    .Y(_09193_));
 BUFx12_ASAP7_75t_R _16327_ (.A(_09192_),
    .Y(_09194_));
 NAND2x1_ASAP7_75t_R _16328_ (.A(_00011_),
    .B(_09194_),
    .Y(_09195_));
 OA21x2_ASAP7_75t_R _16329_ (.A1(_08597_),
    .A2(_09193_),
    .B(_09195_),
    .Y(_01286_));
 BUFx6f_ASAP7_75t_R _16330_ (.A(_08654_),
    .Y(_09196_));
 NAND2x1_ASAP7_75t_R _16331_ (.A(_00743_),
    .B(_09194_),
    .Y(_09197_));
 OA21x2_ASAP7_75t_R _16332_ (.A1(_09196_),
    .A2(_09193_),
    .B(_09197_),
    .Y(_01287_));
 BUFx6f_ASAP7_75t_R _16333_ (.A(_08681_),
    .Y(_09198_));
 NAND2x1_ASAP7_75t_R _16334_ (.A(_00710_),
    .B(_09194_),
    .Y(_09199_));
 OA21x2_ASAP7_75t_R _16335_ (.A1(_09198_),
    .A2(_09193_),
    .B(_09199_),
    .Y(_01288_));
 BUFx4f_ASAP7_75t_R _16336_ (.A(_08697_),
    .Y(_09200_));
 NAND2x1_ASAP7_75t_R _16337_ (.A(_00677_),
    .B(_09194_),
    .Y(_09201_));
 OA21x2_ASAP7_75t_R _16338_ (.A1(_09200_),
    .A2(_09193_),
    .B(_09201_),
    .Y(_01289_));
 AND2x6_ASAP7_75t_R _16339_ (.A(_08606_),
    .B(_09191_),
    .Y(_09202_));
 BUFx6f_ASAP7_75t_R _16340_ (.A(_09202_),
    .Y(_09203_));
 BUFx10_ASAP7_75t_R _16341_ (.A(_09192_),
    .Y(_09204_));
 AND2x2_ASAP7_75t_R _16342_ (.A(_00644_),
    .B(_09204_),
    .Y(_09205_));
 AOI21x1_ASAP7_75t_R _16343_ (.A1(_08725_),
    .A2(_09203_),
    .B(_09205_),
    .Y(_01290_));
 BUFx4f_ASAP7_75t_R _16344_ (.A(_08744_),
    .Y(_09206_));
 NAND2x1_ASAP7_75t_R _16345_ (.A(_00611_),
    .B(_09194_),
    .Y(_09207_));
 OA21x2_ASAP7_75t_R _16346_ (.A1(_09206_),
    .A2(_09193_),
    .B(_09207_),
    .Y(_01291_));
 BUFx4f_ASAP7_75t_R _16347_ (.A(_08607_),
    .Y(_09208_));
 AO21x1_ASAP7_75t_R _16348_ (.A1(_09208_),
    .A2(_09191_),
    .B(_00577_),
    .Y(_09209_));
 OAI21x1_ASAP7_75t_R _16349_ (.A1(_08766_),
    .A2(_09193_),
    .B(_09209_),
    .Y(_01292_));
 BUFx6f_ASAP7_75t_R _16350_ (.A(_08786_),
    .Y(_09210_));
 BUFx6f_ASAP7_75t_R _16351_ (.A(_08794_),
    .Y(_09211_));
 AND3x1_ASAP7_75t_R _16352_ (.A(_09210_),
    .B(_09211_),
    .C(_09203_),
    .Y(_09212_));
 BUFx12f_ASAP7_75t_R _16353_ (.A(_09192_),
    .Y(_09213_));
 INVx1_ASAP7_75t_R _16354_ (.A(_00544_),
    .Y(_09214_));
 AO32x1_ASAP7_75t_R _16355_ (.A1(_08783_),
    .A2(_08785_),
    .A3(_09212_),
    .B1(_09213_),
    .B2(_09214_),
    .Y(_01293_));
 BUFx4f_ASAP7_75t_R _16356_ (.A(_08821_),
    .Y(_09215_));
 BUFx4f_ASAP7_75t_R _16357_ (.A(_09202_),
    .Y(_09216_));
 AND2x2_ASAP7_75t_R _16358_ (.A(_09215_),
    .B(_09216_),
    .Y(_09217_));
 INVx1_ASAP7_75t_R _16359_ (.A(_00511_),
    .Y(_09218_));
 AO32x1_ASAP7_75t_R _16360_ (.A1(_09019_),
    .A2(_08805_),
    .A3(_09217_),
    .B1(_09213_),
    .B2(_09218_),
    .Y(_01294_));
 BUFx6f_ASAP7_75t_R _16361_ (.A(_08834_),
    .Y(_09219_));
 BUFx4f_ASAP7_75t_R _16362_ (.A(_08841_),
    .Y(_09220_));
 AND3x1_ASAP7_75t_R _16363_ (.A(_09219_),
    .B(_09220_),
    .C(_09216_),
    .Y(_09221_));
 INVx1_ASAP7_75t_R _16364_ (.A(_00478_),
    .Y(_09222_));
 AO32x1_ASAP7_75t_R _16365_ (.A1(_09019_),
    .A2(_08830_),
    .A3(_09221_),
    .B1(_09213_),
    .B2(_09222_),
    .Y(_01295_));
 BUFx4f_ASAP7_75t_R _16366_ (.A(_08851_),
    .Y(_09223_));
 BUFx4f_ASAP7_75t_R _16367_ (.A(_08860_),
    .Y(_09224_));
 AND3x1_ASAP7_75t_R _16368_ (.A(_09223_),
    .B(_09224_),
    .C(_09216_),
    .Y(_09225_));
 INVx1_ASAP7_75t_R _16369_ (.A(_00445_),
    .Y(_09226_));
 AO32x1_ASAP7_75t_R _16370_ (.A1(_09019_),
    .A2(_08850_),
    .A3(_09225_),
    .B1(_09213_),
    .B2(_09226_),
    .Y(_01296_));
 BUFx4f_ASAP7_75t_R _16371_ (.A(_08870_),
    .Y(_09227_));
 NAND2x1_ASAP7_75t_R _16372_ (.A(_01042_),
    .B(_09194_),
    .Y(_09228_));
 OA21x2_ASAP7_75t_R _16373_ (.A1(_09227_),
    .A2(_09193_),
    .B(_09228_),
    .Y(_01297_));
 BUFx4f_ASAP7_75t_R _16374_ (.A(_08892_),
    .Y(_09229_));
 AND2x2_ASAP7_75t_R _16375_ (.A(_09229_),
    .B(_09216_),
    .Y(_09230_));
 INVx1_ASAP7_75t_R _16376_ (.A(_00412_),
    .Y(_09231_));
 AO32x1_ASAP7_75t_R _16377_ (.A1(_09019_),
    .A2(_08879_),
    .A3(_09230_),
    .B1(_09213_),
    .B2(_09231_),
    .Y(_01298_));
 BUFx4f_ASAP7_75t_R _16378_ (.A(_08902_),
    .Y(_09232_));
 BUFx4f_ASAP7_75t_R _16379_ (.A(_08910_),
    .Y(_09233_));
 AND3x1_ASAP7_75t_R _16380_ (.A(_09232_),
    .B(_09233_),
    .C(_09216_),
    .Y(_09234_));
 INVx1_ASAP7_75t_R _16381_ (.A(_00379_),
    .Y(_09235_));
 AO32x1_ASAP7_75t_R _16382_ (.A1(_09019_),
    .A2(_08901_),
    .A3(_09234_),
    .B1(_09213_),
    .B2(_09235_),
    .Y(_01299_));
 BUFx4f_ASAP7_75t_R _16383_ (.A(_08929_),
    .Y(_09236_));
 AND2x2_ASAP7_75t_R _16384_ (.A(_09236_),
    .B(_09216_),
    .Y(_09237_));
 INVx1_ASAP7_75t_R _16385_ (.A(_00346_),
    .Y(_09238_));
 AO32x1_ASAP7_75t_R _16386_ (.A1(_09019_),
    .A2(_08918_),
    .A3(_09237_),
    .B1(_09213_),
    .B2(_09238_),
    .Y(_01300_));
 BUFx4f_ASAP7_75t_R _16387_ (.A(_08798_),
    .Y(_09239_));
 BUFx4f_ASAP7_75t_R _16388_ (.A(_08943_),
    .Y(_09240_));
 AND2x2_ASAP7_75t_R _16389_ (.A(_09240_),
    .B(_09216_),
    .Y(_09241_));
 INVx1_ASAP7_75t_R _16390_ (.A(_00312_),
    .Y(_09242_));
 AO32x1_ASAP7_75t_R _16391_ (.A1(_09239_),
    .A2(_08937_),
    .A3(_09241_),
    .B1(_09213_),
    .B2(_09242_),
    .Y(_01301_));
 BUFx4f_ASAP7_75t_R _16392_ (.A(_08962_),
    .Y(_09243_));
 AND2x2_ASAP7_75t_R _16393_ (.A(_09243_),
    .B(_09216_),
    .Y(_09244_));
 INVx1_ASAP7_75t_R _16394_ (.A(_00279_),
    .Y(_09245_));
 AO32x1_ASAP7_75t_R _16395_ (.A1(_09239_),
    .A2(_08951_),
    .A3(_09244_),
    .B1(_09204_),
    .B2(_09245_),
    .Y(_01302_));
 BUFx4f_ASAP7_75t_R _16396_ (.A(_08979_),
    .Y(_09246_));
 AND2x2_ASAP7_75t_R _16397_ (.A(_09246_),
    .B(_09202_),
    .Y(_09247_));
 INVx1_ASAP7_75t_R _16398_ (.A(_00246_),
    .Y(_09248_));
 AO32x1_ASAP7_75t_R _16399_ (.A1(_09239_),
    .A2(_08970_),
    .A3(_09247_),
    .B1(_09204_),
    .B2(_09248_),
    .Y(_01303_));
 NOR2x1_ASAP7_75t_R _16400_ (.A(_08997_),
    .B(_09204_),
    .Y(_09249_));
 INVx1_ASAP7_75t_R _16401_ (.A(_00213_),
    .Y(_09250_));
 AO32x1_ASAP7_75t_R _16402_ (.A1(_09239_),
    .A2(_08987_),
    .A3(_09249_),
    .B1(_09204_),
    .B2(_09250_),
    .Y(_01304_));
 INVx1_ASAP7_75t_R _16403_ (.A(_00179_),
    .Y(_09251_));
 BUFx4f_ASAP7_75t_R _16404_ (.A(_09017_),
    .Y(_09252_));
 AND2x2_ASAP7_75t_R _16405_ (.A(_09252_),
    .B(_09203_),
    .Y(_09253_));
 AO22x1_ASAP7_75t_R _16406_ (.A1(_09251_),
    .A2(_09194_),
    .B1(_09253_),
    .B2(_09006_),
    .Y(_01305_));
 BUFx4f_ASAP7_75t_R _16407_ (.A(_09030_),
    .Y(_09254_));
 BUFx4f_ASAP7_75t_R _16408_ (.A(_09031_),
    .Y(_09255_));
 BUFx4f_ASAP7_75t_R _16409_ (.A(_09035_),
    .Y(_09256_));
 AND4x1_ASAP7_75t_R _16410_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09202_),
    .Y(_09257_));
 INVx1_ASAP7_75t_R _16411_ (.A(_00146_),
    .Y(_09258_));
 AO32x1_ASAP7_75t_R _16412_ (.A1(_09239_),
    .A2(_09025_),
    .A3(_09257_),
    .B1(_09204_),
    .B2(_09258_),
    .Y(_01306_));
 BUFx4f_ASAP7_75t_R _16413_ (.A(_09048_),
    .Y(_09259_));
 BUFx4f_ASAP7_75t_R _16414_ (.A(_09051_),
    .Y(_09260_));
 AND3x1_ASAP7_75t_R _16415_ (.A(_09259_),
    .B(_09260_),
    .C(_09216_),
    .Y(_09261_));
 INVx1_ASAP7_75t_R _16416_ (.A(_00112_),
    .Y(_09262_));
 AO32x1_ASAP7_75t_R _16417_ (.A1(_09239_),
    .A2(_09043_),
    .A3(_09261_),
    .B1(_09204_),
    .B2(_09262_),
    .Y(_01307_));
 BUFx4f_ASAP7_75t_R _16418_ (.A(_09063_),
    .Y(_09263_));
 NAND2x1_ASAP7_75t_R _16419_ (.A(_01009_),
    .B(_09194_),
    .Y(_09264_));
 OA21x2_ASAP7_75t_R _16420_ (.A1(_09263_),
    .A2(_09193_),
    .B(_09264_),
    .Y(_01308_));
 BUFx4f_ASAP7_75t_R _16421_ (.A(_09074_),
    .Y(_09265_));
 BUFx4f_ASAP7_75t_R _16422_ (.A(_09077_),
    .Y(_09266_));
 BUFx4f_ASAP7_75t_R _16423_ (.A(_09078_),
    .Y(_09267_));
 AND4x1_ASAP7_75t_R _16424_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09202_),
    .Y(_09268_));
 INVx1_ASAP7_75t_R _16425_ (.A(_00078_),
    .Y(_09269_));
 AO32x1_ASAP7_75t_R _16426_ (.A1(_09239_),
    .A2(_09070_),
    .A3(_09268_),
    .B1(_09204_),
    .B2(_09269_),
    .Y(_01309_));
 BUFx4f_ASAP7_75t_R _16427_ (.A(_09094_),
    .Y(_09270_));
 BUFx4f_ASAP7_75t_R _16428_ (.A(_09097_),
    .Y(_09271_));
 AND3x1_ASAP7_75t_R _16429_ (.A(_09270_),
    .B(_09271_),
    .C(_09216_),
    .Y(_09272_));
 INVx1_ASAP7_75t_R _16430_ (.A(_00046_),
    .Y(_09273_));
 AO32x1_ASAP7_75t_R _16431_ (.A1(_09239_),
    .A2(_09086_),
    .A3(_09272_),
    .B1(_09204_),
    .B2(_09273_),
    .Y(_01310_));
 BUFx3_ASAP7_75t_R _16432_ (.A(_09109_),
    .Y(_09274_));
 NAND2x1_ASAP7_75t_R _16433_ (.A(_00976_),
    .B(_09194_),
    .Y(_09275_));
 OA21x2_ASAP7_75t_R _16434_ (.A1(_09274_),
    .A2(_09193_),
    .B(_09275_),
    .Y(_01311_));
 BUFx6f_ASAP7_75t_R _16435_ (.A(_09122_),
    .Y(_09276_));
 NAND2x1_ASAP7_75t_R _16436_ (.A(_00943_),
    .B(_09213_),
    .Y(_09277_));
 OA21x2_ASAP7_75t_R _16437_ (.A1(_09276_),
    .A2(_09193_),
    .B(_09277_),
    .Y(_01312_));
 AND2x2_ASAP7_75t_R _16438_ (.A(_00909_),
    .B(_09204_),
    .Y(_09278_));
 AOI21x1_ASAP7_75t_R _16439_ (.A1(_09137_),
    .A2(_09203_),
    .B(_09278_),
    .Y(_01313_));
 BUFx4f_ASAP7_75t_R _16440_ (.A(_09148_),
    .Y(_09279_));
 NOR2x1_ASAP7_75t_R _16441_ (.A(_00876_),
    .B(_09203_),
    .Y(_09280_));
 AO21x1_ASAP7_75t_R _16442_ (.A1(_09279_),
    .A2(_09203_),
    .B(_09280_),
    .Y(_01314_));
 BUFx4f_ASAP7_75t_R _16443_ (.A(_09158_),
    .Y(_09281_));
 NOR2x1_ASAP7_75t_R _16444_ (.A(_00842_),
    .B(_09203_),
    .Y(_09282_));
 AO21x1_ASAP7_75t_R _16445_ (.A1(_09281_),
    .A2(_09203_),
    .B(_09282_),
    .Y(_01315_));
 BUFx4f_ASAP7_75t_R _16446_ (.A(_09173_),
    .Y(_09283_));
 NOR2x1_ASAP7_75t_R _16447_ (.A(_00809_),
    .B(_09203_),
    .Y(_09284_));
 AO21x1_ASAP7_75t_R _16448_ (.A1(_09283_),
    .A2(_09203_),
    .B(_09284_),
    .Y(_01316_));
 BUFx6f_ASAP7_75t_R _16449_ (.A(_09186_),
    .Y(_09285_));
 NAND2x1_ASAP7_75t_R _16450_ (.A(_00775_),
    .B(_09213_),
    .Y(_09286_));
 OA21x2_ASAP7_75t_R _16451_ (.A1(_09285_),
    .A2(_09194_),
    .B(_09286_),
    .Y(_01317_));
 OA21x2_ASAP7_75t_R _16452_ (.A1(net3),
    .A2(net2),
    .B(_03382_),
    .Y(_09287_));
 NOR2x2_ASAP7_75t_R _16453_ (.A(_08603_),
    .B(_09287_),
    .Y(_09288_));
 OR3x4_ASAP7_75t_R _16454_ (.A(_07131_),
    .B(_08601_),
    .C(_09288_),
    .Y(_09289_));
 AO21x1_ASAP7_75t_R _16455_ (.A1(_03566_),
    .A2(_07020_),
    .B(_08605_),
    .Y(_09290_));
 BUFx6f_ASAP7_75t_R _16456_ (.A(_09290_),
    .Y(_09291_));
 OR2x6_ASAP7_75t_R _16457_ (.A(_09289_),
    .B(_09291_),
    .Y(_09292_));
 BUFx6f_ASAP7_75t_R _16458_ (.A(_09292_),
    .Y(_09293_));
 BUFx10_ASAP7_75t_R _16459_ (.A(_09292_),
    .Y(_09294_));
 NAND2x1_ASAP7_75t_R _16460_ (.A(_00012_),
    .B(_09294_),
    .Y(_09295_));
 OA21x2_ASAP7_75t_R _16461_ (.A1(_08597_),
    .A2(_09293_),
    .B(_09295_),
    .Y(_01318_));
 NAND2x1_ASAP7_75t_R _16462_ (.A(_00744_),
    .B(_09294_),
    .Y(_09296_));
 OA21x2_ASAP7_75t_R _16463_ (.A1(_09196_),
    .A2(_09293_),
    .B(_09296_),
    .Y(_01319_));
 NAND2x1_ASAP7_75t_R _16464_ (.A(_00711_),
    .B(_09294_),
    .Y(_09297_));
 OA21x2_ASAP7_75t_R _16465_ (.A1(_09198_),
    .A2(_09293_),
    .B(_09297_),
    .Y(_01320_));
 NAND2x1_ASAP7_75t_R _16466_ (.A(_00678_),
    .B(_09294_),
    .Y(_09298_));
 OA21x2_ASAP7_75t_R _16467_ (.A1(_09200_),
    .A2(_09293_),
    .B(_09298_),
    .Y(_01321_));
 NOR2x2_ASAP7_75t_R _16468_ (.A(_09289_),
    .B(_09291_),
    .Y(_09299_));
 BUFx6f_ASAP7_75t_R _16469_ (.A(_09299_),
    .Y(_09300_));
 BUFx10_ASAP7_75t_R _16470_ (.A(_09292_),
    .Y(_09301_));
 AND2x2_ASAP7_75t_R _16471_ (.A(_00645_),
    .B(_09301_),
    .Y(_09302_));
 AOI21x1_ASAP7_75t_R _16472_ (.A1(_08725_),
    .A2(_09300_),
    .B(_09302_),
    .Y(_01322_));
 NAND2x1_ASAP7_75t_R _16473_ (.A(_00612_),
    .B(_09294_),
    .Y(_09303_));
 OA21x2_ASAP7_75t_R _16474_ (.A1(_09206_),
    .A2(_09293_),
    .B(_09303_),
    .Y(_01323_));
 OR2x2_ASAP7_75t_R _16475_ (.A(_00578_),
    .B(_09300_),
    .Y(_09304_));
 OAI21x1_ASAP7_75t_R _16476_ (.A1(_08766_),
    .A2(_09293_),
    .B(_09304_),
    .Y(_01324_));
 BUFx3_ASAP7_75t_R _16477_ (.A(_09299_),
    .Y(_09305_));
 AND3x4_ASAP7_75t_R _16478_ (.A(_09210_),
    .B(_09211_),
    .C(_09305_),
    .Y(_09306_));
 BUFx10_ASAP7_75t_R _16479_ (.A(_09292_),
    .Y(_09307_));
 INVx1_ASAP7_75t_R _16480_ (.A(_00545_),
    .Y(_09308_));
 AO32x1_ASAP7_75t_R _16481_ (.A1(_08783_),
    .A2(_08785_),
    .A3(_09306_),
    .B1(_09307_),
    .B2(_09308_),
    .Y(_01325_));
 AND2x2_ASAP7_75t_R _16482_ (.A(_09215_),
    .B(_09305_),
    .Y(_09309_));
 INVx1_ASAP7_75t_R _16483_ (.A(_00512_),
    .Y(_09310_));
 AO32x1_ASAP7_75t_R _16484_ (.A1(_09239_),
    .A2(_08805_),
    .A3(_09309_),
    .B1(_09307_),
    .B2(_09310_),
    .Y(_01326_));
 AND3x1_ASAP7_75t_R _16485_ (.A(_09219_),
    .B(_09220_),
    .C(_09305_),
    .Y(_09311_));
 INVx1_ASAP7_75t_R _16486_ (.A(_00479_),
    .Y(_09312_));
 AO32x1_ASAP7_75t_R _16487_ (.A1(_09239_),
    .A2(_08830_),
    .A3(_09311_),
    .B1(_09307_),
    .B2(_09312_),
    .Y(_01327_));
 BUFx3_ASAP7_75t_R _16488_ (.A(_08798_),
    .Y(_09313_));
 AND3x1_ASAP7_75t_R _16489_ (.A(_09223_),
    .B(_09224_),
    .C(_09305_),
    .Y(_09314_));
 INVx1_ASAP7_75t_R _16490_ (.A(_00446_),
    .Y(_09315_));
 AO32x1_ASAP7_75t_R _16491_ (.A1(_09313_),
    .A2(_08850_),
    .A3(_09314_),
    .B1(_09307_),
    .B2(_09315_),
    .Y(_01328_));
 NAND2x1_ASAP7_75t_R _16492_ (.A(_01043_),
    .B(_09294_),
    .Y(_09316_));
 OA21x2_ASAP7_75t_R _16493_ (.A1(_09227_),
    .A2(_09293_),
    .B(_09316_),
    .Y(_01329_));
 AND2x2_ASAP7_75t_R _16494_ (.A(_09229_),
    .B(_09305_),
    .Y(_09317_));
 INVx1_ASAP7_75t_R _16495_ (.A(_00413_),
    .Y(_09318_));
 AO32x1_ASAP7_75t_R _16496_ (.A1(_09313_),
    .A2(_08879_),
    .A3(_09317_),
    .B1(_09307_),
    .B2(_09318_),
    .Y(_01330_));
 AND3x1_ASAP7_75t_R _16497_ (.A(_09232_),
    .B(_09233_),
    .C(_09305_),
    .Y(_09319_));
 INVx1_ASAP7_75t_R _16498_ (.A(_00380_),
    .Y(_09320_));
 AO32x1_ASAP7_75t_R _16499_ (.A1(_09313_),
    .A2(_08901_),
    .A3(_09319_),
    .B1(_09307_),
    .B2(_09320_),
    .Y(_01331_));
 AND2x2_ASAP7_75t_R _16500_ (.A(_09236_),
    .B(_09305_),
    .Y(_09321_));
 INVx1_ASAP7_75t_R _16501_ (.A(_00347_),
    .Y(_09322_));
 AO32x1_ASAP7_75t_R _16502_ (.A1(_09313_),
    .A2(_08918_),
    .A3(_09321_),
    .B1(_09307_),
    .B2(_09322_),
    .Y(_01332_));
 AND2x2_ASAP7_75t_R _16503_ (.A(_09240_),
    .B(_09305_),
    .Y(_09323_));
 INVx1_ASAP7_75t_R _16504_ (.A(_00313_),
    .Y(_09324_));
 AO32x1_ASAP7_75t_R _16505_ (.A1(_09313_),
    .A2(_08937_),
    .A3(_09323_),
    .B1(_09307_),
    .B2(_09324_),
    .Y(_01333_));
 AND2x2_ASAP7_75t_R _16506_ (.A(_09243_),
    .B(_09299_),
    .Y(_09325_));
 INVx1_ASAP7_75t_R _16507_ (.A(_00280_),
    .Y(_09326_));
 AO32x1_ASAP7_75t_R _16508_ (.A1(_09313_),
    .A2(_08951_),
    .A3(_09325_),
    .B1(_09301_),
    .B2(_09326_),
    .Y(_01334_));
 AND2x2_ASAP7_75t_R _16509_ (.A(_09246_),
    .B(_09299_),
    .Y(_09327_));
 INVx1_ASAP7_75t_R _16510_ (.A(_00247_),
    .Y(_09328_));
 AO32x1_ASAP7_75t_R _16511_ (.A1(_09313_),
    .A2(_08970_),
    .A3(_09327_),
    .B1(_09301_),
    .B2(_09328_),
    .Y(_01335_));
 NOR2x1_ASAP7_75t_R _16512_ (.A(_08997_),
    .B(_09301_),
    .Y(_09329_));
 INVx1_ASAP7_75t_R _16513_ (.A(_00214_),
    .Y(_09330_));
 AO32x1_ASAP7_75t_R _16514_ (.A1(_09313_),
    .A2(_08987_),
    .A3(_09329_),
    .B1(_09301_),
    .B2(_09330_),
    .Y(_01336_));
 INVx1_ASAP7_75t_R _16515_ (.A(_00180_),
    .Y(_09331_));
 AND2x2_ASAP7_75t_R _16516_ (.A(_09252_),
    .B(_09300_),
    .Y(_09332_));
 AO22x1_ASAP7_75t_R _16517_ (.A1(_09331_),
    .A2(_09294_),
    .B1(_09332_),
    .B2(_09006_),
    .Y(_01337_));
 AND4x1_ASAP7_75t_R _16518_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09299_),
    .Y(_09333_));
 AO32x1_ASAP7_75t_R _16519_ (.A1(_09313_),
    .A2(_09025_),
    .A3(_09333_),
    .B1(_09301_),
    .B2(_04410_),
    .Y(_01338_));
 AND3x1_ASAP7_75t_R _16520_ (.A(_09259_),
    .B(_09260_),
    .C(_09305_),
    .Y(_09334_));
 INVx1_ASAP7_75t_R _16521_ (.A(_00113_),
    .Y(_09335_));
 AO32x1_ASAP7_75t_R _16522_ (.A1(_09313_),
    .A2(_09043_),
    .A3(_09334_),
    .B1(_09301_),
    .B2(_09335_),
    .Y(_01339_));
 NAND2x1_ASAP7_75t_R _16523_ (.A(_01010_),
    .B(_09294_),
    .Y(_09336_));
 OA21x2_ASAP7_75t_R _16524_ (.A1(_09263_),
    .A2(_09293_),
    .B(_09336_),
    .Y(_01340_));
 BUFx4f_ASAP7_75t_R _16525_ (.A(_08798_),
    .Y(_09337_));
 AND4x1_ASAP7_75t_R _16526_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09299_),
    .Y(_09338_));
 INVx1_ASAP7_75t_R _16527_ (.A(_00079_),
    .Y(_09339_));
 AO32x1_ASAP7_75t_R _16528_ (.A1(_09337_),
    .A2(_09070_),
    .A3(_09338_),
    .B1(_09301_),
    .B2(_09339_),
    .Y(_01341_));
 AND3x1_ASAP7_75t_R _16529_ (.A(_09270_),
    .B(_09271_),
    .C(_09305_),
    .Y(_09340_));
 INVx1_ASAP7_75t_R _16530_ (.A(_00047_),
    .Y(_09341_));
 AO32x1_ASAP7_75t_R _16531_ (.A1(_09337_),
    .A2(_09086_),
    .A3(_09340_),
    .B1(_09301_),
    .B2(_09341_),
    .Y(_01342_));
 NAND2x1_ASAP7_75t_R _16532_ (.A(_00977_),
    .B(_09294_),
    .Y(_09342_));
 OA21x2_ASAP7_75t_R _16533_ (.A1(_09274_),
    .A2(_09293_),
    .B(_09342_),
    .Y(_01343_));
 NAND2x1_ASAP7_75t_R _16534_ (.A(_00944_),
    .B(_09307_),
    .Y(_09343_));
 OA21x2_ASAP7_75t_R _16535_ (.A1(_09276_),
    .A2(_09293_),
    .B(_09343_),
    .Y(_01344_));
 AND2x2_ASAP7_75t_R _16536_ (.A(_00910_),
    .B(_09301_),
    .Y(_09344_));
 AOI21x1_ASAP7_75t_R _16537_ (.A1(_09137_),
    .A2(_09300_),
    .B(_09344_),
    .Y(_01345_));
 NOR2x1_ASAP7_75t_R _16538_ (.A(_00877_),
    .B(_09300_),
    .Y(_09345_));
 AO21x1_ASAP7_75t_R _16539_ (.A1(_09279_),
    .A2(_09300_),
    .B(_09345_),
    .Y(_01346_));
 NOR2x1_ASAP7_75t_R _16540_ (.A(_00843_),
    .B(_09300_),
    .Y(_09346_));
 AO21x1_ASAP7_75t_R _16541_ (.A1(_09281_),
    .A2(_09300_),
    .B(_09346_),
    .Y(_01347_));
 NOR2x1_ASAP7_75t_R _16542_ (.A(_00810_),
    .B(_09300_),
    .Y(_09347_));
 AO21x1_ASAP7_75t_R _16543_ (.A1(_09283_),
    .A2(_09300_),
    .B(_09347_),
    .Y(_01348_));
 NAND2x1_ASAP7_75t_R _16544_ (.A(_00776_),
    .B(_09307_),
    .Y(_09348_));
 OA21x2_ASAP7_75t_R _16545_ (.A1(_09285_),
    .A2(_09294_),
    .B(_09348_),
    .Y(_01349_));
 BUFx4f_ASAP7_75t_R _16546_ (.A(_09189_),
    .Y(_09349_));
 OR3x4_ASAP7_75t_R _16547_ (.A(_07131_),
    .B(_09349_),
    .C(_09291_),
    .Y(_09350_));
 BUFx6f_ASAP7_75t_R _16548_ (.A(_09350_),
    .Y(_09351_));
 BUFx10_ASAP7_75t_R _16549_ (.A(_09350_),
    .Y(_09352_));
 NAND2x1_ASAP7_75t_R _16550_ (.A(_00013_),
    .B(_09352_),
    .Y(_09353_));
 OA21x2_ASAP7_75t_R _16551_ (.A1(_08597_),
    .A2(_09351_),
    .B(_09353_),
    .Y(_01350_));
 NAND2x1_ASAP7_75t_R _16552_ (.A(_00745_),
    .B(_09352_),
    .Y(_09354_));
 OA21x2_ASAP7_75t_R _16553_ (.A1(_09196_),
    .A2(_09351_),
    .B(_09354_),
    .Y(_01351_));
 NAND2x1_ASAP7_75t_R _16554_ (.A(_00712_),
    .B(_09352_),
    .Y(_09355_));
 OA21x2_ASAP7_75t_R _16555_ (.A1(_09198_),
    .A2(_09351_),
    .B(_09355_),
    .Y(_01352_));
 NAND2x1_ASAP7_75t_R _16556_ (.A(_00679_),
    .B(_09352_),
    .Y(_09356_));
 OA21x2_ASAP7_75t_R _16557_ (.A1(_09200_),
    .A2(_09351_),
    .B(_09356_),
    .Y(_01353_));
 OR2x6_ASAP7_75t_R _16558_ (.A(_07131_),
    .B(_09349_),
    .Y(_09357_));
 NOR2x2_ASAP7_75t_R _16559_ (.A(_09291_),
    .B(_09357_),
    .Y(_09358_));
 BUFx6f_ASAP7_75t_R _16560_ (.A(_09358_),
    .Y(_09359_));
 BUFx12_ASAP7_75t_R _16561_ (.A(_09350_),
    .Y(_09360_));
 AND2x2_ASAP7_75t_R _16562_ (.A(_00646_),
    .B(_09360_),
    .Y(_09361_));
 AOI21x1_ASAP7_75t_R _16563_ (.A1(_08725_),
    .A2(_09359_),
    .B(_09361_),
    .Y(_01354_));
 NAND2x1_ASAP7_75t_R _16564_ (.A(_00613_),
    .B(_09352_),
    .Y(_09362_));
 OA21x2_ASAP7_75t_R _16565_ (.A1(_09206_),
    .A2(_09351_),
    .B(_09362_),
    .Y(_01355_));
 OR2x2_ASAP7_75t_R _16566_ (.A(_00579_),
    .B(_09359_),
    .Y(_09363_));
 OAI21x1_ASAP7_75t_R _16567_ (.A1(_08766_),
    .A2(_09351_),
    .B(_09363_),
    .Y(_01356_));
 BUFx4f_ASAP7_75t_R _16568_ (.A(_09358_),
    .Y(_09364_));
 AND3x1_ASAP7_75t_R _16569_ (.A(_09210_),
    .B(_09211_),
    .C(_09364_),
    .Y(_09365_));
 BUFx10_ASAP7_75t_R _16570_ (.A(_09350_),
    .Y(_09366_));
 INVx1_ASAP7_75t_R _16571_ (.A(_00546_),
    .Y(_09367_));
 AO32x1_ASAP7_75t_R _16572_ (.A1(_08783_),
    .A2(_08785_),
    .A3(_09365_),
    .B1(_09366_),
    .B2(_09367_),
    .Y(_01357_));
 AND2x2_ASAP7_75t_R _16573_ (.A(_09215_),
    .B(_09364_),
    .Y(_09368_));
 INVx1_ASAP7_75t_R _16574_ (.A(_00513_),
    .Y(_09369_));
 AO32x1_ASAP7_75t_R _16575_ (.A1(_09337_),
    .A2(_08805_),
    .A3(_09368_),
    .B1(_09366_),
    .B2(_09369_),
    .Y(_01358_));
 AND3x1_ASAP7_75t_R _16576_ (.A(_09219_),
    .B(_09220_),
    .C(_09364_),
    .Y(_09370_));
 INVx1_ASAP7_75t_R _16577_ (.A(_00480_),
    .Y(_09371_));
 AO32x1_ASAP7_75t_R _16578_ (.A1(_09337_),
    .A2(_08830_),
    .A3(_09370_),
    .B1(_09366_),
    .B2(_09371_),
    .Y(_01359_));
 AND3x1_ASAP7_75t_R _16579_ (.A(_09223_),
    .B(_09224_),
    .C(_09364_),
    .Y(_09372_));
 INVx1_ASAP7_75t_R _16580_ (.A(_00447_),
    .Y(_09373_));
 AO32x1_ASAP7_75t_R _16581_ (.A1(_09337_),
    .A2(_08850_),
    .A3(_09372_),
    .B1(_09366_),
    .B2(_09373_),
    .Y(_01360_));
 NAND2x1_ASAP7_75t_R _16582_ (.A(_01044_),
    .B(_09352_),
    .Y(_09374_));
 OA21x2_ASAP7_75t_R _16583_ (.A1(_09227_),
    .A2(_09351_),
    .B(_09374_),
    .Y(_01361_));
 AND2x2_ASAP7_75t_R _16584_ (.A(_09229_),
    .B(_09364_),
    .Y(_09375_));
 INVx1_ASAP7_75t_R _16585_ (.A(_00414_),
    .Y(_09376_));
 AO32x1_ASAP7_75t_R _16586_ (.A1(_09337_),
    .A2(_08879_),
    .A3(_09375_),
    .B1(_09366_),
    .B2(_09376_),
    .Y(_01362_));
 AND3x1_ASAP7_75t_R _16587_ (.A(_09232_),
    .B(_09233_),
    .C(_09364_),
    .Y(_09377_));
 INVx1_ASAP7_75t_R _16588_ (.A(_00381_),
    .Y(_09378_));
 AO32x1_ASAP7_75t_R _16589_ (.A1(_09337_),
    .A2(_08901_),
    .A3(_09377_),
    .B1(_09366_),
    .B2(_09378_),
    .Y(_01363_));
 AND2x2_ASAP7_75t_R _16590_ (.A(_09236_),
    .B(_09364_),
    .Y(_09379_));
 INVx1_ASAP7_75t_R _16591_ (.A(_00348_),
    .Y(_09380_));
 AO32x1_ASAP7_75t_R _16592_ (.A1(_09337_),
    .A2(_08918_),
    .A3(_09379_),
    .B1(_09366_),
    .B2(_09380_),
    .Y(_01364_));
 AND2x2_ASAP7_75t_R _16593_ (.A(_09240_),
    .B(_09364_),
    .Y(_09381_));
 INVx1_ASAP7_75t_R _16594_ (.A(_00314_),
    .Y(_09382_));
 AO32x1_ASAP7_75t_R _16595_ (.A1(_09337_),
    .A2(_08937_),
    .A3(_09381_),
    .B1(_09366_),
    .B2(_09382_),
    .Y(_01365_));
 AND2x2_ASAP7_75t_R _16596_ (.A(_09243_),
    .B(_09358_),
    .Y(_09383_));
 INVx1_ASAP7_75t_R _16597_ (.A(_00281_),
    .Y(_09384_));
 AO32x1_ASAP7_75t_R _16598_ (.A1(_09337_),
    .A2(_08951_),
    .A3(_09383_),
    .B1(_09360_),
    .B2(_09384_),
    .Y(_01366_));
 BUFx6f_ASAP7_75t_R _16599_ (.A(_08784_),
    .Y(_09385_));
 BUFx4f_ASAP7_75t_R _16600_ (.A(_09385_),
    .Y(_09386_));
 AND2x2_ASAP7_75t_R _16601_ (.A(_09246_),
    .B(_09358_),
    .Y(_09387_));
 INVx1_ASAP7_75t_R _16602_ (.A(_00248_),
    .Y(_09388_));
 AO32x1_ASAP7_75t_R _16603_ (.A1(_09386_),
    .A2(_08970_),
    .A3(_09387_),
    .B1(_09360_),
    .B2(_09388_),
    .Y(_01367_));
 NOR2x1_ASAP7_75t_R _16604_ (.A(_08997_),
    .B(_09360_),
    .Y(_09389_));
 INVx1_ASAP7_75t_R _16605_ (.A(_00215_),
    .Y(_09390_));
 AO32x1_ASAP7_75t_R _16606_ (.A1(_09386_),
    .A2(_08987_),
    .A3(_09389_),
    .B1(_09360_),
    .B2(_09390_),
    .Y(_01368_));
 INVx1_ASAP7_75t_R _16607_ (.A(_00181_),
    .Y(_09391_));
 AND2x2_ASAP7_75t_R _16608_ (.A(_09252_),
    .B(_09359_),
    .Y(_09392_));
 AO22x1_ASAP7_75t_R _16609_ (.A1(_09391_),
    .A2(_09352_),
    .B1(_09392_),
    .B2(_09006_),
    .Y(_01369_));
 AND4x1_ASAP7_75t_R _16610_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09358_),
    .Y(_09393_));
 AO32x1_ASAP7_75t_R _16611_ (.A1(_09386_),
    .A2(_09025_),
    .A3(_09393_),
    .B1(_09360_),
    .B2(_04408_),
    .Y(_01370_));
 AND3x1_ASAP7_75t_R _16612_ (.A(_09259_),
    .B(_09260_),
    .C(_09364_),
    .Y(_09394_));
 INVx1_ASAP7_75t_R _16613_ (.A(_00114_),
    .Y(_09395_));
 AO32x1_ASAP7_75t_R _16614_ (.A1(_09386_),
    .A2(_09043_),
    .A3(_09394_),
    .B1(_09360_),
    .B2(_09395_),
    .Y(_01371_));
 NAND2x1_ASAP7_75t_R _16615_ (.A(_01011_),
    .B(_09352_),
    .Y(_09396_));
 OA21x2_ASAP7_75t_R _16616_ (.A1(_09263_),
    .A2(_09351_),
    .B(_09396_),
    .Y(_01372_));
 AND4x1_ASAP7_75t_R _16617_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09358_),
    .Y(_09397_));
 INVx1_ASAP7_75t_R _16618_ (.A(_00080_),
    .Y(_09398_));
 AO32x1_ASAP7_75t_R _16619_ (.A1(_09386_),
    .A2(_09070_),
    .A3(_09397_),
    .B1(_09360_),
    .B2(_09398_),
    .Y(_01373_));
 AND3x1_ASAP7_75t_R _16620_ (.A(_09270_),
    .B(_09271_),
    .C(_09364_),
    .Y(_09399_));
 INVx1_ASAP7_75t_R _16621_ (.A(_00048_),
    .Y(_09400_));
 AO32x1_ASAP7_75t_R _16622_ (.A1(_09386_),
    .A2(_09086_),
    .A3(_09399_),
    .B1(_09360_),
    .B2(_09400_),
    .Y(_01374_));
 NAND2x1_ASAP7_75t_R _16623_ (.A(_00978_),
    .B(_09352_),
    .Y(_09401_));
 OA21x2_ASAP7_75t_R _16624_ (.A1(_09274_),
    .A2(_09351_),
    .B(_09401_),
    .Y(_01375_));
 NAND2x1_ASAP7_75t_R _16625_ (.A(_00945_),
    .B(_09366_),
    .Y(_09402_));
 OA21x2_ASAP7_75t_R _16626_ (.A1(_09276_),
    .A2(_09351_),
    .B(_09402_),
    .Y(_01376_));
 AND2x2_ASAP7_75t_R _16627_ (.A(_00911_),
    .B(_09360_),
    .Y(_09403_));
 AOI21x1_ASAP7_75t_R _16628_ (.A1(_09137_),
    .A2(_09359_),
    .B(_09403_),
    .Y(_01377_));
 NOR2x1_ASAP7_75t_R _16629_ (.A(_00878_),
    .B(_09359_),
    .Y(_09404_));
 AO21x1_ASAP7_75t_R _16630_ (.A1(_09279_),
    .A2(_09359_),
    .B(_09404_),
    .Y(_01378_));
 NOR2x1_ASAP7_75t_R _16631_ (.A(_00844_),
    .B(_09359_),
    .Y(_09405_));
 AO21x1_ASAP7_75t_R _16632_ (.A1(_09281_),
    .A2(_09359_),
    .B(_09405_),
    .Y(_01379_));
 NOR2x1_ASAP7_75t_R _16633_ (.A(_00811_),
    .B(_09359_),
    .Y(_09406_));
 AO21x1_ASAP7_75t_R _16634_ (.A1(_09283_),
    .A2(_09359_),
    .B(_09406_),
    .Y(_01380_));
 NAND2x1_ASAP7_75t_R _16635_ (.A(_00777_),
    .B(_09366_),
    .Y(_09407_));
 OA21x2_ASAP7_75t_R _16636_ (.A1(_09285_),
    .A2(_09352_),
    .B(_09407_),
    .Y(_01381_));
 BUFx4f_ASAP7_75t_R _16637_ (.A(_08598_),
    .Y(_09408_));
 OR3x4_ASAP7_75t_R _16638_ (.A(_09408_),
    .B(_08601_),
    .C(_09291_),
    .Y(_09409_));
 BUFx10_ASAP7_75t_R _16639_ (.A(_09409_),
    .Y(_09410_));
 BUFx12_ASAP7_75t_R _16640_ (.A(_09409_),
    .Y(_09411_));
 NAND2x1_ASAP7_75t_R _16641_ (.A(_00014_),
    .B(_09411_),
    .Y(_09412_));
 OA21x2_ASAP7_75t_R _16642_ (.A1(_08597_),
    .A2(_09410_),
    .B(_09412_),
    .Y(_01382_));
 NAND2x1_ASAP7_75t_R _16643_ (.A(_00746_),
    .B(_09411_),
    .Y(_09413_));
 OA21x2_ASAP7_75t_R _16644_ (.A1(_09196_),
    .A2(_09410_),
    .B(_09413_),
    .Y(_01383_));
 NAND2x1_ASAP7_75t_R _16645_ (.A(_00713_),
    .B(_09411_),
    .Y(_09414_));
 OA21x2_ASAP7_75t_R _16646_ (.A1(_09198_),
    .A2(_09410_),
    .B(_09414_),
    .Y(_01384_));
 NAND2x1_ASAP7_75t_R _16647_ (.A(_00680_),
    .B(_09411_),
    .Y(_09415_));
 OA21x2_ASAP7_75t_R _16648_ (.A1(_09200_),
    .A2(_09410_),
    .B(_09415_),
    .Y(_01385_));
 OR2x6_ASAP7_75t_R _16649_ (.A(_09408_),
    .B(_08601_),
    .Y(_09416_));
 NOR2x2_ASAP7_75t_R _16650_ (.A(_09416_),
    .B(_09291_),
    .Y(_09417_));
 BUFx6f_ASAP7_75t_R _16651_ (.A(_09417_),
    .Y(_09418_));
 BUFx10_ASAP7_75t_R _16652_ (.A(_09409_),
    .Y(_09419_));
 AND2x2_ASAP7_75t_R _16653_ (.A(_00647_),
    .B(_09419_),
    .Y(_09420_));
 AOI21x1_ASAP7_75t_R _16654_ (.A1(_08725_),
    .A2(_09418_),
    .B(_09420_),
    .Y(_01386_));
 NAND2x1_ASAP7_75t_R _16655_ (.A(_00614_),
    .B(_09411_),
    .Y(_09421_));
 OA21x2_ASAP7_75t_R _16656_ (.A1(_09206_),
    .A2(_09410_),
    .B(_09421_),
    .Y(_01387_));
 OR2x2_ASAP7_75t_R _16657_ (.A(_00580_),
    .B(_09418_),
    .Y(_09422_));
 OAI21x1_ASAP7_75t_R _16658_ (.A1(_08766_),
    .A2(_09410_),
    .B(_09422_),
    .Y(_01388_));
 BUFx4f_ASAP7_75t_R _16659_ (.A(_09417_),
    .Y(_09423_));
 AND3x1_ASAP7_75t_R _16660_ (.A(_09210_),
    .B(_09211_),
    .C(_09423_),
    .Y(_09424_));
 BUFx10_ASAP7_75t_R _16661_ (.A(_09409_),
    .Y(_09425_));
 INVx1_ASAP7_75t_R _16662_ (.A(_00547_),
    .Y(_09426_));
 AO32x1_ASAP7_75t_R _16663_ (.A1(_08783_),
    .A2(_08785_),
    .A3(_09424_),
    .B1(_09425_),
    .B2(_09426_),
    .Y(_01389_));
 AND2x2_ASAP7_75t_R _16664_ (.A(_09215_),
    .B(_09423_),
    .Y(_09427_));
 INVx1_ASAP7_75t_R _16665_ (.A(_00514_),
    .Y(_09428_));
 AO32x1_ASAP7_75t_R _16666_ (.A1(_09386_),
    .A2(_08805_),
    .A3(_09427_),
    .B1(_09425_),
    .B2(_09428_),
    .Y(_01390_));
 AND3x1_ASAP7_75t_R _16667_ (.A(_09219_),
    .B(_09220_),
    .C(_09423_),
    .Y(_09429_));
 INVx1_ASAP7_75t_R _16668_ (.A(_00481_),
    .Y(_09430_));
 AO32x1_ASAP7_75t_R _16669_ (.A1(_09386_),
    .A2(_08830_),
    .A3(_09429_),
    .B1(_09425_),
    .B2(_09430_),
    .Y(_01391_));
 AND3x1_ASAP7_75t_R _16670_ (.A(_09223_),
    .B(_09224_),
    .C(_09423_),
    .Y(_09431_));
 INVx1_ASAP7_75t_R _16671_ (.A(_00448_),
    .Y(_09432_));
 AO32x1_ASAP7_75t_R _16672_ (.A1(_09386_),
    .A2(_08850_),
    .A3(_09431_),
    .B1(_09425_),
    .B2(_09432_),
    .Y(_01392_));
 NAND2x1_ASAP7_75t_R _16673_ (.A(_01045_),
    .B(_09411_),
    .Y(_09433_));
 OA21x2_ASAP7_75t_R _16674_ (.A1(_09227_),
    .A2(_09410_),
    .B(_09433_),
    .Y(_01393_));
 AND2x2_ASAP7_75t_R _16675_ (.A(_09229_),
    .B(_09423_),
    .Y(_09434_));
 INVx1_ASAP7_75t_R _16676_ (.A(_00415_),
    .Y(_09435_));
 AO32x1_ASAP7_75t_R _16677_ (.A1(_09386_),
    .A2(_08879_),
    .A3(_09434_),
    .B1(_09425_),
    .B2(_09435_),
    .Y(_01394_));
 BUFx3_ASAP7_75t_R _16678_ (.A(_09385_),
    .Y(_09436_));
 AND3x1_ASAP7_75t_R _16679_ (.A(_09232_),
    .B(_09233_),
    .C(_09423_),
    .Y(_09437_));
 INVx1_ASAP7_75t_R _16680_ (.A(_00382_),
    .Y(_09438_));
 AO32x1_ASAP7_75t_R _16681_ (.A1(_09436_),
    .A2(_08901_),
    .A3(_09437_),
    .B1(_09425_),
    .B2(_09438_),
    .Y(_01395_));
 AND2x2_ASAP7_75t_R _16682_ (.A(_09236_),
    .B(_09423_),
    .Y(_09439_));
 INVx1_ASAP7_75t_R _16683_ (.A(_00349_),
    .Y(_09440_));
 AO32x1_ASAP7_75t_R _16684_ (.A1(_09436_),
    .A2(_08918_),
    .A3(_09439_),
    .B1(_09425_),
    .B2(_09440_),
    .Y(_01396_));
 AND2x2_ASAP7_75t_R _16685_ (.A(_09240_),
    .B(_09423_),
    .Y(_09441_));
 INVx1_ASAP7_75t_R _16686_ (.A(_00315_),
    .Y(_09442_));
 AO32x1_ASAP7_75t_R _16687_ (.A1(_09436_),
    .A2(_08937_),
    .A3(_09441_),
    .B1(_09425_),
    .B2(_09442_),
    .Y(_01397_));
 AND2x2_ASAP7_75t_R _16688_ (.A(_09243_),
    .B(_09417_),
    .Y(_09443_));
 INVx1_ASAP7_75t_R _16689_ (.A(_00282_),
    .Y(_09444_));
 AO32x1_ASAP7_75t_R _16690_ (.A1(_09436_),
    .A2(_08951_),
    .A3(_09443_),
    .B1(_09419_),
    .B2(_09444_),
    .Y(_01398_));
 AND2x2_ASAP7_75t_R _16691_ (.A(_09246_),
    .B(_09417_),
    .Y(_09445_));
 INVx1_ASAP7_75t_R _16692_ (.A(_00249_),
    .Y(_09446_));
 AO32x1_ASAP7_75t_R _16693_ (.A1(_09436_),
    .A2(_08970_),
    .A3(_09445_),
    .B1(_09419_),
    .B2(_09446_),
    .Y(_01399_));
 NOR2x1_ASAP7_75t_R _16694_ (.A(_08997_),
    .B(_09419_),
    .Y(_09447_));
 INVx1_ASAP7_75t_R _16695_ (.A(_00216_),
    .Y(_09448_));
 AO32x1_ASAP7_75t_R _16696_ (.A1(_09436_),
    .A2(_08987_),
    .A3(_09447_),
    .B1(_09419_),
    .B2(_09448_),
    .Y(_01400_));
 INVx1_ASAP7_75t_R _16697_ (.A(_00182_),
    .Y(_09449_));
 AND2x2_ASAP7_75t_R _16698_ (.A(_09252_),
    .B(_09418_),
    .Y(_09450_));
 AO22x1_ASAP7_75t_R _16699_ (.A1(_09449_),
    .A2(_09411_),
    .B1(_09450_),
    .B2(_09006_),
    .Y(_01401_));
 AND4x1_ASAP7_75t_R _16700_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09417_),
    .Y(_09451_));
 AO32x1_ASAP7_75t_R _16701_ (.A1(_09436_),
    .A2(_09025_),
    .A3(_09451_),
    .B1(_09419_),
    .B2(_04402_),
    .Y(_01402_));
 AND3x1_ASAP7_75t_R _16702_ (.A(_09259_),
    .B(_09260_),
    .C(_09423_),
    .Y(_09452_));
 INVx1_ASAP7_75t_R _16703_ (.A(_00115_),
    .Y(_09453_));
 AO32x1_ASAP7_75t_R _16704_ (.A1(_09436_),
    .A2(_09043_),
    .A3(_09452_),
    .B1(_09419_),
    .B2(_09453_),
    .Y(_01403_));
 NAND2x1_ASAP7_75t_R _16705_ (.A(_01012_),
    .B(_09411_),
    .Y(_09454_));
 OA21x2_ASAP7_75t_R _16706_ (.A1(_09263_),
    .A2(_09410_),
    .B(_09454_),
    .Y(_01404_));
 AND4x1_ASAP7_75t_R _16707_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09417_),
    .Y(_09455_));
 INVx1_ASAP7_75t_R _16708_ (.A(_00081_),
    .Y(_09456_));
 AO32x1_ASAP7_75t_R _16709_ (.A1(_09436_),
    .A2(_09070_),
    .A3(_09455_),
    .B1(_09419_),
    .B2(_09456_),
    .Y(_01405_));
 AND3x1_ASAP7_75t_R _16710_ (.A(_09270_),
    .B(_09271_),
    .C(_09423_),
    .Y(_09457_));
 INVx1_ASAP7_75t_R _16711_ (.A(_00049_),
    .Y(_09458_));
 AO32x1_ASAP7_75t_R _16712_ (.A1(_09436_),
    .A2(_09086_),
    .A3(_09457_),
    .B1(_09419_),
    .B2(_09458_),
    .Y(_01406_));
 NAND2x1_ASAP7_75t_R _16713_ (.A(_00979_),
    .B(_09411_),
    .Y(_09459_));
 OA21x2_ASAP7_75t_R _16714_ (.A1(_09274_),
    .A2(_09410_),
    .B(_09459_),
    .Y(_01407_));
 NAND2x1_ASAP7_75t_R _16715_ (.A(_00946_),
    .B(_09425_),
    .Y(_09460_));
 OA21x2_ASAP7_75t_R _16716_ (.A1(_09276_),
    .A2(_09410_),
    .B(_09460_),
    .Y(_01408_));
 AND2x2_ASAP7_75t_R _16717_ (.A(_00912_),
    .B(_09419_),
    .Y(_09461_));
 AOI21x1_ASAP7_75t_R _16718_ (.A1(_09137_),
    .A2(_09418_),
    .B(_09461_),
    .Y(_01409_));
 NOR2x1_ASAP7_75t_R _16719_ (.A(_00879_),
    .B(_09418_),
    .Y(_09462_));
 AO21x1_ASAP7_75t_R _16720_ (.A1(_09279_),
    .A2(_09418_),
    .B(_09462_),
    .Y(_01410_));
 NOR2x1_ASAP7_75t_R _16721_ (.A(_00845_),
    .B(_09418_),
    .Y(_09463_));
 AO21x1_ASAP7_75t_R _16722_ (.A1(_09281_),
    .A2(_09418_),
    .B(_09463_),
    .Y(_01411_));
 NOR2x1_ASAP7_75t_R _16723_ (.A(_00812_),
    .B(_09418_),
    .Y(_09464_));
 AO21x1_ASAP7_75t_R _16724_ (.A1(_09283_),
    .A2(_09418_),
    .B(_09464_),
    .Y(_01412_));
 NAND2x1_ASAP7_75t_R _16725_ (.A(_00778_),
    .B(_09425_),
    .Y(_09465_));
 OA21x2_ASAP7_75t_R _16726_ (.A1(_09285_),
    .A2(_09411_),
    .B(_09465_),
    .Y(_01413_));
 OR3x4_ASAP7_75t_R _16727_ (.A(_09408_),
    .B(_09349_),
    .C(_09291_),
    .Y(_09466_));
 BUFx6f_ASAP7_75t_R _16728_ (.A(_09466_),
    .Y(_09467_));
 BUFx10_ASAP7_75t_R _16729_ (.A(_09466_),
    .Y(_09468_));
 NAND2x1_ASAP7_75t_R _16730_ (.A(_00015_),
    .B(_09468_),
    .Y(_09469_));
 OA21x2_ASAP7_75t_R _16731_ (.A1(_08597_),
    .A2(_09467_),
    .B(_09469_),
    .Y(_01414_));
 NAND2x1_ASAP7_75t_R _16732_ (.A(_00747_),
    .B(_09468_),
    .Y(_09470_));
 OA21x2_ASAP7_75t_R _16733_ (.A1(_09196_),
    .A2(_09467_),
    .B(_09470_),
    .Y(_01415_));
 NAND2x1_ASAP7_75t_R _16734_ (.A(_00714_),
    .B(_09468_),
    .Y(_09471_));
 OA21x2_ASAP7_75t_R _16735_ (.A1(_09198_),
    .A2(_09467_),
    .B(_09471_),
    .Y(_01416_));
 NAND2x1_ASAP7_75t_R _16736_ (.A(_00681_),
    .B(_09468_),
    .Y(_09472_));
 OA21x2_ASAP7_75t_R _16737_ (.A1(_09200_),
    .A2(_09467_),
    .B(_09472_),
    .Y(_01417_));
 OR2x6_ASAP7_75t_R _16738_ (.A(_09408_),
    .B(_09349_),
    .Y(_09473_));
 NOR2x2_ASAP7_75t_R _16739_ (.A(_09473_),
    .B(_09291_),
    .Y(_09474_));
 BUFx6f_ASAP7_75t_R _16740_ (.A(_09474_),
    .Y(_09475_));
 BUFx10_ASAP7_75t_R _16741_ (.A(_09466_),
    .Y(_09476_));
 AND2x2_ASAP7_75t_R _16742_ (.A(_00648_),
    .B(_09476_),
    .Y(_09477_));
 AOI21x1_ASAP7_75t_R _16743_ (.A1(_08725_),
    .A2(_09475_),
    .B(_09477_),
    .Y(_01418_));
 NAND2x1_ASAP7_75t_R _16744_ (.A(_00615_),
    .B(_09468_),
    .Y(_09478_));
 OA21x2_ASAP7_75t_R _16745_ (.A1(_09206_),
    .A2(_09467_),
    .B(_09478_),
    .Y(_01419_));
 OR2x2_ASAP7_75t_R _16746_ (.A(_00581_),
    .B(_09475_),
    .Y(_09479_));
 OAI21x1_ASAP7_75t_R _16747_ (.A1(_08766_),
    .A2(_09467_),
    .B(_09479_),
    .Y(_01420_));
 BUFx4f_ASAP7_75t_R _16748_ (.A(_09474_),
    .Y(_09480_));
 AND3x1_ASAP7_75t_R _16749_ (.A(_09210_),
    .B(_09211_),
    .C(_09480_),
    .Y(_09481_));
 BUFx10_ASAP7_75t_R _16750_ (.A(_09466_),
    .Y(_09482_));
 INVx1_ASAP7_75t_R _16751_ (.A(_00548_),
    .Y(_09483_));
 AO32x1_ASAP7_75t_R _16752_ (.A1(_08783_),
    .A2(_08785_),
    .A3(_09481_),
    .B1(_09482_),
    .B2(_09483_),
    .Y(_01421_));
 BUFx3_ASAP7_75t_R _16753_ (.A(_09385_),
    .Y(_09484_));
 AND2x2_ASAP7_75t_R _16754_ (.A(_09215_),
    .B(_09480_),
    .Y(_09485_));
 INVx1_ASAP7_75t_R _16755_ (.A(_00515_),
    .Y(_09486_));
 AO32x1_ASAP7_75t_R _16756_ (.A1(_09484_),
    .A2(_08805_),
    .A3(_09485_),
    .B1(_09482_),
    .B2(_09486_),
    .Y(_01422_));
 AND3x1_ASAP7_75t_R _16757_ (.A(_09219_),
    .B(_09220_),
    .C(_09480_),
    .Y(_09487_));
 INVx1_ASAP7_75t_R _16758_ (.A(_00482_),
    .Y(_09488_));
 AO32x1_ASAP7_75t_R _16759_ (.A1(_09484_),
    .A2(_08830_),
    .A3(_09487_),
    .B1(_09482_),
    .B2(_09488_),
    .Y(_01423_));
 AND3x1_ASAP7_75t_R _16760_ (.A(_09223_),
    .B(_09224_),
    .C(_09480_),
    .Y(_09489_));
 INVx1_ASAP7_75t_R _16761_ (.A(_00449_),
    .Y(_09490_));
 AO32x1_ASAP7_75t_R _16762_ (.A1(_09484_),
    .A2(_08850_),
    .A3(_09489_),
    .B1(_09482_),
    .B2(_09490_),
    .Y(_01424_));
 NAND2x1_ASAP7_75t_R _16763_ (.A(_01046_),
    .B(_09468_),
    .Y(_09491_));
 OA21x2_ASAP7_75t_R _16764_ (.A1(_09227_),
    .A2(_09467_),
    .B(_09491_),
    .Y(_01425_));
 AND2x2_ASAP7_75t_R _16765_ (.A(_09229_),
    .B(_09480_),
    .Y(_09492_));
 INVx1_ASAP7_75t_R _16766_ (.A(_00416_),
    .Y(_09493_));
 AO32x1_ASAP7_75t_R _16767_ (.A1(_09484_),
    .A2(_08879_),
    .A3(_09492_),
    .B1(_09482_),
    .B2(_09493_),
    .Y(_01426_));
 AND3x1_ASAP7_75t_R _16768_ (.A(_09232_),
    .B(_09233_),
    .C(_09480_),
    .Y(_09494_));
 INVx1_ASAP7_75t_R _16769_ (.A(_00383_),
    .Y(_09495_));
 AO32x1_ASAP7_75t_R _16770_ (.A1(_09484_),
    .A2(_08901_),
    .A3(_09494_),
    .B1(_09482_),
    .B2(_09495_),
    .Y(_01427_));
 AND2x2_ASAP7_75t_R _16771_ (.A(_09236_),
    .B(_09480_),
    .Y(_09496_));
 INVx1_ASAP7_75t_R _16772_ (.A(_00350_),
    .Y(_09497_));
 AO32x1_ASAP7_75t_R _16773_ (.A1(_09484_),
    .A2(_08918_),
    .A3(_09496_),
    .B1(_09482_),
    .B2(_09497_),
    .Y(_01428_));
 AND2x2_ASAP7_75t_R _16774_ (.A(_09240_),
    .B(_09480_),
    .Y(_09498_));
 INVx1_ASAP7_75t_R _16775_ (.A(_00316_),
    .Y(_09499_));
 AO32x1_ASAP7_75t_R _16776_ (.A1(_09484_),
    .A2(_08937_),
    .A3(_09498_),
    .B1(_09482_),
    .B2(_09499_),
    .Y(_01429_));
 AND2x2_ASAP7_75t_R _16777_ (.A(_09243_),
    .B(_09474_),
    .Y(_09500_));
 INVx1_ASAP7_75t_R _16778_ (.A(_00283_),
    .Y(_09501_));
 AO32x1_ASAP7_75t_R _16779_ (.A1(_09484_),
    .A2(_08951_),
    .A3(_09500_),
    .B1(_09476_),
    .B2(_09501_),
    .Y(_01430_));
 AND2x2_ASAP7_75t_R _16780_ (.A(_09246_),
    .B(_09474_),
    .Y(_09502_));
 INVx1_ASAP7_75t_R _16781_ (.A(_00250_),
    .Y(_09503_));
 AO32x1_ASAP7_75t_R _16782_ (.A1(_09484_),
    .A2(_08970_),
    .A3(_09502_),
    .B1(_09476_),
    .B2(_09503_),
    .Y(_01431_));
 NOR2x1_ASAP7_75t_R _16783_ (.A(_08997_),
    .B(_09476_),
    .Y(_09504_));
 INVx1_ASAP7_75t_R _16784_ (.A(_00217_),
    .Y(_09505_));
 AO32x1_ASAP7_75t_R _16785_ (.A1(_09484_),
    .A2(_08987_),
    .A3(_09504_),
    .B1(_09476_),
    .B2(_09505_),
    .Y(_01432_));
 INVx1_ASAP7_75t_R _16786_ (.A(_00183_),
    .Y(_09506_));
 AND2x2_ASAP7_75t_R _16787_ (.A(_09252_),
    .B(_09475_),
    .Y(_09507_));
 AO22x1_ASAP7_75t_R _16788_ (.A1(_09506_),
    .A2(_09468_),
    .B1(_09507_),
    .B2(_09006_),
    .Y(_01433_));
 BUFx4f_ASAP7_75t_R _16789_ (.A(_09385_),
    .Y(_09508_));
 AND4x1_ASAP7_75t_R _16790_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09474_),
    .Y(_09509_));
 INVx1_ASAP7_75t_R _16791_ (.A(_00150_),
    .Y(_09510_));
 AO32x1_ASAP7_75t_R _16792_ (.A1(_09508_),
    .A2(_09025_),
    .A3(_09509_),
    .B1(_09476_),
    .B2(_09510_),
    .Y(_01434_));
 AND3x1_ASAP7_75t_R _16793_ (.A(_09259_),
    .B(_09260_),
    .C(_09480_),
    .Y(_09511_));
 INVx1_ASAP7_75t_R _16794_ (.A(_00116_),
    .Y(_09512_));
 AO32x1_ASAP7_75t_R _16795_ (.A1(_09508_),
    .A2(_09043_),
    .A3(_09511_),
    .B1(_09476_),
    .B2(_09512_),
    .Y(_01435_));
 NAND2x1_ASAP7_75t_R _16796_ (.A(_01013_),
    .B(_09468_),
    .Y(_09513_));
 OA21x2_ASAP7_75t_R _16797_ (.A1(_09263_),
    .A2(_09467_),
    .B(_09513_),
    .Y(_01436_));
 AND4x1_ASAP7_75t_R _16798_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09474_),
    .Y(_09514_));
 INVx1_ASAP7_75t_R _16799_ (.A(_00082_),
    .Y(_09515_));
 AO32x1_ASAP7_75t_R _16800_ (.A1(_09508_),
    .A2(_09070_),
    .A3(_09514_),
    .B1(_09476_),
    .B2(_09515_),
    .Y(_01437_));
 AND3x1_ASAP7_75t_R _16801_ (.A(_09270_),
    .B(_09271_),
    .C(_09480_),
    .Y(_09516_));
 INVx1_ASAP7_75t_R _16802_ (.A(_00050_),
    .Y(_09517_));
 AO32x1_ASAP7_75t_R _16803_ (.A1(_09508_),
    .A2(_09086_),
    .A3(_09516_),
    .B1(_09476_),
    .B2(_09517_),
    .Y(_01438_));
 NAND2x1_ASAP7_75t_R _16804_ (.A(_00980_),
    .B(_09468_),
    .Y(_09518_));
 OA21x2_ASAP7_75t_R _16805_ (.A1(_09274_),
    .A2(_09467_),
    .B(_09518_),
    .Y(_01439_));
 NAND2x1_ASAP7_75t_R _16806_ (.A(_00947_),
    .B(_09482_),
    .Y(_09519_));
 OA21x2_ASAP7_75t_R _16807_ (.A1(_09276_),
    .A2(_09467_),
    .B(_09519_),
    .Y(_01440_));
 AND2x2_ASAP7_75t_R _16808_ (.A(_00913_),
    .B(_09476_),
    .Y(_09520_));
 AOI21x1_ASAP7_75t_R _16809_ (.A1(_09137_),
    .A2(_09475_),
    .B(_09520_),
    .Y(_01441_));
 NOR2x1_ASAP7_75t_R _16810_ (.A(_00880_),
    .B(_09475_),
    .Y(_09521_));
 AO21x1_ASAP7_75t_R _16811_ (.A1(_09279_),
    .A2(_09475_),
    .B(_09521_),
    .Y(_01442_));
 NOR2x1_ASAP7_75t_R _16812_ (.A(_00846_),
    .B(_09475_),
    .Y(_09522_));
 AO21x1_ASAP7_75t_R _16813_ (.A1(_09281_),
    .A2(_09475_),
    .B(_09522_),
    .Y(_01443_));
 NOR2x1_ASAP7_75t_R _16814_ (.A(_00813_),
    .B(_09475_),
    .Y(_09523_));
 AO21x1_ASAP7_75t_R _16815_ (.A1(_09283_),
    .A2(_09475_),
    .B(_09523_),
    .Y(_01444_));
 NAND2x1_ASAP7_75t_R _16816_ (.A(_00779_),
    .B(_09482_),
    .Y(_09524_));
 OA21x2_ASAP7_75t_R _16817_ (.A1(_09285_),
    .A2(_09468_),
    .B(_09524_),
    .Y(_01445_));
 NAND2x1_ASAP7_75t_R _16818_ (.A(_03574_),
    .B(_08600_),
    .Y(_09525_));
 INVx2_ASAP7_75t_R _16819_ (.A(_09288_),
    .Y(_09526_));
 AND4x2_ASAP7_75t_R _16820_ (.A(_09188_),
    .B(_08598_),
    .C(_09525_),
    .D(_09526_),
    .Y(_09527_));
 BUFx12f_ASAP7_75t_R _16821_ (.A(_09527_),
    .Y(_09528_));
 BUFx10_ASAP7_75t_R _16822_ (.A(_09528_),
    .Y(_09529_));
 AND2x2_ASAP7_75t_R _16823_ (.A(_03566_),
    .B(_07020_),
    .Y(_09530_));
 AND3x4_ASAP7_75t_R _16824_ (.A(_08604_),
    .B(_06807_),
    .C(_09530_),
    .Y(_09531_));
 BUFx12f_ASAP7_75t_R _16825_ (.A(_09531_),
    .Y(_09532_));
 NAND2x2_ASAP7_75t_R _16826_ (.A(_09529_),
    .B(_09532_),
    .Y(_09533_));
 BUFx6f_ASAP7_75t_R _16827_ (.A(_09533_),
    .Y(_09534_));
 BUFx12_ASAP7_75t_R _16828_ (.A(_09533_),
    .Y(_09535_));
 NAND2x1_ASAP7_75t_R _16829_ (.A(_00016_),
    .B(_09535_),
    .Y(_09536_));
 OA21x2_ASAP7_75t_R _16830_ (.A1(_08597_),
    .A2(_09534_),
    .B(_09536_),
    .Y(_01446_));
 NAND2x1_ASAP7_75t_R _16831_ (.A(_00748_),
    .B(_09535_),
    .Y(_09537_));
 OA21x2_ASAP7_75t_R _16832_ (.A1(_09196_),
    .A2(_09534_),
    .B(_09537_),
    .Y(_01447_));
 NAND2x1_ASAP7_75t_R _16833_ (.A(_00715_),
    .B(_09535_),
    .Y(_09538_));
 OA21x2_ASAP7_75t_R _16834_ (.A1(_09198_),
    .A2(_09534_),
    .B(_09538_),
    .Y(_01448_));
 NAND2x1_ASAP7_75t_R _16835_ (.A(_00682_),
    .B(_09535_),
    .Y(_09539_));
 OA21x2_ASAP7_75t_R _16836_ (.A1(_09200_),
    .A2(_09534_),
    .B(_09539_),
    .Y(_01449_));
 AND2x6_ASAP7_75t_R _16837_ (.A(_09528_),
    .B(_09531_),
    .Y(_09540_));
 BUFx6f_ASAP7_75t_R _16838_ (.A(_09540_),
    .Y(_09541_));
 AND2x2_ASAP7_75t_R _16839_ (.A(_00649_),
    .B(_09533_),
    .Y(_09542_));
 AOI21x1_ASAP7_75t_R _16840_ (.A1(_08725_),
    .A2(_09541_),
    .B(_09542_),
    .Y(_01450_));
 BUFx6f_ASAP7_75t_R _16841_ (.A(_09529_),
    .Y(_09543_));
 BUFx6f_ASAP7_75t_R _16842_ (.A(_09532_),
    .Y(_09544_));
 AO21x1_ASAP7_75t_R _16843_ (.A1(_09543_),
    .A2(_09544_),
    .B(_05892_),
    .Y(_09545_));
 OA21x2_ASAP7_75t_R _16844_ (.A1(_09206_),
    .A2(_09534_),
    .B(_09545_),
    .Y(_01451_));
 AO21x1_ASAP7_75t_R _16845_ (.A1(_09543_),
    .A2(_09544_),
    .B(_00582_),
    .Y(_09546_));
 OAI21x1_ASAP7_75t_R _16846_ (.A1(_08766_),
    .A2(_09534_),
    .B(_09546_),
    .Y(_01452_));
 BUFx6f_ASAP7_75t_R _16847_ (.A(_08784_),
    .Y(_09547_));
 BUFx6f_ASAP7_75t_R _16848_ (.A(_09547_),
    .Y(_09548_));
 AND3x1_ASAP7_75t_R _16849_ (.A(_09210_),
    .B(_09211_),
    .C(_09541_),
    .Y(_09549_));
 AO32x1_ASAP7_75t_R _16850_ (.A1(_08783_),
    .A2(_09548_),
    .A3(_09549_),
    .B1(_09535_),
    .B2(_05660_),
    .Y(_01453_));
 BUFx4f_ASAP7_75t_R _16851_ (.A(_09540_),
    .Y(_09550_));
 AND2x2_ASAP7_75t_R _16852_ (.A(_09215_),
    .B(_09550_),
    .Y(_09551_));
 BUFx3_ASAP7_75t_R _16853_ (.A(_09533_),
    .Y(_09552_));
 INVx1_ASAP7_75t_R _16854_ (.A(_00516_),
    .Y(_09553_));
 AO32x1_ASAP7_75t_R _16855_ (.A1(_09508_),
    .A2(_08805_),
    .A3(_09551_),
    .B1(_09552_),
    .B2(_09553_),
    .Y(_01454_));
 AND3x1_ASAP7_75t_R _16856_ (.A(_09219_),
    .B(_09220_),
    .C(_09550_),
    .Y(_09554_));
 INVx1_ASAP7_75t_R _16857_ (.A(_00483_),
    .Y(_09555_));
 AO32x1_ASAP7_75t_R _16858_ (.A1(_09508_),
    .A2(_08830_),
    .A3(_09554_),
    .B1(_09552_),
    .B2(_09555_),
    .Y(_01455_));
 AND3x1_ASAP7_75t_R _16859_ (.A(_09223_),
    .B(_09224_),
    .C(_09550_),
    .Y(_09556_));
 INVx1_ASAP7_75t_R _16860_ (.A(_00450_),
    .Y(_09557_));
 AO32x1_ASAP7_75t_R _16861_ (.A1(_09508_),
    .A2(_08850_),
    .A3(_09556_),
    .B1(_09552_),
    .B2(_09557_),
    .Y(_01456_));
 AO21x1_ASAP7_75t_R _16862_ (.A1(_09543_),
    .A2(_09544_),
    .B(_07213_),
    .Y(_09558_));
 OA21x2_ASAP7_75t_R _16863_ (.A1(_09227_),
    .A2(_09534_),
    .B(_09558_),
    .Y(_01457_));
 AND2x2_ASAP7_75t_R _16864_ (.A(_09229_),
    .B(_09550_),
    .Y(_09559_));
 INVx1_ASAP7_75t_R _16865_ (.A(_00417_),
    .Y(_09560_));
 AO32x1_ASAP7_75t_R _16866_ (.A1(_09508_),
    .A2(_08879_),
    .A3(_09559_),
    .B1(_09552_),
    .B2(_09560_),
    .Y(_01458_));
 AND3x1_ASAP7_75t_R _16867_ (.A(_09232_),
    .B(_09233_),
    .C(_09550_),
    .Y(_09561_));
 AO32x1_ASAP7_75t_R _16868_ (.A1(_09508_),
    .A2(_08901_),
    .A3(_09561_),
    .B1(_09552_),
    .B2(_05175_),
    .Y(_01459_));
 AND2x2_ASAP7_75t_R _16869_ (.A(_09236_),
    .B(_09550_),
    .Y(_09562_));
 INVx1_ASAP7_75t_R _16870_ (.A(_00351_),
    .Y(_09563_));
 AO32x1_ASAP7_75t_R _16871_ (.A1(_09508_),
    .A2(_08918_),
    .A3(_09562_),
    .B1(_09552_),
    .B2(_09563_),
    .Y(_01460_));
 BUFx4f_ASAP7_75t_R _16872_ (.A(_09385_),
    .Y(_09564_));
 AND2x2_ASAP7_75t_R _16873_ (.A(_09240_),
    .B(_09550_),
    .Y(_09565_));
 INVx1_ASAP7_75t_R _16874_ (.A(_00317_),
    .Y(_09566_));
 AO32x1_ASAP7_75t_R _16875_ (.A1(_09564_),
    .A2(_08937_),
    .A3(_09565_),
    .B1(_09552_),
    .B2(_09566_),
    .Y(_01461_));
 AND2x2_ASAP7_75t_R _16876_ (.A(_09243_),
    .B(_09550_),
    .Y(_09567_));
 INVx1_ASAP7_75t_R _16877_ (.A(_00284_),
    .Y(_09568_));
 AO32x1_ASAP7_75t_R _16878_ (.A1(_09564_),
    .A2(_08951_),
    .A3(_09567_),
    .B1(_09552_),
    .B2(_09568_),
    .Y(_01462_));
 AND2x2_ASAP7_75t_R _16879_ (.A(_09246_),
    .B(_09540_),
    .Y(_09569_));
 INVx1_ASAP7_75t_R _16880_ (.A(_00251_),
    .Y(_09570_));
 AO32x1_ASAP7_75t_R _16881_ (.A1(_09564_),
    .A2(_08970_),
    .A3(_09569_),
    .B1(_09552_),
    .B2(_09570_),
    .Y(_01463_));
 NOR2x1_ASAP7_75t_R _16882_ (.A(_08997_),
    .B(_09533_),
    .Y(_09571_));
 INVx1_ASAP7_75t_R _16883_ (.A(_00218_),
    .Y(_09572_));
 AO32x1_ASAP7_75t_R _16884_ (.A1(_09564_),
    .A2(_08987_),
    .A3(_09571_),
    .B1(_09552_),
    .B2(_09572_),
    .Y(_01464_));
 INVx1_ASAP7_75t_R _16885_ (.A(_00184_),
    .Y(_09573_));
 AND2x2_ASAP7_75t_R _16886_ (.A(_09252_),
    .B(_09541_),
    .Y(_09574_));
 AO22x1_ASAP7_75t_R _16887_ (.A1(_09573_),
    .A2(_09535_),
    .B1(_09574_),
    .B2(_09006_),
    .Y(_01465_));
 AND4x1_ASAP7_75t_R _16888_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09540_),
    .Y(_09575_));
 AO32x1_ASAP7_75t_R _16889_ (.A1(_09564_),
    .A2(_09025_),
    .A3(_09575_),
    .B1(_09533_),
    .B2(_04497_),
    .Y(_01466_));
 AND3x1_ASAP7_75t_R _16890_ (.A(_09259_),
    .B(_09260_),
    .C(_09550_),
    .Y(_09576_));
 INVx1_ASAP7_75t_R _16891_ (.A(_00117_),
    .Y(_09577_));
 AO32x1_ASAP7_75t_R _16892_ (.A1(_09564_),
    .A2(_09043_),
    .A3(_09576_),
    .B1(_09533_),
    .B2(_09577_),
    .Y(_01467_));
 AO21x1_ASAP7_75t_R _16893_ (.A1(_09543_),
    .A2(_09544_),
    .B(_07068_),
    .Y(_09578_));
 OA21x2_ASAP7_75t_R _16894_ (.A1(_09263_),
    .A2(_09534_),
    .B(_09578_),
    .Y(_01468_));
 AND4x1_ASAP7_75t_R _16895_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09540_),
    .Y(_09579_));
 INVx1_ASAP7_75t_R _16896_ (.A(_00083_),
    .Y(_09580_));
 AO32x1_ASAP7_75t_R _16897_ (.A1(_09564_),
    .A2(_09070_),
    .A3(_09579_),
    .B1(_09533_),
    .B2(_09580_),
    .Y(_01469_));
 AND3x1_ASAP7_75t_R _16898_ (.A(_09270_),
    .B(_09271_),
    .C(_09550_),
    .Y(_09581_));
 AO32x1_ASAP7_75t_R _16899_ (.A1(_09564_),
    .A2(_09086_),
    .A3(_09581_),
    .B1(_09533_),
    .B2(_03788_),
    .Y(_01470_));
 NAND2x1_ASAP7_75t_R _16900_ (.A(_00981_),
    .B(_09535_),
    .Y(_09582_));
 OA21x2_ASAP7_75t_R _16901_ (.A1(_09274_),
    .A2(_09534_),
    .B(_09582_),
    .Y(_01471_));
 NAND2x1_ASAP7_75t_R _16902_ (.A(_00948_),
    .B(_09535_),
    .Y(_09583_));
 OA21x2_ASAP7_75t_R _16903_ (.A1(_09276_),
    .A2(_09534_),
    .B(_09583_),
    .Y(_01472_));
 AND2x2_ASAP7_75t_R _16904_ (.A(_00914_),
    .B(_09533_),
    .Y(_09584_));
 AOI21x1_ASAP7_75t_R _16905_ (.A1(_09137_),
    .A2(_09541_),
    .B(_09584_),
    .Y(_01473_));
 NOR2x1_ASAP7_75t_R _16906_ (.A(_00881_),
    .B(_09541_),
    .Y(_09585_));
 AO21x1_ASAP7_75t_R _16907_ (.A1(_09279_),
    .A2(_09541_),
    .B(_09585_),
    .Y(_01474_));
 NOR2x1_ASAP7_75t_R _16908_ (.A(_00847_),
    .B(_09541_),
    .Y(_09586_));
 AO21x1_ASAP7_75t_R _16909_ (.A1(_09281_),
    .A2(_09541_),
    .B(_09586_),
    .Y(_01475_));
 NOR2x1_ASAP7_75t_R _16910_ (.A(_00814_),
    .B(_09541_),
    .Y(_09587_));
 AO21x1_ASAP7_75t_R _16911_ (.A1(_09283_),
    .A2(_09541_),
    .B(_09587_),
    .Y(_01476_));
 NAND2x1_ASAP7_75t_R _16912_ (.A(_00780_),
    .B(_09535_),
    .Y(_09588_));
 OA21x2_ASAP7_75t_R _16913_ (.A1(_09285_),
    .A2(_09535_),
    .B(_09588_),
    .Y(_01477_));
 NOR2x2_ASAP7_75t_R _16914_ (.A(_07131_),
    .B(_09189_),
    .Y(_09589_));
 BUFx16f_ASAP7_75t_R _16915_ (.A(_09589_),
    .Y(_09590_));
 NAND2x2_ASAP7_75t_R _16916_ (.A(_09590_),
    .B(_09532_),
    .Y(_09591_));
 BUFx10_ASAP7_75t_R _16917_ (.A(_09591_),
    .Y(_09592_));
 BUFx6f_ASAP7_75t_R _16918_ (.A(_09592_),
    .Y(_09593_));
 BUFx12f_ASAP7_75t_R _16919_ (.A(_09591_),
    .Y(_09594_));
 NAND2x1_ASAP7_75t_R _16920_ (.A(_00017_),
    .B(_09594_),
    .Y(_09595_));
 OA21x2_ASAP7_75t_R _16921_ (.A1(_08597_),
    .A2(_09593_),
    .B(_09595_),
    .Y(_01478_));
 NAND2x1_ASAP7_75t_R _16922_ (.A(_00749_),
    .B(_09594_),
    .Y(_09596_));
 OA21x2_ASAP7_75t_R _16923_ (.A1(_09196_),
    .A2(_09593_),
    .B(_09596_),
    .Y(_01479_));
 BUFx6f_ASAP7_75t_R _16924_ (.A(_09590_),
    .Y(_09597_));
 AO21x1_ASAP7_75t_R _16925_ (.A1(_09597_),
    .A2(_09544_),
    .B(_06221_),
    .Y(_09598_));
 OA21x2_ASAP7_75t_R _16926_ (.A1(_09198_),
    .A2(_09593_),
    .B(_09598_),
    .Y(_01480_));
 AO21x1_ASAP7_75t_R _16927_ (.A1(_09597_),
    .A2(_09544_),
    .B(_06104_),
    .Y(_09599_));
 OA21x2_ASAP7_75t_R _16928_ (.A1(_09200_),
    .A2(_09593_),
    .B(_09599_),
    .Y(_01481_));
 AND2x4_ASAP7_75t_R _16929_ (.A(_09589_),
    .B(_09531_),
    .Y(_09600_));
 BUFx6f_ASAP7_75t_R _16930_ (.A(_09600_),
    .Y(_09601_));
 AND2x2_ASAP7_75t_R _16931_ (.A(_00650_),
    .B(_09592_),
    .Y(_09602_));
 AOI21x1_ASAP7_75t_R _16932_ (.A1(_08725_),
    .A2(_09601_),
    .B(_09602_),
    .Y(_01482_));
 NAND2x1_ASAP7_75t_R _16933_ (.A(_00617_),
    .B(_09594_),
    .Y(_09603_));
 OA21x2_ASAP7_75t_R _16934_ (.A1(_09206_),
    .A2(_09593_),
    .B(_09603_),
    .Y(_01483_));
 AO21x1_ASAP7_75t_R _16935_ (.A1(_09597_),
    .A2(_09544_),
    .B(_00583_),
    .Y(_09604_));
 OAI21x1_ASAP7_75t_R _16936_ (.A1(_08766_),
    .A2(_09593_),
    .B(_09604_),
    .Y(_01484_));
 AND3x1_ASAP7_75t_R _16937_ (.A(_09210_),
    .B(_09211_),
    .C(_09601_),
    .Y(_09605_));
 AO32x1_ASAP7_75t_R _16938_ (.A1(_08783_),
    .A2(_09548_),
    .A3(_09605_),
    .B1(_09594_),
    .B2(_05665_),
    .Y(_01485_));
 BUFx4f_ASAP7_75t_R _16939_ (.A(_09600_),
    .Y(_09606_));
 AND2x2_ASAP7_75t_R _16940_ (.A(_09215_),
    .B(_09606_),
    .Y(_09607_));
 INVx1_ASAP7_75t_R _16941_ (.A(_00517_),
    .Y(_09608_));
 AO32x1_ASAP7_75t_R _16942_ (.A1(_09564_),
    .A2(_08805_),
    .A3(_09607_),
    .B1(_09594_),
    .B2(_09608_),
    .Y(_01486_));
 AND3x1_ASAP7_75t_R _16943_ (.A(_09219_),
    .B(_09220_),
    .C(_09601_),
    .Y(_09609_));
 BUFx3_ASAP7_75t_R _16944_ (.A(_09592_),
    .Y(_09610_));
 AO32x1_ASAP7_75t_R _16945_ (.A1(_09564_),
    .A2(_08830_),
    .A3(_09609_),
    .B1(_09610_),
    .B2(_05503_),
    .Y(_01487_));
 BUFx4f_ASAP7_75t_R _16946_ (.A(_09385_),
    .Y(_09611_));
 AND3x1_ASAP7_75t_R _16947_ (.A(_09223_),
    .B(_09224_),
    .C(_09601_),
    .Y(_09612_));
 INVx1_ASAP7_75t_R _16948_ (.A(_00451_),
    .Y(_09613_));
 AO32x1_ASAP7_75t_R _16949_ (.A1(_09611_),
    .A2(_08850_),
    .A3(_09612_),
    .B1(_09610_),
    .B2(_09613_),
    .Y(_01488_));
 NAND2x1_ASAP7_75t_R _16950_ (.A(_01048_),
    .B(_09594_),
    .Y(_09614_));
 OA21x2_ASAP7_75t_R _16951_ (.A1(_09227_),
    .A2(_09593_),
    .B(_09614_),
    .Y(_01489_));
 AND2x2_ASAP7_75t_R _16952_ (.A(_09229_),
    .B(_09606_),
    .Y(_09615_));
 INVx1_ASAP7_75t_R _16953_ (.A(_00418_),
    .Y(_09616_));
 AO32x1_ASAP7_75t_R _16954_ (.A1(_09611_),
    .A2(_08879_),
    .A3(_09615_),
    .B1(_09610_),
    .B2(_09616_),
    .Y(_01490_));
 AND3x1_ASAP7_75t_R _16955_ (.A(_09232_),
    .B(_09233_),
    .C(_09606_),
    .Y(_09617_));
 AO32x1_ASAP7_75t_R _16956_ (.A1(_09611_),
    .A2(_08901_),
    .A3(_09617_),
    .B1(_09610_),
    .B2(_05180_),
    .Y(_01491_));
 AND2x2_ASAP7_75t_R _16957_ (.A(_09236_),
    .B(_09606_),
    .Y(_09618_));
 INVx1_ASAP7_75t_R _16958_ (.A(_00352_),
    .Y(_09619_));
 AO32x1_ASAP7_75t_R _16959_ (.A1(_09611_),
    .A2(_08918_),
    .A3(_09618_),
    .B1(_09610_),
    .B2(_09619_),
    .Y(_01492_));
 AND2x2_ASAP7_75t_R _16960_ (.A(_09240_),
    .B(_09606_),
    .Y(_09620_));
 INVx1_ASAP7_75t_R _16961_ (.A(_00318_),
    .Y(_09621_));
 AO32x1_ASAP7_75t_R _16962_ (.A1(_09611_),
    .A2(_08937_),
    .A3(_09620_),
    .B1(_09610_),
    .B2(_09621_),
    .Y(_01493_));
 AND2x2_ASAP7_75t_R _16963_ (.A(_09243_),
    .B(_09606_),
    .Y(_09622_));
 INVx1_ASAP7_75t_R _16964_ (.A(_00285_),
    .Y(_09623_));
 AO32x1_ASAP7_75t_R _16965_ (.A1(_09611_),
    .A2(_08951_),
    .A3(_09622_),
    .B1(_09610_),
    .B2(_09623_),
    .Y(_01494_));
 AND2x2_ASAP7_75t_R _16966_ (.A(_09246_),
    .B(_09606_),
    .Y(_09624_));
 AO32x1_ASAP7_75t_R _16967_ (.A1(_09611_),
    .A2(_08970_),
    .A3(_09624_),
    .B1(_09610_),
    .B2(_04813_),
    .Y(_01495_));
 NOR2x1_ASAP7_75t_R _16968_ (.A(_08997_),
    .B(_09592_),
    .Y(_09625_));
 INVx1_ASAP7_75t_R _16969_ (.A(_00219_),
    .Y(_09626_));
 AO32x1_ASAP7_75t_R _16970_ (.A1(_09611_),
    .A2(_08987_),
    .A3(_09625_),
    .B1(_09610_),
    .B2(_09626_),
    .Y(_01496_));
 INVx1_ASAP7_75t_R _16971_ (.A(_00185_),
    .Y(_09627_));
 AND2x2_ASAP7_75t_R _16972_ (.A(_09252_),
    .B(_09601_),
    .Y(_09628_));
 AO22x1_ASAP7_75t_R _16973_ (.A1(_09627_),
    .A2(_09594_),
    .B1(_09628_),
    .B2(_09006_),
    .Y(_01497_));
 AND4x1_ASAP7_75t_R _16974_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09606_),
    .Y(_09629_));
 INVx1_ASAP7_75t_R _16975_ (.A(_00152_),
    .Y(_09630_));
 AO32x1_ASAP7_75t_R _16976_ (.A1(_09611_),
    .A2(_09025_),
    .A3(_09629_),
    .B1(_09610_),
    .B2(_09630_),
    .Y(_01498_));
 AND3x1_ASAP7_75t_R _16977_ (.A(_09259_),
    .B(_09260_),
    .C(_09606_),
    .Y(_09631_));
 INVx1_ASAP7_75t_R _16978_ (.A(_00118_),
    .Y(_09632_));
 AO32x1_ASAP7_75t_R _16979_ (.A1(_09611_),
    .A2(_09043_),
    .A3(_09631_),
    .B1(_09592_),
    .B2(_09632_),
    .Y(_01499_));
 NAND2x1_ASAP7_75t_R _16980_ (.A(_01015_),
    .B(_09594_),
    .Y(_09633_));
 OA21x2_ASAP7_75t_R _16981_ (.A1(_09263_),
    .A2(_09593_),
    .B(_09633_),
    .Y(_01500_));
 BUFx3_ASAP7_75t_R _16982_ (.A(_09385_),
    .Y(_09634_));
 AND4x1_ASAP7_75t_R _16983_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09600_),
    .Y(_09635_));
 INVx1_ASAP7_75t_R _16984_ (.A(_00084_),
    .Y(_09636_));
 AO32x1_ASAP7_75t_R _16985_ (.A1(_09634_),
    .A2(_09070_),
    .A3(_09635_),
    .B1(_09592_),
    .B2(_09636_),
    .Y(_01501_));
 AND3x1_ASAP7_75t_R _16986_ (.A(_09270_),
    .B(_09271_),
    .C(_09606_),
    .Y(_09637_));
 INVx1_ASAP7_75t_R _16987_ (.A(_00052_),
    .Y(_09638_));
 AO32x1_ASAP7_75t_R _16988_ (.A1(_09634_),
    .A2(_09086_),
    .A3(_09637_),
    .B1(_09592_),
    .B2(_09638_),
    .Y(_01502_));
 AO21x1_ASAP7_75t_R _16989_ (.A1(_09597_),
    .A2(_09544_),
    .B(_06988_),
    .Y(_09639_));
 OA21x2_ASAP7_75t_R _16990_ (.A1(_09274_),
    .A2(_09593_),
    .B(_09639_),
    .Y(_01503_));
 NAND2x1_ASAP7_75t_R _16991_ (.A(_00949_),
    .B(_09594_),
    .Y(_09640_));
 OA21x2_ASAP7_75t_R _16992_ (.A1(_09276_),
    .A2(_09593_),
    .B(_09640_),
    .Y(_01504_));
 AND2x2_ASAP7_75t_R _16993_ (.A(_00915_),
    .B(_09592_),
    .Y(_09641_));
 AOI21x1_ASAP7_75t_R _16994_ (.A1(_09137_),
    .A2(_09601_),
    .B(_09641_),
    .Y(_01505_));
 AND2x2_ASAP7_75t_R _16995_ (.A(_06709_),
    .B(_09592_),
    .Y(_09642_));
 AO21x1_ASAP7_75t_R _16996_ (.A1(_09279_),
    .A2(_09601_),
    .B(_09642_),
    .Y(_01506_));
 NOR2x1_ASAP7_75t_R _16997_ (.A(_00848_),
    .B(_09601_),
    .Y(_09643_));
 AO21x1_ASAP7_75t_R _16998_ (.A1(_09281_),
    .A2(_09601_),
    .B(_09643_),
    .Y(_01507_));
 AND2x2_ASAP7_75t_R _16999_ (.A(_06484_),
    .B(_09592_),
    .Y(_09644_));
 AO21x1_ASAP7_75t_R _17000_ (.A1(_09283_),
    .A2(_09601_),
    .B(_09644_),
    .Y(_01508_));
 AO21x1_ASAP7_75t_R _17001_ (.A1(_09597_),
    .A2(_09532_),
    .B(_06387_),
    .Y(_09645_));
 OA21x2_ASAP7_75t_R _17002_ (.A1(_09285_),
    .A2(_09594_),
    .B(_09645_),
    .Y(_01509_));
 NAND2x2_ASAP7_75t_R _17003_ (.A(_08602_),
    .B(_09532_),
    .Y(_09646_));
 BUFx10_ASAP7_75t_R _17004_ (.A(_09646_),
    .Y(_09647_));
 BUFx6f_ASAP7_75t_R _17005_ (.A(_09647_),
    .Y(_09648_));
 BUFx12f_ASAP7_75t_R _17006_ (.A(_09646_),
    .Y(_09649_));
 NAND2x1_ASAP7_75t_R _17007_ (.A(_00018_),
    .B(_09649_),
    .Y(_09650_));
 OA21x2_ASAP7_75t_R _17008_ (.A1(_08597_),
    .A2(_09648_),
    .B(_09650_),
    .Y(_01510_));
 NAND2x1_ASAP7_75t_R _17009_ (.A(_00750_),
    .B(_09649_),
    .Y(_09651_));
 OA21x2_ASAP7_75t_R _17010_ (.A1(_09196_),
    .A2(_09648_),
    .B(_09651_),
    .Y(_01511_));
 AO21x1_ASAP7_75t_R _17011_ (.A1(_08871_),
    .A2(_09532_),
    .B(_06220_),
    .Y(_09652_));
 OA21x2_ASAP7_75t_R _17012_ (.A1(_09198_),
    .A2(_09648_),
    .B(_09652_),
    .Y(_01512_));
 AO21x1_ASAP7_75t_R _17013_ (.A1(_08871_),
    .A2(_09532_),
    .B(_06103_),
    .Y(_09653_));
 OA21x2_ASAP7_75t_R _17014_ (.A1(_09200_),
    .A2(_09648_),
    .B(_09653_),
    .Y(_01513_));
 AND2x4_ASAP7_75t_R _17015_ (.A(_08602_),
    .B(_09531_),
    .Y(_09654_));
 BUFx10_ASAP7_75t_R _17016_ (.A(_09654_),
    .Y(_09655_));
 AND2x2_ASAP7_75t_R _17017_ (.A(_00651_),
    .B(_09647_),
    .Y(_09656_));
 AOI21x1_ASAP7_75t_R _17018_ (.A1(_08725_),
    .A2(_09655_),
    .B(_09656_),
    .Y(_01514_));
 NAND2x1_ASAP7_75t_R _17019_ (.A(_00618_),
    .B(_09649_),
    .Y(_09657_));
 OA21x2_ASAP7_75t_R _17020_ (.A1(_09206_),
    .A2(_09648_),
    .B(_09657_),
    .Y(_01515_));
 AO21x1_ASAP7_75t_R _17021_ (.A1(_08871_),
    .A2(_09544_),
    .B(_00584_),
    .Y(_09658_));
 OAI21x1_ASAP7_75t_R _17022_ (.A1(_08766_),
    .A2(_09648_),
    .B(_09658_),
    .Y(_01516_));
 AND3x1_ASAP7_75t_R _17023_ (.A(_09210_),
    .B(_09211_),
    .C(_09655_),
    .Y(_09659_));
 INVx1_ASAP7_75t_R _17024_ (.A(_00551_),
    .Y(_09660_));
 AO32x1_ASAP7_75t_R _17025_ (.A1(_08783_),
    .A2(_09548_),
    .A3(_09659_),
    .B1(_09649_),
    .B2(_09660_),
    .Y(_01517_));
 BUFx3_ASAP7_75t_R _17026_ (.A(_09654_),
    .Y(_09661_));
 AND2x2_ASAP7_75t_R _17027_ (.A(_09215_),
    .B(_09661_),
    .Y(_09662_));
 INVx1_ASAP7_75t_R _17028_ (.A(_00518_),
    .Y(_09663_));
 AO32x1_ASAP7_75t_R _17029_ (.A1(_09634_),
    .A2(_08805_),
    .A3(_09662_),
    .B1(_09649_),
    .B2(_09663_),
    .Y(_01518_));
 AND3x1_ASAP7_75t_R _17030_ (.A(_09219_),
    .B(_09220_),
    .C(_09655_),
    .Y(_09664_));
 BUFx3_ASAP7_75t_R _17031_ (.A(_09647_),
    .Y(_09665_));
 AO32x1_ASAP7_75t_R _17032_ (.A1(_09634_),
    .A2(_08830_),
    .A3(_09664_),
    .B1(_09665_),
    .B2(_05502_),
    .Y(_01519_));
 AND3x1_ASAP7_75t_R _17033_ (.A(_09223_),
    .B(_09224_),
    .C(_09655_),
    .Y(_09666_));
 INVx1_ASAP7_75t_R _17034_ (.A(_00452_),
    .Y(_09667_));
 AO32x1_ASAP7_75t_R _17035_ (.A1(_09634_),
    .A2(_08850_),
    .A3(_09666_),
    .B1(_09665_),
    .B2(_09667_),
    .Y(_01520_));
 NAND2x1_ASAP7_75t_R _17036_ (.A(_01049_),
    .B(_09649_),
    .Y(_09668_));
 OA21x2_ASAP7_75t_R _17037_ (.A1(_09227_),
    .A2(_09648_),
    .B(_09668_),
    .Y(_01521_));
 AND2x2_ASAP7_75t_R _17038_ (.A(_09229_),
    .B(_09661_),
    .Y(_09669_));
 INVx1_ASAP7_75t_R _17039_ (.A(_00419_),
    .Y(_09670_));
 AO32x1_ASAP7_75t_R _17040_ (.A1(_09634_),
    .A2(_08879_),
    .A3(_09669_),
    .B1(_09665_),
    .B2(_09670_),
    .Y(_01522_));
 AND3x1_ASAP7_75t_R _17041_ (.A(_09232_),
    .B(_09233_),
    .C(_09661_),
    .Y(_09671_));
 INVx1_ASAP7_75t_R _17042_ (.A(_00386_),
    .Y(_09672_));
 AO32x1_ASAP7_75t_R _17043_ (.A1(_09634_),
    .A2(_08901_),
    .A3(_09671_),
    .B1(_09665_),
    .B2(_09672_),
    .Y(_01523_));
 AND2x2_ASAP7_75t_R _17044_ (.A(_09236_),
    .B(_09661_),
    .Y(_09673_));
 INVx1_ASAP7_75t_R _17045_ (.A(_00353_),
    .Y(_09674_));
 AO32x1_ASAP7_75t_R _17046_ (.A1(_09634_),
    .A2(_08918_),
    .A3(_09673_),
    .B1(_09665_),
    .B2(_09674_),
    .Y(_01524_));
 AND2x2_ASAP7_75t_R _17047_ (.A(_09240_),
    .B(_09661_),
    .Y(_09675_));
 INVx1_ASAP7_75t_R _17048_ (.A(_00319_),
    .Y(_09676_));
 AO32x1_ASAP7_75t_R _17049_ (.A1(_09634_),
    .A2(_08937_),
    .A3(_09675_),
    .B1(_09665_),
    .B2(_09676_),
    .Y(_01525_));
 AND2x2_ASAP7_75t_R _17050_ (.A(_09243_),
    .B(_09661_),
    .Y(_09677_));
 AO32x1_ASAP7_75t_R _17051_ (.A1(_09634_),
    .A2(_08951_),
    .A3(_09677_),
    .B1(_09665_),
    .B2(_04887_),
    .Y(_01526_));
 BUFx4f_ASAP7_75t_R _17052_ (.A(_09385_),
    .Y(_09678_));
 AND2x2_ASAP7_75t_R _17053_ (.A(_09246_),
    .B(_09661_),
    .Y(_09679_));
 AO32x1_ASAP7_75t_R _17054_ (.A1(_09678_),
    .A2(_08970_),
    .A3(_09679_),
    .B1(_09665_),
    .B2(_04812_),
    .Y(_01527_));
 NOR2x1_ASAP7_75t_R _17055_ (.A(_08997_),
    .B(_09647_),
    .Y(_09680_));
 INVx1_ASAP7_75t_R _17056_ (.A(_00220_),
    .Y(_09681_));
 AO32x1_ASAP7_75t_R _17057_ (.A1(_09678_),
    .A2(_08987_),
    .A3(_09680_),
    .B1(_09665_),
    .B2(_09681_),
    .Y(_01528_));
 INVx1_ASAP7_75t_R _17058_ (.A(_00186_),
    .Y(_09682_));
 AND2x2_ASAP7_75t_R _17059_ (.A(_09252_),
    .B(_09655_),
    .Y(_09683_));
 AO22x1_ASAP7_75t_R _17060_ (.A1(_09682_),
    .A2(_09649_),
    .B1(_09683_),
    .B2(_09006_),
    .Y(_01529_));
 AND4x1_ASAP7_75t_R _17061_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09661_),
    .Y(_09684_));
 INVx1_ASAP7_75t_R _17062_ (.A(_00153_),
    .Y(_09685_));
 AO32x1_ASAP7_75t_R _17063_ (.A1(_09678_),
    .A2(_09025_),
    .A3(_09684_),
    .B1(_09665_),
    .B2(_09685_),
    .Y(_01530_));
 AND3x1_ASAP7_75t_R _17064_ (.A(_09259_),
    .B(_09260_),
    .C(_09661_),
    .Y(_09686_));
 INVx1_ASAP7_75t_R _17065_ (.A(_00119_),
    .Y(_09687_));
 AO32x1_ASAP7_75t_R _17066_ (.A1(_09678_),
    .A2(_09043_),
    .A3(_09686_),
    .B1(_09647_),
    .B2(_09687_),
    .Y(_01531_));
 NAND2x1_ASAP7_75t_R _17067_ (.A(_01016_),
    .B(_09649_),
    .Y(_09688_));
 OA21x2_ASAP7_75t_R _17068_ (.A1(_09263_),
    .A2(_09648_),
    .B(_09688_),
    .Y(_01532_));
 AND4x1_ASAP7_75t_R _17069_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09654_),
    .Y(_09689_));
 INVx1_ASAP7_75t_R _17070_ (.A(_00085_),
    .Y(_09690_));
 AO32x1_ASAP7_75t_R _17071_ (.A1(_09678_),
    .A2(_09070_),
    .A3(_09689_),
    .B1(_09647_),
    .B2(_09690_),
    .Y(_01533_));
 AND3x1_ASAP7_75t_R _17072_ (.A(_09270_),
    .B(_09271_),
    .C(_09661_),
    .Y(_09691_));
 INVx1_ASAP7_75t_R _17073_ (.A(_00053_),
    .Y(_09692_));
 AO32x1_ASAP7_75t_R _17074_ (.A1(_09678_),
    .A2(_09086_),
    .A3(_09691_),
    .B1(_09647_),
    .B2(_09692_),
    .Y(_01534_));
 AO21x1_ASAP7_75t_R _17075_ (.A1(_08871_),
    .A2(_09532_),
    .B(_06987_),
    .Y(_09693_));
 OA21x2_ASAP7_75t_R _17076_ (.A1(_09274_),
    .A2(_09648_),
    .B(_09693_),
    .Y(_01535_));
 NAND2x1_ASAP7_75t_R _17077_ (.A(_00950_),
    .B(_09649_),
    .Y(_09694_));
 OA21x2_ASAP7_75t_R _17078_ (.A1(_09276_),
    .A2(_09648_),
    .B(_09694_),
    .Y(_01536_));
 AND2x2_ASAP7_75t_R _17079_ (.A(_00916_),
    .B(_09647_),
    .Y(_09695_));
 AOI21x1_ASAP7_75t_R _17080_ (.A1(_09137_),
    .A2(_09655_),
    .B(_09695_),
    .Y(_01537_));
 AND2x2_ASAP7_75t_R _17081_ (.A(_06708_),
    .B(_09647_),
    .Y(_09696_));
 AO21x1_ASAP7_75t_R _17082_ (.A1(_09279_),
    .A2(_09655_),
    .B(_09696_),
    .Y(_01538_));
 NOR2x1_ASAP7_75t_R _17083_ (.A(_00849_),
    .B(_09655_),
    .Y(_09697_));
 AO21x1_ASAP7_75t_R _17084_ (.A1(_09281_),
    .A2(_09655_),
    .B(_09697_),
    .Y(_01539_));
 AND2x2_ASAP7_75t_R _17085_ (.A(_06483_),
    .B(_09647_),
    .Y(_09698_));
 AO21x1_ASAP7_75t_R _17086_ (.A1(_09283_),
    .A2(_09655_),
    .B(_09698_),
    .Y(_01540_));
 AO21x1_ASAP7_75t_R _17087_ (.A1(_08871_),
    .A2(_09532_),
    .B(_06386_),
    .Y(_09699_));
 OA21x2_ASAP7_75t_R _17088_ (.A1(_09285_),
    .A2(_09649_),
    .B(_09699_),
    .Y(_01541_));
 NAND2x2_ASAP7_75t_R _17089_ (.A(_09191_),
    .B(_09532_),
    .Y(_09700_));
 BUFx10_ASAP7_75t_R _17090_ (.A(_09700_),
    .Y(_09701_));
 BUFx12_ASAP7_75t_R _17091_ (.A(_09700_),
    .Y(_09702_));
 NAND2x1_ASAP7_75t_R _17092_ (.A(_00019_),
    .B(_09702_),
    .Y(_09703_));
 OA21x2_ASAP7_75t_R _17093_ (.A1(_08597_),
    .A2(_09701_),
    .B(_09703_),
    .Y(_01542_));
 NAND2x1_ASAP7_75t_R _17094_ (.A(_00751_),
    .B(_09702_),
    .Y(_09704_));
 OA21x2_ASAP7_75t_R _17095_ (.A1(_09196_),
    .A2(_09701_),
    .B(_09704_),
    .Y(_01543_));
 NAND2x1_ASAP7_75t_R _17096_ (.A(_00718_),
    .B(_09702_),
    .Y(_09705_));
 OA21x2_ASAP7_75t_R _17097_ (.A1(_09198_),
    .A2(_09701_),
    .B(_09705_),
    .Y(_01544_));
 NAND2x1_ASAP7_75t_R _17098_ (.A(_00685_),
    .B(_09702_),
    .Y(_09706_));
 OA21x2_ASAP7_75t_R _17099_ (.A1(_09200_),
    .A2(_09701_),
    .B(_09706_),
    .Y(_01545_));
 AND2x6_ASAP7_75t_R _17100_ (.A(_09191_),
    .B(_09531_),
    .Y(_09707_));
 BUFx6f_ASAP7_75t_R _17101_ (.A(_09707_),
    .Y(_09708_));
 BUFx6f_ASAP7_75t_R _17102_ (.A(_09700_),
    .Y(_09709_));
 AND2x2_ASAP7_75t_R _17103_ (.A(_00652_),
    .B(_09709_),
    .Y(_09710_));
 AOI21x1_ASAP7_75t_R _17104_ (.A1(_08725_),
    .A2(_09708_),
    .B(_09710_),
    .Y(_01546_));
 NAND2x1_ASAP7_75t_R _17105_ (.A(_00619_),
    .B(_09702_),
    .Y(_09711_));
 OA21x2_ASAP7_75t_R _17106_ (.A1(_09206_),
    .A2(_09701_),
    .B(_09711_),
    .Y(_01547_));
 AO21x1_ASAP7_75t_R _17107_ (.A1(_09191_),
    .A2(_09544_),
    .B(_00585_),
    .Y(_09712_));
 OAI21x1_ASAP7_75t_R _17108_ (.A1(_08766_),
    .A2(_09701_),
    .B(_09712_),
    .Y(_01548_));
 AND3x1_ASAP7_75t_R _17109_ (.A(_09210_),
    .B(_09211_),
    .C(_09708_),
    .Y(_09713_));
 BUFx12_ASAP7_75t_R _17110_ (.A(_09700_),
    .Y(_09714_));
 AO32x1_ASAP7_75t_R _17111_ (.A1(_08783_),
    .A2(_09548_),
    .A3(_09713_),
    .B1(_09714_),
    .B2(_05663_),
    .Y(_01549_));
 BUFx3_ASAP7_75t_R _17112_ (.A(_09707_),
    .Y(_09715_));
 AND2x2_ASAP7_75t_R _17113_ (.A(_09215_),
    .B(_09715_),
    .Y(_09716_));
 INVx1_ASAP7_75t_R _17114_ (.A(_00519_),
    .Y(_09717_));
 AO32x1_ASAP7_75t_R _17115_ (.A1(_09678_),
    .A2(_08805_),
    .A3(_09716_),
    .B1(_09714_),
    .B2(_09717_),
    .Y(_01550_));
 AND3x1_ASAP7_75t_R _17116_ (.A(_09219_),
    .B(_09220_),
    .C(_09715_),
    .Y(_09718_));
 INVx1_ASAP7_75t_R _17117_ (.A(_00486_),
    .Y(_09719_));
 AO32x1_ASAP7_75t_R _17118_ (.A1(_09678_),
    .A2(_08830_),
    .A3(_09718_),
    .B1(_09714_),
    .B2(_09719_),
    .Y(_01551_));
 AND3x1_ASAP7_75t_R _17119_ (.A(_09223_),
    .B(_09224_),
    .C(_09715_),
    .Y(_09720_));
 INVx1_ASAP7_75t_R _17120_ (.A(_00453_),
    .Y(_09721_));
 AO32x1_ASAP7_75t_R _17121_ (.A1(_09678_),
    .A2(_08850_),
    .A3(_09720_),
    .B1(_09714_),
    .B2(_09721_),
    .Y(_01552_));
 NAND2x1_ASAP7_75t_R _17122_ (.A(_01050_),
    .B(_09702_),
    .Y(_09722_));
 OA21x2_ASAP7_75t_R _17123_ (.A1(_09227_),
    .A2(_09701_),
    .B(_09722_),
    .Y(_01553_));
 AND2x2_ASAP7_75t_R _17124_ (.A(_09229_),
    .B(_09715_),
    .Y(_09723_));
 INVx1_ASAP7_75t_R _17125_ (.A(_00420_),
    .Y(_09724_));
 AO32x1_ASAP7_75t_R _17126_ (.A1(_09678_),
    .A2(_08879_),
    .A3(_09723_),
    .B1(_09714_),
    .B2(_09724_),
    .Y(_01554_));
 BUFx3_ASAP7_75t_R _17127_ (.A(_09385_),
    .Y(_09725_));
 AND3x1_ASAP7_75t_R _17128_ (.A(_09232_),
    .B(_09233_),
    .C(_09715_),
    .Y(_09726_));
 AO32x1_ASAP7_75t_R _17129_ (.A1(_09725_),
    .A2(_08901_),
    .A3(_09726_),
    .B1(_09714_),
    .B2(_05178_),
    .Y(_01555_));
 AND2x2_ASAP7_75t_R _17130_ (.A(_09236_),
    .B(_09715_),
    .Y(_09727_));
 INVx1_ASAP7_75t_R _17131_ (.A(_00354_),
    .Y(_09728_));
 AO32x1_ASAP7_75t_R _17132_ (.A1(_09725_),
    .A2(_08918_),
    .A3(_09727_),
    .B1(_09714_),
    .B2(_09728_),
    .Y(_01556_));
 AND2x2_ASAP7_75t_R _17133_ (.A(_09240_),
    .B(_09715_),
    .Y(_09729_));
 INVx1_ASAP7_75t_R _17134_ (.A(_00320_),
    .Y(_09730_));
 AO32x1_ASAP7_75t_R _17135_ (.A1(_09725_),
    .A2(_08937_),
    .A3(_09729_),
    .B1(_09714_),
    .B2(_09730_),
    .Y(_01557_));
 AND2x2_ASAP7_75t_R _17136_ (.A(_09243_),
    .B(_09715_),
    .Y(_09731_));
 INVx1_ASAP7_75t_R _17137_ (.A(_00287_),
    .Y(_09732_));
 AO32x1_ASAP7_75t_R _17138_ (.A1(_09725_),
    .A2(_08951_),
    .A3(_09731_),
    .B1(_09709_),
    .B2(_09732_),
    .Y(_01558_));
 AND2x2_ASAP7_75t_R _17139_ (.A(_09246_),
    .B(_09707_),
    .Y(_09733_));
 INVx1_ASAP7_75t_R _17140_ (.A(_00254_),
    .Y(_09734_));
 AO32x1_ASAP7_75t_R _17141_ (.A1(_09725_),
    .A2(_08970_),
    .A3(_09733_),
    .B1(_09709_),
    .B2(_09734_),
    .Y(_01559_));
 NOR2x1_ASAP7_75t_R _17142_ (.A(_08997_),
    .B(_09709_),
    .Y(_09735_));
 INVx1_ASAP7_75t_R _17143_ (.A(_00221_),
    .Y(_09736_));
 AO32x1_ASAP7_75t_R _17144_ (.A1(_09725_),
    .A2(_08987_),
    .A3(_09735_),
    .B1(_09709_),
    .B2(_09736_),
    .Y(_01560_));
 INVx1_ASAP7_75t_R _17145_ (.A(_00187_),
    .Y(_09737_));
 AND2x2_ASAP7_75t_R _17146_ (.A(_09252_),
    .B(_09708_),
    .Y(_09738_));
 AO22x1_ASAP7_75t_R _17147_ (.A1(_09737_),
    .A2(_09702_),
    .B1(_09738_),
    .B2(_09006_),
    .Y(_01561_));
 AND4x1_ASAP7_75t_R _17148_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09707_),
    .Y(_09739_));
 INVx1_ASAP7_75t_R _17149_ (.A(_00154_),
    .Y(_09740_));
 AO32x1_ASAP7_75t_R _17150_ (.A1(_09725_),
    .A2(_09025_),
    .A3(_09739_),
    .B1(_09709_),
    .B2(_09740_),
    .Y(_01562_));
 AND3x1_ASAP7_75t_R _17151_ (.A(_09259_),
    .B(_09260_),
    .C(_09715_),
    .Y(_09741_));
 INVx1_ASAP7_75t_R _17152_ (.A(_00120_),
    .Y(_09742_));
 AO32x1_ASAP7_75t_R _17153_ (.A1(_09725_),
    .A2(_09043_),
    .A3(_09741_),
    .B1(_09709_),
    .B2(_09742_),
    .Y(_01563_));
 NAND2x1_ASAP7_75t_R _17154_ (.A(_01017_),
    .B(_09702_),
    .Y(_09743_));
 OA21x2_ASAP7_75t_R _17155_ (.A1(_09263_),
    .A2(_09701_),
    .B(_09743_),
    .Y(_01564_));
 AND4x1_ASAP7_75t_R _17156_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09707_),
    .Y(_09744_));
 INVx1_ASAP7_75t_R _17157_ (.A(_00086_),
    .Y(_09745_));
 AO32x1_ASAP7_75t_R _17158_ (.A1(_09725_),
    .A2(_09070_),
    .A3(_09744_),
    .B1(_09709_),
    .B2(_09745_),
    .Y(_01565_));
 AND3x1_ASAP7_75t_R _17159_ (.A(_09270_),
    .B(_09271_),
    .C(_09715_),
    .Y(_09746_));
 INVx1_ASAP7_75t_R _17160_ (.A(_00054_),
    .Y(_09747_));
 AO32x1_ASAP7_75t_R _17161_ (.A1(_09725_),
    .A2(_09086_),
    .A3(_09746_),
    .B1(_09709_),
    .B2(_09747_),
    .Y(_01566_));
 NAND2x1_ASAP7_75t_R _17162_ (.A(_00984_),
    .B(_09702_),
    .Y(_09748_));
 OA21x2_ASAP7_75t_R _17163_ (.A1(_09274_),
    .A2(_09701_),
    .B(_09748_),
    .Y(_01567_));
 NAND2x1_ASAP7_75t_R _17164_ (.A(_00951_),
    .B(_09714_),
    .Y(_09749_));
 OA21x2_ASAP7_75t_R _17165_ (.A1(_09276_),
    .A2(_09701_),
    .B(_09749_),
    .Y(_01568_));
 AND2x2_ASAP7_75t_R _17166_ (.A(_00917_),
    .B(_09709_),
    .Y(_09750_));
 AOI21x1_ASAP7_75t_R _17167_ (.A1(_09137_),
    .A2(_09708_),
    .B(_09750_),
    .Y(_01569_));
 NOR2x1_ASAP7_75t_R _17168_ (.A(_00884_),
    .B(_09708_),
    .Y(_09751_));
 AO21x1_ASAP7_75t_R _17169_ (.A1(_09279_),
    .A2(_09708_),
    .B(_09751_),
    .Y(_01570_));
 NOR2x1_ASAP7_75t_R _17170_ (.A(_00850_),
    .B(_09708_),
    .Y(_09752_));
 AO21x1_ASAP7_75t_R _17171_ (.A1(_09281_),
    .A2(_09708_),
    .B(_09752_),
    .Y(_01571_));
 NOR2x1_ASAP7_75t_R _17172_ (.A(_00817_),
    .B(_09708_),
    .Y(_09753_));
 AO21x1_ASAP7_75t_R _17173_ (.A1(_09283_),
    .A2(_09708_),
    .B(_09753_),
    .Y(_01572_));
 NAND2x1_ASAP7_75t_R _17174_ (.A(_00783_),
    .B(_09714_),
    .Y(_09754_));
 OA21x2_ASAP7_75t_R _17175_ (.A1(_09285_),
    .A2(_09702_),
    .B(_09754_),
    .Y(_01573_));
 BUFx6f_ASAP7_75t_R _17176_ (.A(_08596_),
    .Y(_09755_));
 OR3x4_ASAP7_75t_R _17177_ (.A(_07131_),
    .B(_09349_),
    .C(_09526_),
    .Y(_09756_));
 BUFx10_ASAP7_75t_R _17178_ (.A(_09756_),
    .Y(_09757_));
 BUFx12f_ASAP7_75t_R _17179_ (.A(_09756_),
    .Y(_09758_));
 NAND2x1_ASAP7_75t_R _17180_ (.A(_00001_),
    .B(_09758_),
    .Y(_09759_));
 OA21x2_ASAP7_75t_R _17181_ (.A1(_09755_),
    .A2(_09757_),
    .B(_09759_),
    .Y(_01574_));
 NAND2x1_ASAP7_75t_R _17182_ (.A(_00733_),
    .B(_09758_),
    .Y(_09760_));
 OA21x2_ASAP7_75t_R _17183_ (.A1(_09196_),
    .A2(_09757_),
    .B(_09760_),
    .Y(_01575_));
 NAND2x1_ASAP7_75t_R _17184_ (.A(_00700_),
    .B(_09758_),
    .Y(_09761_));
 OA21x2_ASAP7_75t_R _17185_ (.A1(_09198_),
    .A2(_09757_),
    .B(_09761_),
    .Y(_01576_));
 NAND2x1_ASAP7_75t_R _17186_ (.A(_00667_),
    .B(_09758_),
    .Y(_09762_));
 OA21x2_ASAP7_75t_R _17187_ (.A1(_09200_),
    .A2(_09757_),
    .B(_09762_),
    .Y(_01577_));
 BUFx10_ASAP7_75t_R _17188_ (.A(_08724_),
    .Y(_09763_));
 AND2x6_ASAP7_75t_R _17189_ (.A(_09288_),
    .B(_09589_),
    .Y(_09764_));
 BUFx6f_ASAP7_75t_R _17190_ (.A(_09764_),
    .Y(_09765_));
 BUFx10_ASAP7_75t_R _17191_ (.A(_09756_),
    .Y(_09766_));
 AND2x2_ASAP7_75t_R _17192_ (.A(_00634_),
    .B(_09766_),
    .Y(_09767_));
 AOI21x1_ASAP7_75t_R _17193_ (.A1(_09763_),
    .A2(_09765_),
    .B(_09767_),
    .Y(_01578_));
 NAND2x1_ASAP7_75t_R _17194_ (.A(_00601_),
    .B(_09758_),
    .Y(_09768_));
 OA21x2_ASAP7_75t_R _17195_ (.A1(_09206_),
    .A2(_09757_),
    .B(_09768_),
    .Y(_01579_));
 BUFx12f_ASAP7_75t_R _17196_ (.A(_08765_),
    .Y(_09769_));
 AND2x2_ASAP7_75t_R _17197_ (.A(_00567_),
    .B(_09766_),
    .Y(_09770_));
 AOI21x1_ASAP7_75t_R _17198_ (.A1(_09769_),
    .A2(_09765_),
    .B(_09770_),
    .Y(_01580_));
 BUFx4f_ASAP7_75t_R _17199_ (.A(_08782_),
    .Y(_09771_));
 BUFx4f_ASAP7_75t_R _17200_ (.A(_09764_),
    .Y(_09772_));
 AND3x2_ASAP7_75t_R _17201_ (.A(_09210_),
    .B(_09211_),
    .C(_09772_),
    .Y(_09773_));
 BUFx6f_ASAP7_75t_R _17202_ (.A(_09756_),
    .Y(_09774_));
 AO32x1_ASAP7_75t_R _17203_ (.A1(_09771_),
    .A2(_09548_),
    .A3(_09773_),
    .B1(_09774_),
    .B2(_05709_),
    .Y(_01581_));
 BUFx4f_ASAP7_75t_R _17204_ (.A(_09385_),
    .Y(_09775_));
 BUFx4f_ASAP7_75t_R _17205_ (.A(_08804_),
    .Y(_09776_));
 AND2x2_ASAP7_75t_R _17206_ (.A(_09215_),
    .B(_09772_),
    .Y(_09777_));
 INVx1_ASAP7_75t_R _17207_ (.A(_00501_),
    .Y(_09778_));
 AO32x1_ASAP7_75t_R _17208_ (.A1(_09775_),
    .A2(_09776_),
    .A3(_09777_),
    .B1(_09774_),
    .B2(_09778_),
    .Y(_01582_));
 BUFx4f_ASAP7_75t_R _17209_ (.A(_08829_),
    .Y(_09779_));
 AND3x1_ASAP7_75t_R _17210_ (.A(_09219_),
    .B(_09220_),
    .C(_09772_),
    .Y(_09780_));
 INVx1_ASAP7_75t_R _17211_ (.A(_00468_),
    .Y(_09781_));
 AO32x1_ASAP7_75t_R _17212_ (.A1(_09775_),
    .A2(_09779_),
    .A3(_09780_),
    .B1(_09774_),
    .B2(_09781_),
    .Y(_01583_));
 BUFx4f_ASAP7_75t_R _17213_ (.A(_08849_),
    .Y(_09782_));
 AND3x1_ASAP7_75t_R _17214_ (.A(_09223_),
    .B(_09224_),
    .C(_09772_),
    .Y(_09783_));
 INVx1_ASAP7_75t_R _17215_ (.A(_00435_),
    .Y(_09784_));
 AO32x1_ASAP7_75t_R _17216_ (.A1(_09775_),
    .A2(_09782_),
    .A3(_09783_),
    .B1(_09774_),
    .B2(_09784_),
    .Y(_01584_));
 NAND2x1_ASAP7_75t_R _17217_ (.A(_01032_),
    .B(_09758_),
    .Y(_09785_));
 OA21x2_ASAP7_75t_R _17218_ (.A1(_09227_),
    .A2(_09757_),
    .B(_09785_),
    .Y(_01585_));
 BUFx4f_ASAP7_75t_R _17219_ (.A(_08878_),
    .Y(_09786_));
 AND2x2_ASAP7_75t_R _17220_ (.A(_09229_),
    .B(_09772_),
    .Y(_09787_));
 INVx1_ASAP7_75t_R _17221_ (.A(_00402_),
    .Y(_09788_));
 AO32x1_ASAP7_75t_R _17222_ (.A1(_09775_),
    .A2(_09786_),
    .A3(_09787_),
    .B1(_09774_),
    .B2(_09788_),
    .Y(_01586_));
 BUFx4f_ASAP7_75t_R _17223_ (.A(_08900_),
    .Y(_09789_));
 AND3x1_ASAP7_75t_R _17224_ (.A(_09232_),
    .B(_09233_),
    .C(_09772_),
    .Y(_09790_));
 INVx1_ASAP7_75t_R _17225_ (.A(_00369_),
    .Y(_09791_));
 AO32x1_ASAP7_75t_R _17226_ (.A1(_09775_),
    .A2(_09789_),
    .A3(_09790_),
    .B1(_09774_),
    .B2(_09791_),
    .Y(_01587_));
 BUFx3_ASAP7_75t_R _17227_ (.A(_08917_),
    .Y(_09792_));
 AND2x2_ASAP7_75t_R _17228_ (.A(_09236_),
    .B(_09772_),
    .Y(_09793_));
 AO32x1_ASAP7_75t_R _17229_ (.A1(_09775_),
    .A2(_09792_),
    .A3(_09793_),
    .B1(_09774_),
    .B2(_05149_),
    .Y(_01588_));
 BUFx3_ASAP7_75t_R _17230_ (.A(_08936_),
    .Y(_09794_));
 AND2x2_ASAP7_75t_R _17231_ (.A(_09240_),
    .B(_09772_),
    .Y(_09795_));
 INVx1_ASAP7_75t_R _17232_ (.A(_00302_),
    .Y(_09796_));
 AO32x1_ASAP7_75t_R _17233_ (.A1(_09775_),
    .A2(_09794_),
    .A3(_09795_),
    .B1(_09774_),
    .B2(_09796_),
    .Y(_01589_));
 BUFx4f_ASAP7_75t_R _17234_ (.A(_08950_),
    .Y(_09797_));
 AND2x2_ASAP7_75t_R _17235_ (.A(_09243_),
    .B(_09764_),
    .Y(_09798_));
 INVx1_ASAP7_75t_R _17236_ (.A(_00269_),
    .Y(_09799_));
 AO32x1_ASAP7_75t_R _17237_ (.A1(_09775_),
    .A2(_09797_),
    .A3(_09798_),
    .B1(_09774_),
    .B2(_09799_),
    .Y(_01590_));
 BUFx6f_ASAP7_75t_R _17238_ (.A(_08969_),
    .Y(_09800_));
 AND2x2_ASAP7_75t_R _17239_ (.A(_09246_),
    .B(_09764_),
    .Y(_09801_));
 INVx1_ASAP7_75t_R _17240_ (.A(_00236_),
    .Y(_09802_));
 AO32x1_ASAP7_75t_R _17241_ (.A1(_09775_),
    .A2(_09800_),
    .A3(_09801_),
    .B1(_09766_),
    .B2(_09802_),
    .Y(_01591_));
 BUFx4f_ASAP7_75t_R _17242_ (.A(_08986_),
    .Y(_09803_));
 BUFx10_ASAP7_75t_R _17243_ (.A(_08996_),
    .Y(_09804_));
 NOR2x1_ASAP7_75t_R _17244_ (.A(_09804_),
    .B(_09766_),
    .Y(_09805_));
 AO32x1_ASAP7_75t_R _17245_ (.A1(_09775_),
    .A2(_09803_),
    .A3(_09805_),
    .B1(_09766_),
    .B2(_04732_),
    .Y(_01592_));
 INVx1_ASAP7_75t_R _17246_ (.A(_00169_),
    .Y(_09806_));
 AND2x2_ASAP7_75t_R _17247_ (.A(_09252_),
    .B(_09765_),
    .Y(_09807_));
 BUFx3_ASAP7_75t_R _17248_ (.A(_09005_),
    .Y(_09808_));
 AO22x1_ASAP7_75t_R _17249_ (.A1(_09806_),
    .A2(_09758_),
    .B1(_09807_),
    .B2(_09808_),
    .Y(_01593_));
 BUFx6f_ASAP7_75t_R _17250_ (.A(_08784_),
    .Y(_09809_));
 BUFx6f_ASAP7_75t_R _17251_ (.A(_09809_),
    .Y(_09810_));
 BUFx4f_ASAP7_75t_R _17252_ (.A(_09024_),
    .Y(_09811_));
 AND4x1_ASAP7_75t_R _17253_ (.A(_09254_),
    .B(_09255_),
    .C(_09256_),
    .D(_09764_),
    .Y(_09812_));
 AO32x1_ASAP7_75t_R _17254_ (.A1(_09810_),
    .A2(_09811_),
    .A3(_09812_),
    .B1(_09766_),
    .B2(_04443_),
    .Y(_01594_));
 BUFx4f_ASAP7_75t_R _17255_ (.A(_09042_),
    .Y(_09813_));
 AND3x1_ASAP7_75t_R _17256_ (.A(_09259_),
    .B(_09260_),
    .C(_09772_),
    .Y(_09814_));
 AO32x1_ASAP7_75t_R _17257_ (.A1(_09810_),
    .A2(_09813_),
    .A3(_09814_),
    .B1(_09766_),
    .B2(_04368_),
    .Y(_01595_));
 NAND2x1_ASAP7_75t_R _17258_ (.A(_00999_),
    .B(_09758_),
    .Y(_09815_));
 OA21x2_ASAP7_75t_R _17259_ (.A1(_09263_),
    .A2(_09757_),
    .B(_09815_),
    .Y(_01596_));
 BUFx4f_ASAP7_75t_R _17260_ (.A(_09069_),
    .Y(_09816_));
 AND4x1_ASAP7_75t_R _17261_ (.A(_09265_),
    .B(_09266_),
    .C(_09267_),
    .D(_09764_),
    .Y(_09817_));
 AO32x1_ASAP7_75t_R _17262_ (.A1(_09810_),
    .A2(_09816_),
    .A3(_09817_),
    .B1(_09766_),
    .B2(_04186_),
    .Y(_01597_));
 BUFx4f_ASAP7_75t_R _17263_ (.A(_09085_),
    .Y(_09818_));
 AND3x1_ASAP7_75t_R _17264_ (.A(_09270_),
    .B(_09271_),
    .C(_09772_),
    .Y(_09819_));
 AO32x1_ASAP7_75t_R _17265_ (.A1(_09810_),
    .A2(_09818_),
    .A3(_09819_),
    .B1(_09766_),
    .B2(_03903_),
    .Y(_01598_));
 NAND2x1_ASAP7_75t_R _17266_ (.A(_00966_),
    .B(_09758_),
    .Y(_09820_));
 OA21x2_ASAP7_75t_R _17267_ (.A1(_09274_),
    .A2(_09757_),
    .B(_09820_),
    .Y(_01599_));
 NAND2x1_ASAP7_75t_R _17268_ (.A(_00933_),
    .B(_09758_),
    .Y(_09821_));
 OA21x2_ASAP7_75t_R _17269_ (.A1(_09276_),
    .A2(_09757_),
    .B(_09821_),
    .Y(_01600_));
 BUFx6f_ASAP7_75t_R _17270_ (.A(_09136_),
    .Y(_09822_));
 AND2x2_ASAP7_75t_R _17271_ (.A(_00899_),
    .B(_09766_),
    .Y(_09823_));
 AOI21x1_ASAP7_75t_R _17272_ (.A1(_09822_),
    .A2(_09765_),
    .B(_09823_),
    .Y(_01601_));
 NOR2x1_ASAP7_75t_R _17273_ (.A(_00866_),
    .B(_09765_),
    .Y(_09824_));
 AO21x1_ASAP7_75t_R _17274_ (.A1(_09279_),
    .A2(_09765_),
    .B(_09824_),
    .Y(_01602_));
 NOR2x1_ASAP7_75t_R _17275_ (.A(_00832_),
    .B(_09765_),
    .Y(_09825_));
 AO21x1_ASAP7_75t_R _17276_ (.A1(_09281_),
    .A2(_09765_),
    .B(_09825_),
    .Y(_01603_));
 NOR2x1_ASAP7_75t_R _17277_ (.A(_00799_),
    .B(_09765_),
    .Y(_09826_));
 AO21x1_ASAP7_75t_R _17278_ (.A1(_09283_),
    .A2(_09765_),
    .B(_09826_),
    .Y(_01604_));
 NAND2x1_ASAP7_75t_R _17279_ (.A(_00765_),
    .B(_09774_),
    .Y(_09827_));
 OA21x2_ASAP7_75t_R _17280_ (.A1(_09285_),
    .A2(_09757_),
    .B(_09827_),
    .Y(_01605_));
 INVx1_ASAP7_75t_R _17281_ (.A(net3),
    .Y(_09828_));
 OR4x1_ASAP7_75t_R _17282_ (.A(_04072_),
    .B(_09828_),
    .C(net2),
    .D(_09530_),
    .Y(_09829_));
 BUFx10_ASAP7_75t_R _17283_ (.A(_09829_),
    .Y(_09830_));
 OR2x6_ASAP7_75t_R _17284_ (.A(_09289_),
    .B(_09830_),
    .Y(_09831_));
 BUFx4f_ASAP7_75t_R _17285_ (.A(_09831_),
    .Y(_09832_));
 BUFx6f_ASAP7_75t_R _17286_ (.A(_09831_),
    .Y(_09833_));
 NAND2x1_ASAP7_75t_R _17287_ (.A(_00020_),
    .B(_09833_),
    .Y(_09834_));
 OA21x2_ASAP7_75t_R _17288_ (.A1(_09755_),
    .A2(_09832_),
    .B(_09834_),
    .Y(_01606_));
 BUFx4f_ASAP7_75t_R _17289_ (.A(_08654_),
    .Y(_09835_));
 NAND2x1_ASAP7_75t_R _17290_ (.A(_00752_),
    .B(_09833_),
    .Y(_09836_));
 OA21x2_ASAP7_75t_R _17291_ (.A1(_09835_),
    .A2(_09832_),
    .B(_09836_),
    .Y(_01607_));
 BUFx4f_ASAP7_75t_R _17292_ (.A(_08681_),
    .Y(_09837_));
 NAND2x1_ASAP7_75t_R _17293_ (.A(_00719_),
    .B(_09833_),
    .Y(_09838_));
 OA21x2_ASAP7_75t_R _17294_ (.A1(_09837_),
    .A2(_09832_),
    .B(_09838_),
    .Y(_01608_));
 BUFx4f_ASAP7_75t_R _17295_ (.A(_08697_),
    .Y(_09839_));
 NAND2x1_ASAP7_75t_R _17296_ (.A(_00686_),
    .B(_09833_),
    .Y(_09840_));
 OA21x2_ASAP7_75t_R _17297_ (.A1(_09839_),
    .A2(_09832_),
    .B(_09840_),
    .Y(_01609_));
 NOR2x2_ASAP7_75t_R _17298_ (.A(_09289_),
    .B(_09830_),
    .Y(_09841_));
 BUFx6f_ASAP7_75t_R _17299_ (.A(_09841_),
    .Y(_09842_));
 BUFx6f_ASAP7_75t_R _17300_ (.A(_09831_),
    .Y(_09843_));
 AND2x2_ASAP7_75t_R _17301_ (.A(_00653_),
    .B(_09843_),
    .Y(_09844_));
 AOI21x1_ASAP7_75t_R _17302_ (.A1(_09763_),
    .A2(_09842_),
    .B(_09844_),
    .Y(_01610_));
 BUFx4f_ASAP7_75t_R _17303_ (.A(_08744_),
    .Y(_09845_));
 NAND2x1_ASAP7_75t_R _17304_ (.A(_00620_),
    .B(_09833_),
    .Y(_09846_));
 OA21x2_ASAP7_75t_R _17305_ (.A1(_09845_),
    .A2(_09832_),
    .B(_09846_),
    .Y(_01611_));
 AND2x2_ASAP7_75t_R _17306_ (.A(_00586_),
    .B(_09843_),
    .Y(_09847_));
 AOI21x1_ASAP7_75t_R _17307_ (.A1(_09769_),
    .A2(_09842_),
    .B(_09847_),
    .Y(_01612_));
 BUFx4f_ASAP7_75t_R _17308_ (.A(_08786_),
    .Y(_09848_));
 BUFx3_ASAP7_75t_R _17309_ (.A(_08794_),
    .Y(_09849_));
 BUFx4f_ASAP7_75t_R _17310_ (.A(_09841_),
    .Y(_09850_));
 AND3x1_ASAP7_75t_R _17311_ (.A(_09848_),
    .B(_09849_),
    .C(_09850_),
    .Y(_09851_));
 BUFx6f_ASAP7_75t_R _17312_ (.A(_09831_),
    .Y(_09852_));
 INVx1_ASAP7_75t_R _17313_ (.A(_00553_),
    .Y(_09853_));
 AO32x1_ASAP7_75t_R _17314_ (.A1(_09771_),
    .A2(_09548_),
    .A3(_09851_),
    .B1(_09852_),
    .B2(_09853_),
    .Y(_01613_));
 BUFx4f_ASAP7_75t_R _17315_ (.A(_08821_),
    .Y(_09854_));
 AND2x2_ASAP7_75t_R _17316_ (.A(_09854_),
    .B(_09850_),
    .Y(_09855_));
 INVx1_ASAP7_75t_R _17317_ (.A(_00520_),
    .Y(_09856_));
 AO32x1_ASAP7_75t_R _17318_ (.A1(_09810_),
    .A2(_09776_),
    .A3(_09855_),
    .B1(_09852_),
    .B2(_09856_),
    .Y(_01614_));
 BUFx6f_ASAP7_75t_R _17319_ (.A(_08834_),
    .Y(_09857_));
 BUFx4f_ASAP7_75t_R _17320_ (.A(_08841_),
    .Y(_09858_));
 AND3x1_ASAP7_75t_R _17321_ (.A(_09857_),
    .B(_09858_),
    .C(_09850_),
    .Y(_09859_));
 INVx1_ASAP7_75t_R _17322_ (.A(_00487_),
    .Y(_09860_));
 AO32x1_ASAP7_75t_R _17323_ (.A1(_09810_),
    .A2(_09779_),
    .A3(_09859_),
    .B1(_09852_),
    .B2(_09860_),
    .Y(_01615_));
 BUFx4f_ASAP7_75t_R _17324_ (.A(_08851_),
    .Y(_09861_));
 BUFx4f_ASAP7_75t_R _17325_ (.A(_08860_),
    .Y(_09862_));
 AND3x1_ASAP7_75t_R _17326_ (.A(_09861_),
    .B(_09862_),
    .C(_09850_),
    .Y(_09863_));
 INVx1_ASAP7_75t_R _17327_ (.A(_00454_),
    .Y(_09864_));
 AO32x1_ASAP7_75t_R _17328_ (.A1(_09810_),
    .A2(_09782_),
    .A3(_09863_),
    .B1(_09852_),
    .B2(_09864_),
    .Y(_01616_));
 BUFx4f_ASAP7_75t_R _17329_ (.A(_08870_),
    .Y(_09865_));
 NAND2x1_ASAP7_75t_R _17330_ (.A(_01051_),
    .B(_09833_),
    .Y(_09866_));
 OA21x2_ASAP7_75t_R _17331_ (.A1(_09865_),
    .A2(_09832_),
    .B(_09866_),
    .Y(_01617_));
 BUFx4f_ASAP7_75t_R _17332_ (.A(_08892_),
    .Y(_09867_));
 AND2x2_ASAP7_75t_R _17333_ (.A(_09867_),
    .B(_09850_),
    .Y(_09868_));
 INVx1_ASAP7_75t_R _17334_ (.A(_00421_),
    .Y(_09869_));
 AO32x1_ASAP7_75t_R _17335_ (.A1(_09810_),
    .A2(_09786_),
    .A3(_09868_),
    .B1(_09852_),
    .B2(_09869_),
    .Y(_01618_));
 BUFx4f_ASAP7_75t_R _17336_ (.A(_08902_),
    .Y(_09870_));
 BUFx4f_ASAP7_75t_R _17337_ (.A(_08910_),
    .Y(_09871_));
 AND3x1_ASAP7_75t_R _17338_ (.A(_09870_),
    .B(_09871_),
    .C(_09850_),
    .Y(_09872_));
 INVx1_ASAP7_75t_R _17339_ (.A(_00388_),
    .Y(_09873_));
 AO32x1_ASAP7_75t_R _17340_ (.A1(_09810_),
    .A2(_09789_),
    .A3(_09872_),
    .B1(_09852_),
    .B2(_09873_),
    .Y(_01619_));
 BUFx3_ASAP7_75t_R _17341_ (.A(_08929_),
    .Y(_09874_));
 AND2x2_ASAP7_75t_R _17342_ (.A(_09874_),
    .B(_09850_),
    .Y(_09875_));
 INVx1_ASAP7_75t_R _17343_ (.A(_00355_),
    .Y(_09876_));
 AO32x1_ASAP7_75t_R _17344_ (.A1(_09810_),
    .A2(_09792_),
    .A3(_09875_),
    .B1(_09852_),
    .B2(_09876_),
    .Y(_01620_));
 BUFx4f_ASAP7_75t_R _17345_ (.A(_09809_),
    .Y(_09877_));
 BUFx3_ASAP7_75t_R _17346_ (.A(_08943_),
    .Y(_09878_));
 AND2x2_ASAP7_75t_R _17347_ (.A(_09878_),
    .B(_09850_),
    .Y(_09879_));
 INVx1_ASAP7_75t_R _17348_ (.A(_00321_),
    .Y(_09880_));
 AO32x1_ASAP7_75t_R _17349_ (.A1(_09877_),
    .A2(_09794_),
    .A3(_09879_),
    .B1(_09852_),
    .B2(_09880_),
    .Y(_01621_));
 BUFx4f_ASAP7_75t_R _17350_ (.A(_08962_),
    .Y(_09881_));
 AND2x2_ASAP7_75t_R _17351_ (.A(_09881_),
    .B(_09841_),
    .Y(_09882_));
 INVx1_ASAP7_75t_R _17352_ (.A(_00288_),
    .Y(_09883_));
 AO32x1_ASAP7_75t_R _17353_ (.A1(_09877_),
    .A2(_09797_),
    .A3(_09882_),
    .B1(_09852_),
    .B2(_09883_),
    .Y(_01622_));
 BUFx6f_ASAP7_75t_R _17354_ (.A(_08979_),
    .Y(_09884_));
 AND2x2_ASAP7_75t_R _17355_ (.A(_09884_),
    .B(_09841_),
    .Y(_09885_));
 INVx1_ASAP7_75t_R _17356_ (.A(_00255_),
    .Y(_09886_));
 AO32x1_ASAP7_75t_R _17357_ (.A1(_09877_),
    .A2(_09800_),
    .A3(_09885_),
    .B1(_09843_),
    .B2(_09886_),
    .Y(_01623_));
 NOR2x1_ASAP7_75t_R _17358_ (.A(_09804_),
    .B(_09843_),
    .Y(_09887_));
 INVx1_ASAP7_75t_R _17359_ (.A(_00222_),
    .Y(_09888_));
 AO32x1_ASAP7_75t_R _17360_ (.A1(_09877_),
    .A2(_09803_),
    .A3(_09887_),
    .B1(_09843_),
    .B2(_09888_),
    .Y(_01624_));
 INVx1_ASAP7_75t_R _17361_ (.A(_00188_),
    .Y(_09889_));
 BUFx3_ASAP7_75t_R _17362_ (.A(_09017_),
    .Y(_09890_));
 AND2x2_ASAP7_75t_R _17363_ (.A(_09890_),
    .B(_09842_),
    .Y(_09891_));
 AO22x1_ASAP7_75t_R _17364_ (.A1(_09889_),
    .A2(_09833_),
    .B1(_09891_),
    .B2(_09808_),
    .Y(_01625_));
 BUFx6f_ASAP7_75t_R _17365_ (.A(_09030_),
    .Y(_09892_));
 BUFx6f_ASAP7_75t_R _17366_ (.A(_09031_),
    .Y(_09893_));
 BUFx6f_ASAP7_75t_R _17367_ (.A(_09035_),
    .Y(_09894_));
 AND4x1_ASAP7_75t_R _17368_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_09841_),
    .Y(_09895_));
 INVx1_ASAP7_75t_R _17369_ (.A(_00155_),
    .Y(_09896_));
 AO32x1_ASAP7_75t_R _17370_ (.A1(_09877_),
    .A2(_09811_),
    .A3(_09895_),
    .B1(_09843_),
    .B2(_09896_),
    .Y(_01626_));
 BUFx4f_ASAP7_75t_R _17371_ (.A(_09048_),
    .Y(_09897_));
 BUFx3_ASAP7_75t_R _17372_ (.A(_09051_),
    .Y(_09898_));
 AND3x1_ASAP7_75t_R _17373_ (.A(_09897_),
    .B(_09898_),
    .C(_09850_),
    .Y(_09899_));
 INVx1_ASAP7_75t_R _17374_ (.A(_00121_),
    .Y(_09900_));
 AO32x1_ASAP7_75t_R _17375_ (.A1(_09877_),
    .A2(_09813_),
    .A3(_09899_),
    .B1(_09843_),
    .B2(_09900_),
    .Y(_01627_));
 BUFx4f_ASAP7_75t_R _17376_ (.A(_09063_),
    .Y(_09901_));
 NAND2x1_ASAP7_75t_R _17377_ (.A(_01018_),
    .B(_09833_),
    .Y(_09902_));
 OA21x2_ASAP7_75t_R _17378_ (.A1(_09901_),
    .A2(_09832_),
    .B(_09902_),
    .Y(_01628_));
 BUFx4f_ASAP7_75t_R _17379_ (.A(_09074_),
    .Y(_09903_));
 BUFx4f_ASAP7_75t_R _17380_ (.A(_09077_),
    .Y(_09904_));
 BUFx4f_ASAP7_75t_R _17381_ (.A(_09078_),
    .Y(_09905_));
 AND4x1_ASAP7_75t_R _17382_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_09841_),
    .Y(_09906_));
 INVx1_ASAP7_75t_R _17383_ (.A(_00087_),
    .Y(_09907_));
 AO32x1_ASAP7_75t_R _17384_ (.A1(_09877_),
    .A2(_09816_),
    .A3(_09906_),
    .B1(_09843_),
    .B2(_09907_),
    .Y(_01629_));
 BUFx4f_ASAP7_75t_R _17385_ (.A(_09094_),
    .Y(_09908_));
 BUFx4f_ASAP7_75t_R _17386_ (.A(_09097_),
    .Y(_09909_));
 AND3x1_ASAP7_75t_R _17387_ (.A(_09908_),
    .B(_09909_),
    .C(_09850_),
    .Y(_09910_));
 INVx1_ASAP7_75t_R _17388_ (.A(_00055_),
    .Y(_09911_));
 AO32x1_ASAP7_75t_R _17389_ (.A1(_09877_),
    .A2(_09818_),
    .A3(_09910_),
    .B1(_09843_),
    .B2(_09911_),
    .Y(_01630_));
 BUFx4f_ASAP7_75t_R _17390_ (.A(_09109_),
    .Y(_09912_));
 NAND2x1_ASAP7_75t_R _17391_ (.A(_00985_),
    .B(_09833_),
    .Y(_09913_));
 OA21x2_ASAP7_75t_R _17392_ (.A1(_09912_),
    .A2(_09832_),
    .B(_09913_),
    .Y(_01631_));
 BUFx4f_ASAP7_75t_R _17393_ (.A(_09122_),
    .Y(_09914_));
 NAND2x1_ASAP7_75t_R _17394_ (.A(_00952_),
    .B(_09833_),
    .Y(_09915_));
 OA21x2_ASAP7_75t_R _17395_ (.A1(_09914_),
    .A2(_09832_),
    .B(_09915_),
    .Y(_01632_));
 AND2x2_ASAP7_75t_R _17396_ (.A(_00918_),
    .B(_09843_),
    .Y(_09916_));
 AOI21x1_ASAP7_75t_R _17397_ (.A1(_09822_),
    .A2(_09842_),
    .B(_09916_),
    .Y(_01633_));
 BUFx3_ASAP7_75t_R _17398_ (.A(_09148_),
    .Y(_09917_));
 NOR2x1_ASAP7_75t_R _17399_ (.A(_00885_),
    .B(_09842_),
    .Y(_09918_));
 AO21x1_ASAP7_75t_R _17400_ (.A1(_09917_),
    .A2(_09842_),
    .B(_09918_),
    .Y(_01634_));
 BUFx4f_ASAP7_75t_R _17401_ (.A(_09158_),
    .Y(_09919_));
 NOR2x1_ASAP7_75t_R _17402_ (.A(_00851_),
    .B(_09842_),
    .Y(_09920_));
 AO21x1_ASAP7_75t_R _17403_ (.A1(_09919_),
    .A2(_09842_),
    .B(_09920_),
    .Y(_01635_));
 BUFx4f_ASAP7_75t_R _17404_ (.A(_09173_),
    .Y(_09921_));
 NOR2x1_ASAP7_75t_R _17405_ (.A(_00818_),
    .B(_09842_),
    .Y(_09922_));
 AO21x1_ASAP7_75t_R _17406_ (.A1(_09921_),
    .A2(_09842_),
    .B(_09922_),
    .Y(_01636_));
 BUFx6f_ASAP7_75t_R _17407_ (.A(_09186_),
    .Y(_09923_));
 NAND2x1_ASAP7_75t_R _17408_ (.A(_00784_),
    .B(_09852_),
    .Y(_09924_));
 OA21x2_ASAP7_75t_R _17409_ (.A1(_09923_),
    .A2(_09832_),
    .B(_09924_),
    .Y(_01637_));
 OR3x4_ASAP7_75t_R _17410_ (.A(_07131_),
    .B(_09349_),
    .C(_09830_),
    .Y(_09925_));
 BUFx6f_ASAP7_75t_R _17411_ (.A(_09925_),
    .Y(_09926_));
 BUFx12_ASAP7_75t_R _17412_ (.A(_09925_),
    .Y(_09927_));
 NAND2x1_ASAP7_75t_R _17413_ (.A(_00021_),
    .B(_09927_),
    .Y(_09928_));
 OA21x2_ASAP7_75t_R _17414_ (.A1(_09755_),
    .A2(_09926_),
    .B(_09928_),
    .Y(_01638_));
 NAND2x1_ASAP7_75t_R _17415_ (.A(_00753_),
    .B(_09927_),
    .Y(_09929_));
 OA21x2_ASAP7_75t_R _17416_ (.A1(_09835_),
    .A2(_09926_),
    .B(_09929_),
    .Y(_01639_));
 NAND2x1_ASAP7_75t_R _17417_ (.A(_00720_),
    .B(_09927_),
    .Y(_09930_));
 OA21x2_ASAP7_75t_R _17418_ (.A1(_09837_),
    .A2(_09926_),
    .B(_09930_),
    .Y(_01640_));
 NAND2x1_ASAP7_75t_R _17419_ (.A(_00687_),
    .B(_09927_),
    .Y(_09931_));
 OA21x2_ASAP7_75t_R _17420_ (.A1(_09839_),
    .A2(_09926_),
    .B(_09931_),
    .Y(_01641_));
 NOR2x2_ASAP7_75t_R _17421_ (.A(_09357_),
    .B(_09830_),
    .Y(_09932_));
 BUFx6f_ASAP7_75t_R _17422_ (.A(_09932_),
    .Y(_09933_));
 BUFx6f_ASAP7_75t_R _17423_ (.A(_09925_),
    .Y(_09934_));
 AND2x2_ASAP7_75t_R _17424_ (.A(_00654_),
    .B(_09934_),
    .Y(_09935_));
 AOI21x1_ASAP7_75t_R _17425_ (.A1(_09763_),
    .A2(_09933_),
    .B(_09935_),
    .Y(_01642_));
 NAND2x1_ASAP7_75t_R _17426_ (.A(_00621_),
    .B(_09927_),
    .Y(_09936_));
 OA21x2_ASAP7_75t_R _17427_ (.A1(_09845_),
    .A2(_09926_),
    .B(_09936_),
    .Y(_01643_));
 BUFx12f_ASAP7_75t_R _17428_ (.A(_08765_),
    .Y(_09937_));
 OR2x2_ASAP7_75t_R _17429_ (.A(_00587_),
    .B(_09933_),
    .Y(_09938_));
 OAI21x1_ASAP7_75t_R _17430_ (.A1(_09937_),
    .A2(_09926_),
    .B(_09938_),
    .Y(_01644_));
 BUFx4f_ASAP7_75t_R _17431_ (.A(_09932_),
    .Y(_09939_));
 AND3x1_ASAP7_75t_R _17432_ (.A(_09848_),
    .B(_09849_),
    .C(_09939_),
    .Y(_02246_));
 BUFx10_ASAP7_75t_R _17433_ (.A(_09925_),
    .Y(_02247_));
 INVx1_ASAP7_75t_R _17434_ (.A(_00554_),
    .Y(_02248_));
 AO32x1_ASAP7_75t_R _17435_ (.A1(_09771_),
    .A2(_09548_),
    .A3(_02246_),
    .B1(_02247_),
    .B2(_02248_),
    .Y(_01645_));
 AND2x2_ASAP7_75t_R _17436_ (.A(_09854_),
    .B(_09939_),
    .Y(_02249_));
 INVx1_ASAP7_75t_R _17437_ (.A(_00521_),
    .Y(_02250_));
 AO32x1_ASAP7_75t_R _17438_ (.A1(_09877_),
    .A2(_09776_),
    .A3(_02249_),
    .B1(_02247_),
    .B2(_02250_),
    .Y(_01646_));
 AND3x1_ASAP7_75t_R _17439_ (.A(_09857_),
    .B(_09858_),
    .C(_09939_),
    .Y(_02251_));
 INVx1_ASAP7_75t_R _17440_ (.A(_00488_),
    .Y(_02252_));
 AO32x1_ASAP7_75t_R _17441_ (.A1(_09877_),
    .A2(_09779_),
    .A3(_02251_),
    .B1(_02247_),
    .B2(_02252_),
    .Y(_01647_));
 BUFx4f_ASAP7_75t_R _17442_ (.A(_09809_),
    .Y(_02253_));
 AND3x1_ASAP7_75t_R _17443_ (.A(_09861_),
    .B(_09862_),
    .C(_09939_),
    .Y(_02254_));
 INVx1_ASAP7_75t_R _17444_ (.A(_00455_),
    .Y(_02255_));
 AO32x1_ASAP7_75t_R _17445_ (.A1(_02253_),
    .A2(_09782_),
    .A3(_02254_),
    .B1(_02247_),
    .B2(_02255_),
    .Y(_01648_));
 NAND2x1_ASAP7_75t_R _17446_ (.A(_01052_),
    .B(_09927_),
    .Y(_02256_));
 OA21x2_ASAP7_75t_R _17447_ (.A1(_09865_),
    .A2(_09926_),
    .B(_02256_),
    .Y(_01649_));
 AND2x2_ASAP7_75t_R _17448_ (.A(_09867_),
    .B(_09939_),
    .Y(_02257_));
 INVx1_ASAP7_75t_R _17449_ (.A(_00422_),
    .Y(_02258_));
 AO32x1_ASAP7_75t_R _17450_ (.A1(_02253_),
    .A2(_09786_),
    .A3(_02257_),
    .B1(_02247_),
    .B2(_02258_),
    .Y(_01650_));
 AND3x1_ASAP7_75t_R _17451_ (.A(_09870_),
    .B(_09871_),
    .C(_09939_),
    .Y(_02259_));
 INVx1_ASAP7_75t_R _17452_ (.A(_00389_),
    .Y(_02260_));
 AO32x1_ASAP7_75t_R _17453_ (.A1(_02253_),
    .A2(_09789_),
    .A3(_02259_),
    .B1(_02247_),
    .B2(_02260_),
    .Y(_01651_));
 AND2x2_ASAP7_75t_R _17454_ (.A(_09874_),
    .B(_09939_),
    .Y(_02261_));
 INVx1_ASAP7_75t_R _17455_ (.A(_00356_),
    .Y(_02262_));
 AO32x1_ASAP7_75t_R _17456_ (.A1(_02253_),
    .A2(_09792_),
    .A3(_02261_),
    .B1(_02247_),
    .B2(_02262_),
    .Y(_01652_));
 AND2x2_ASAP7_75t_R _17457_ (.A(_09878_),
    .B(_09939_),
    .Y(_02263_));
 INVx1_ASAP7_75t_R _17458_ (.A(_00322_),
    .Y(_02264_));
 AO32x1_ASAP7_75t_R _17459_ (.A1(_02253_),
    .A2(_09794_),
    .A3(_02263_),
    .B1(_02247_),
    .B2(_02264_),
    .Y(_01653_));
 AND2x2_ASAP7_75t_R _17460_ (.A(_09881_),
    .B(_09932_),
    .Y(_02265_));
 INVx1_ASAP7_75t_R _17461_ (.A(_00289_),
    .Y(_02266_));
 AO32x1_ASAP7_75t_R _17462_ (.A1(_02253_),
    .A2(_09797_),
    .A3(_02265_),
    .B1(_09934_),
    .B2(_02266_),
    .Y(_01654_));
 AND2x2_ASAP7_75t_R _17463_ (.A(_09884_),
    .B(_09932_),
    .Y(_02267_));
 INVx1_ASAP7_75t_R _17464_ (.A(_00256_),
    .Y(_02268_));
 AO32x1_ASAP7_75t_R _17465_ (.A1(_02253_),
    .A2(_09800_),
    .A3(_02267_),
    .B1(_09934_),
    .B2(_02268_),
    .Y(_01655_));
 NOR2x1_ASAP7_75t_R _17466_ (.A(_09804_),
    .B(_09934_),
    .Y(_02269_));
 INVx1_ASAP7_75t_R _17467_ (.A(_00223_),
    .Y(_02270_));
 AO32x1_ASAP7_75t_R _17468_ (.A1(_02253_),
    .A2(_09803_),
    .A3(_02269_),
    .B1(_09934_),
    .B2(_02270_),
    .Y(_01656_));
 INVx1_ASAP7_75t_R _17469_ (.A(_00189_),
    .Y(_02271_));
 AND2x2_ASAP7_75t_R _17470_ (.A(_09890_),
    .B(_09933_),
    .Y(_02272_));
 AO22x1_ASAP7_75t_R _17471_ (.A1(_02271_),
    .A2(_09927_),
    .B1(_02272_),
    .B2(_09808_),
    .Y(_01657_));
 AND4x1_ASAP7_75t_R _17472_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_09932_),
    .Y(_02273_));
 INVx1_ASAP7_75t_R _17473_ (.A(_00156_),
    .Y(_02274_));
 AO32x1_ASAP7_75t_R _17474_ (.A1(_02253_),
    .A2(_09811_),
    .A3(_02273_),
    .B1(_09934_),
    .B2(_02274_),
    .Y(_01658_));
 AND3x1_ASAP7_75t_R _17475_ (.A(_09897_),
    .B(_09898_),
    .C(_09939_),
    .Y(_02275_));
 INVx1_ASAP7_75t_R _17476_ (.A(_00122_),
    .Y(_02276_));
 AO32x1_ASAP7_75t_R _17477_ (.A1(_02253_),
    .A2(_09813_),
    .A3(_02275_),
    .B1(_09934_),
    .B2(_02276_),
    .Y(_01659_));
 NAND2x1_ASAP7_75t_R _17478_ (.A(_01019_),
    .B(_09927_),
    .Y(_02277_));
 OA21x2_ASAP7_75t_R _17479_ (.A1(_09901_),
    .A2(_09926_),
    .B(_02277_),
    .Y(_01660_));
 BUFx4f_ASAP7_75t_R _17480_ (.A(_09809_),
    .Y(_02278_));
 AND4x1_ASAP7_75t_R _17481_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_09932_),
    .Y(_02279_));
 INVx1_ASAP7_75t_R _17482_ (.A(_00088_),
    .Y(_02280_));
 AO32x1_ASAP7_75t_R _17483_ (.A1(_02278_),
    .A2(_09816_),
    .A3(_02279_),
    .B1(_09934_),
    .B2(_02280_),
    .Y(_01661_));
 AND3x1_ASAP7_75t_R _17484_ (.A(_09908_),
    .B(_09909_),
    .C(_09939_),
    .Y(_02281_));
 INVx1_ASAP7_75t_R _17485_ (.A(_00056_),
    .Y(_02282_));
 AO32x1_ASAP7_75t_R _17486_ (.A1(_02278_),
    .A2(_09818_),
    .A3(_02281_),
    .B1(_09934_),
    .B2(_02282_),
    .Y(_01662_));
 NAND2x1_ASAP7_75t_R _17487_ (.A(_00986_),
    .B(_09927_),
    .Y(_02283_));
 OA21x2_ASAP7_75t_R _17488_ (.A1(_09912_),
    .A2(_09926_),
    .B(_02283_),
    .Y(_01663_));
 NAND2x1_ASAP7_75t_R _17489_ (.A(_00953_),
    .B(_02247_),
    .Y(_02284_));
 OA21x2_ASAP7_75t_R _17490_ (.A1(_09914_),
    .A2(_09926_),
    .B(_02284_),
    .Y(_01664_));
 AND2x2_ASAP7_75t_R _17491_ (.A(_00919_),
    .B(_09934_),
    .Y(_02285_));
 AOI21x1_ASAP7_75t_R _17492_ (.A1(_09822_),
    .A2(_09933_),
    .B(_02285_),
    .Y(_01665_));
 NOR2x1_ASAP7_75t_R _17493_ (.A(_00886_),
    .B(_09933_),
    .Y(_02286_));
 AO21x1_ASAP7_75t_R _17494_ (.A1(_09917_),
    .A2(_09933_),
    .B(_02286_),
    .Y(_01666_));
 NOR2x1_ASAP7_75t_R _17495_ (.A(_00852_),
    .B(_09933_),
    .Y(_02287_));
 AO21x1_ASAP7_75t_R _17496_ (.A1(_09919_),
    .A2(_09933_),
    .B(_02287_),
    .Y(_01667_));
 NOR2x1_ASAP7_75t_R _17497_ (.A(_00819_),
    .B(_09933_),
    .Y(_02288_));
 AO21x1_ASAP7_75t_R _17498_ (.A1(_09921_),
    .A2(_09933_),
    .B(_02288_),
    .Y(_01668_));
 NAND2x1_ASAP7_75t_R _17499_ (.A(_00785_),
    .B(_02247_),
    .Y(_02289_));
 OA21x2_ASAP7_75t_R _17500_ (.A1(_09923_),
    .A2(_09927_),
    .B(_02289_),
    .Y(_01669_));
 OR3x4_ASAP7_75t_R _17501_ (.A(_09408_),
    .B(_08601_),
    .C(_09830_),
    .Y(_02290_));
 BUFx4f_ASAP7_75t_R _17502_ (.A(_02290_),
    .Y(_02291_));
 BUFx6f_ASAP7_75t_R _17503_ (.A(_02290_),
    .Y(_02292_));
 NAND2x1_ASAP7_75t_R _17504_ (.A(_00022_),
    .B(_02292_),
    .Y(_02293_));
 OA21x2_ASAP7_75t_R _17505_ (.A1(_09755_),
    .A2(_02291_),
    .B(_02293_),
    .Y(_01670_));
 NAND2x1_ASAP7_75t_R _17506_ (.A(_00754_),
    .B(_02292_),
    .Y(_02294_));
 OA21x2_ASAP7_75t_R _17507_ (.A1(_09835_),
    .A2(_02291_),
    .B(_02294_),
    .Y(_01671_));
 NAND2x1_ASAP7_75t_R _17508_ (.A(_00721_),
    .B(_02292_),
    .Y(_02295_));
 OA21x2_ASAP7_75t_R _17509_ (.A1(_09837_),
    .A2(_02291_),
    .B(_02295_),
    .Y(_01672_));
 NAND2x1_ASAP7_75t_R _17510_ (.A(_00688_),
    .B(_02292_),
    .Y(_02296_));
 OA21x2_ASAP7_75t_R _17511_ (.A1(_09839_),
    .A2(_02291_),
    .B(_02296_),
    .Y(_01673_));
 NOR2x2_ASAP7_75t_R _17512_ (.A(_09416_),
    .B(_09830_),
    .Y(_02297_));
 BUFx6f_ASAP7_75t_R _17513_ (.A(_02297_),
    .Y(_02298_));
 BUFx6f_ASAP7_75t_R _17514_ (.A(_02290_),
    .Y(_02299_));
 AND2x2_ASAP7_75t_R _17515_ (.A(_00655_),
    .B(_02299_),
    .Y(_02300_));
 AOI21x1_ASAP7_75t_R _17516_ (.A1(_09763_),
    .A2(_02298_),
    .B(_02300_),
    .Y(_01674_));
 NAND2x1_ASAP7_75t_R _17517_ (.A(_00622_),
    .B(_02292_),
    .Y(_02301_));
 OA21x2_ASAP7_75t_R _17518_ (.A1(_09845_),
    .A2(_02291_),
    .B(_02301_),
    .Y(_01675_));
 OR2x2_ASAP7_75t_R _17519_ (.A(_00588_),
    .B(_02298_),
    .Y(_02302_));
 OAI21x1_ASAP7_75t_R _17520_ (.A1(_09937_),
    .A2(_02291_),
    .B(_02302_),
    .Y(_01676_));
 AND3x1_ASAP7_75t_R _17521_ (.A(_09848_),
    .B(_09849_),
    .C(_02298_),
    .Y(_02303_));
 BUFx10_ASAP7_75t_R _17522_ (.A(_02290_),
    .Y(_02304_));
 AO32x1_ASAP7_75t_R _17523_ (.A1(_09771_),
    .A2(_09548_),
    .A3(_02303_),
    .B1(_02304_),
    .B2(_05742_),
    .Y(_01677_));
 BUFx4f_ASAP7_75t_R _17524_ (.A(_02297_),
    .Y(_02305_));
 AND2x2_ASAP7_75t_R _17525_ (.A(_09854_),
    .B(_02305_),
    .Y(_02306_));
 INVx1_ASAP7_75t_R _17526_ (.A(_00522_),
    .Y(_02307_));
 AO32x1_ASAP7_75t_R _17527_ (.A1(_02278_),
    .A2(_09776_),
    .A3(_02306_),
    .B1(_02304_),
    .B2(_02307_),
    .Y(_01678_));
 AND3x1_ASAP7_75t_R _17528_ (.A(_09857_),
    .B(_09858_),
    .C(_02305_),
    .Y(_02308_));
 INVx1_ASAP7_75t_R _17529_ (.A(_00489_),
    .Y(_02309_));
 AO32x1_ASAP7_75t_R _17530_ (.A1(_02278_),
    .A2(_09779_),
    .A3(_02308_),
    .B1(_02304_),
    .B2(_02309_),
    .Y(_01679_));
 AND3x1_ASAP7_75t_R _17531_ (.A(_09861_),
    .B(_09862_),
    .C(_02305_),
    .Y(_02310_));
 INVx1_ASAP7_75t_R _17532_ (.A(_00456_),
    .Y(_02311_));
 AO32x1_ASAP7_75t_R _17533_ (.A1(_02278_),
    .A2(_09782_),
    .A3(_02310_),
    .B1(_02304_),
    .B2(_02311_),
    .Y(_01680_));
 NAND2x1_ASAP7_75t_R _17534_ (.A(_01053_),
    .B(_02292_),
    .Y(_02312_));
 OA21x2_ASAP7_75t_R _17535_ (.A1(_09865_),
    .A2(_02291_),
    .B(_02312_),
    .Y(_01681_));
 AND2x2_ASAP7_75t_R _17536_ (.A(_09867_),
    .B(_02305_),
    .Y(_02313_));
 INVx1_ASAP7_75t_R _17537_ (.A(_00423_),
    .Y(_02314_));
 AO32x1_ASAP7_75t_R _17538_ (.A1(_02278_),
    .A2(_09786_),
    .A3(_02313_),
    .B1(_02304_),
    .B2(_02314_),
    .Y(_01682_));
 AND3x1_ASAP7_75t_R _17539_ (.A(_09870_),
    .B(_09871_),
    .C(_02305_),
    .Y(_02315_));
 INVx1_ASAP7_75t_R _17540_ (.A(_00390_),
    .Y(_02316_));
 AO32x1_ASAP7_75t_R _17541_ (.A1(_02278_),
    .A2(_09789_),
    .A3(_02315_),
    .B1(_02304_),
    .B2(_02316_),
    .Y(_01683_));
 AND2x2_ASAP7_75t_R _17542_ (.A(_09874_),
    .B(_02305_),
    .Y(_02317_));
 INVx1_ASAP7_75t_R _17543_ (.A(_00357_),
    .Y(_02318_));
 AO32x1_ASAP7_75t_R _17544_ (.A1(_02278_),
    .A2(_09792_),
    .A3(_02317_),
    .B1(_02304_),
    .B2(_02318_),
    .Y(_01684_));
 AND2x2_ASAP7_75t_R _17545_ (.A(_09878_),
    .B(_02305_),
    .Y(_02319_));
 INVx1_ASAP7_75t_R _17546_ (.A(_00323_),
    .Y(_02320_));
 AO32x1_ASAP7_75t_R _17547_ (.A1(_02278_),
    .A2(_09794_),
    .A3(_02319_),
    .B1(_02304_),
    .B2(_02320_),
    .Y(_01685_));
 AND2x2_ASAP7_75t_R _17548_ (.A(_09881_),
    .B(_02305_),
    .Y(_02321_));
 INVx1_ASAP7_75t_R _17549_ (.A(_00290_),
    .Y(_02322_));
 AO32x1_ASAP7_75t_R _17550_ (.A1(_02278_),
    .A2(_09797_),
    .A3(_02321_),
    .B1(_02299_),
    .B2(_02322_),
    .Y(_01686_));
 BUFx4f_ASAP7_75t_R _17551_ (.A(_09809_),
    .Y(_02323_));
 AND2x2_ASAP7_75t_R _17552_ (.A(_09884_),
    .B(_02297_),
    .Y(_02324_));
 INVx1_ASAP7_75t_R _17553_ (.A(_00257_),
    .Y(_02325_));
 AO32x1_ASAP7_75t_R _17554_ (.A1(_02323_),
    .A2(_09800_),
    .A3(_02324_),
    .B1(_02299_),
    .B2(_02325_),
    .Y(_01687_));
 NOR2x1_ASAP7_75t_R _17555_ (.A(_09804_),
    .B(_02299_),
    .Y(_02326_));
 INVx1_ASAP7_75t_R _17556_ (.A(_00224_),
    .Y(_02327_));
 AO32x1_ASAP7_75t_R _17557_ (.A1(_02323_),
    .A2(_09803_),
    .A3(_02326_),
    .B1(_02299_),
    .B2(_02327_),
    .Y(_01688_));
 INVx1_ASAP7_75t_R _17558_ (.A(_00190_),
    .Y(_02328_));
 AND2x2_ASAP7_75t_R _17559_ (.A(_09890_),
    .B(_02298_),
    .Y(_02329_));
 AO22x1_ASAP7_75t_R _17560_ (.A1(_02328_),
    .A2(_02292_),
    .B1(_02329_),
    .B2(_09808_),
    .Y(_01689_));
 AND4x1_ASAP7_75t_R _17561_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02297_),
    .Y(_02330_));
 AO32x1_ASAP7_75t_R _17562_ (.A1(_02323_),
    .A2(_09811_),
    .A3(_02330_),
    .B1(_02299_),
    .B2(_04485_),
    .Y(_01690_));
 AND3x1_ASAP7_75t_R _17563_ (.A(_09897_),
    .B(_09898_),
    .C(_02305_),
    .Y(_02331_));
 INVx1_ASAP7_75t_R _17564_ (.A(_00123_),
    .Y(_02332_));
 AO32x1_ASAP7_75t_R _17565_ (.A1(_02323_),
    .A2(_09813_),
    .A3(_02331_),
    .B1(_02299_),
    .B2(_02332_),
    .Y(_01691_));
 NAND2x1_ASAP7_75t_R _17566_ (.A(_01020_),
    .B(_02292_),
    .Y(_02333_));
 OA21x2_ASAP7_75t_R _17567_ (.A1(_09901_),
    .A2(_02291_),
    .B(_02333_),
    .Y(_01692_));
 AND4x1_ASAP7_75t_R _17568_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02297_),
    .Y(_02334_));
 INVx1_ASAP7_75t_R _17569_ (.A(_00089_),
    .Y(_02335_));
 AO32x1_ASAP7_75t_R _17570_ (.A1(_02323_),
    .A2(_09816_),
    .A3(_02334_),
    .B1(_02299_),
    .B2(_02335_),
    .Y(_01693_));
 AND3x1_ASAP7_75t_R _17571_ (.A(_09908_),
    .B(_09909_),
    .C(_02305_),
    .Y(_02336_));
 INVx1_ASAP7_75t_R _17572_ (.A(_00057_),
    .Y(_02337_));
 AO32x1_ASAP7_75t_R _17573_ (.A1(_02323_),
    .A2(_09818_),
    .A3(_02336_),
    .B1(_02299_),
    .B2(_02337_),
    .Y(_01694_));
 NAND2x1_ASAP7_75t_R _17574_ (.A(_00987_),
    .B(_02292_),
    .Y(_02338_));
 OA21x2_ASAP7_75t_R _17575_ (.A1(_09912_),
    .A2(_02291_),
    .B(_02338_),
    .Y(_01695_));
 NAND2x1_ASAP7_75t_R _17576_ (.A(_00954_),
    .B(_02304_),
    .Y(_02339_));
 OA21x2_ASAP7_75t_R _17577_ (.A1(_09914_),
    .A2(_02291_),
    .B(_02339_),
    .Y(_01696_));
 AND2x2_ASAP7_75t_R _17578_ (.A(_00920_),
    .B(_02299_),
    .Y(_02340_));
 AOI21x1_ASAP7_75t_R _17579_ (.A1(_09822_),
    .A2(_02298_),
    .B(_02340_),
    .Y(_01697_));
 NOR2x1_ASAP7_75t_R _17580_ (.A(_00887_),
    .B(_02298_),
    .Y(_02341_));
 AO21x1_ASAP7_75t_R _17581_ (.A1(_09917_),
    .A2(_02298_),
    .B(_02341_),
    .Y(_01698_));
 AND2x2_ASAP7_75t_R _17582_ (.A(_06541_),
    .B(_02290_),
    .Y(_02342_));
 AO21x1_ASAP7_75t_R _17583_ (.A1(_09919_),
    .A2(_02298_),
    .B(_02342_),
    .Y(_01699_));
 NOR2x1_ASAP7_75t_R _17584_ (.A(_00820_),
    .B(_02298_),
    .Y(_02343_));
 AO21x1_ASAP7_75t_R _17585_ (.A1(_09921_),
    .A2(_02298_),
    .B(_02343_),
    .Y(_01700_));
 NAND2x1_ASAP7_75t_R _17586_ (.A(_00786_),
    .B(_02304_),
    .Y(_02344_));
 OA21x2_ASAP7_75t_R _17587_ (.A1(_09923_),
    .A2(_02292_),
    .B(_02344_),
    .Y(_01701_));
 OR3x4_ASAP7_75t_R _17588_ (.A(_09408_),
    .B(_09349_),
    .C(_09830_),
    .Y(_02345_));
 BUFx6f_ASAP7_75t_R _17589_ (.A(_02345_),
    .Y(_02346_));
 BUFx6f_ASAP7_75t_R _17590_ (.A(_02345_),
    .Y(_02347_));
 NAND2x1_ASAP7_75t_R _17591_ (.A(_00023_),
    .B(_02347_),
    .Y(_02348_));
 OA21x2_ASAP7_75t_R _17592_ (.A1(_09755_),
    .A2(_02346_),
    .B(_02348_),
    .Y(_01702_));
 NAND2x1_ASAP7_75t_R _17593_ (.A(_00755_),
    .B(_02347_),
    .Y(_02349_));
 OA21x2_ASAP7_75t_R _17594_ (.A1(_09835_),
    .A2(_02346_),
    .B(_02349_),
    .Y(_01703_));
 NAND2x1_ASAP7_75t_R _17595_ (.A(_00722_),
    .B(_02347_),
    .Y(_02350_));
 OA21x2_ASAP7_75t_R _17596_ (.A1(_09837_),
    .A2(_02346_),
    .B(_02350_),
    .Y(_01704_));
 NAND2x1_ASAP7_75t_R _17597_ (.A(_00689_),
    .B(_02347_),
    .Y(_02351_));
 OA21x2_ASAP7_75t_R _17598_ (.A1(_09839_),
    .A2(_02346_),
    .B(_02351_),
    .Y(_01705_));
 NOR2x2_ASAP7_75t_R _17599_ (.A(_09473_),
    .B(_09830_),
    .Y(_02352_));
 BUFx6f_ASAP7_75t_R _17600_ (.A(_02352_),
    .Y(_02353_));
 BUFx6f_ASAP7_75t_R _17601_ (.A(_02345_),
    .Y(_02354_));
 AND2x2_ASAP7_75t_R _17602_ (.A(_00656_),
    .B(_02354_),
    .Y(_02355_));
 AOI21x1_ASAP7_75t_R _17603_ (.A1(_09763_),
    .A2(_02353_),
    .B(_02355_),
    .Y(_01706_));
 NAND2x1_ASAP7_75t_R _17604_ (.A(_00623_),
    .B(_02347_),
    .Y(_02356_));
 OA21x2_ASAP7_75t_R _17605_ (.A1(_09845_),
    .A2(_02346_),
    .B(_02356_),
    .Y(_01707_));
 OR2x2_ASAP7_75t_R _17606_ (.A(_00589_),
    .B(_02353_),
    .Y(_02357_));
 OAI21x1_ASAP7_75t_R _17607_ (.A1(_09937_),
    .A2(_02346_),
    .B(_02357_),
    .Y(_01708_));
 BUFx4f_ASAP7_75t_R _17608_ (.A(_02352_),
    .Y(_02358_));
 AND3x1_ASAP7_75t_R _17609_ (.A(_09848_),
    .B(_09849_),
    .C(_02358_),
    .Y(_02359_));
 BUFx10_ASAP7_75t_R _17610_ (.A(_02345_),
    .Y(_02360_));
 AO32x1_ASAP7_75t_R _17611_ (.A1(_09771_),
    .A2(_09548_),
    .A3(_02359_),
    .B1(_02360_),
    .B2(_05744_),
    .Y(_01709_));
 AND2x2_ASAP7_75t_R _17612_ (.A(_09854_),
    .B(_02358_),
    .Y(_02361_));
 INVx1_ASAP7_75t_R _17613_ (.A(_00523_),
    .Y(_02362_));
 AO32x1_ASAP7_75t_R _17614_ (.A1(_02323_),
    .A2(_09776_),
    .A3(_02361_),
    .B1(_02360_),
    .B2(_02362_),
    .Y(_01710_));
 AND3x1_ASAP7_75t_R _17615_ (.A(_09857_),
    .B(_09858_),
    .C(_02358_),
    .Y(_02363_));
 INVx1_ASAP7_75t_R _17616_ (.A(_00490_),
    .Y(_02364_));
 AO32x1_ASAP7_75t_R _17617_ (.A1(_02323_),
    .A2(_09779_),
    .A3(_02363_),
    .B1(_02360_),
    .B2(_02364_),
    .Y(_01711_));
 AND3x1_ASAP7_75t_R _17618_ (.A(_09861_),
    .B(_09862_),
    .C(_02358_),
    .Y(_02365_));
 INVx1_ASAP7_75t_R _17619_ (.A(_00457_),
    .Y(_02366_));
 AO32x1_ASAP7_75t_R _17620_ (.A1(_02323_),
    .A2(_09782_),
    .A3(_02365_),
    .B1(_02360_),
    .B2(_02366_),
    .Y(_01712_));
 NAND2x1_ASAP7_75t_R _17621_ (.A(_01054_),
    .B(_02347_),
    .Y(_02367_));
 OA21x2_ASAP7_75t_R _17622_ (.A1(_09865_),
    .A2(_02346_),
    .B(_02367_),
    .Y(_01713_));
 AND2x2_ASAP7_75t_R _17623_ (.A(_09867_),
    .B(_02358_),
    .Y(_02368_));
 INVx1_ASAP7_75t_R _17624_ (.A(_00424_),
    .Y(_02369_));
 AO32x1_ASAP7_75t_R _17625_ (.A1(_02323_),
    .A2(_09786_),
    .A3(_02368_),
    .B1(_02360_),
    .B2(_02369_),
    .Y(_01714_));
 BUFx4f_ASAP7_75t_R _17626_ (.A(_09809_),
    .Y(_02370_));
 AND3x1_ASAP7_75t_R _17627_ (.A(_09870_),
    .B(_09871_),
    .C(_02358_),
    .Y(_02371_));
 INVx1_ASAP7_75t_R _17628_ (.A(_00391_),
    .Y(_02372_));
 AO32x1_ASAP7_75t_R _17629_ (.A1(_02370_),
    .A2(_09789_),
    .A3(_02371_),
    .B1(_02360_),
    .B2(_02372_),
    .Y(_01715_));
 AND2x2_ASAP7_75t_R _17630_ (.A(_09874_),
    .B(_02358_),
    .Y(_02373_));
 INVx1_ASAP7_75t_R _17631_ (.A(_00358_),
    .Y(_02374_));
 AO32x1_ASAP7_75t_R _17632_ (.A1(_02370_),
    .A2(_09792_),
    .A3(_02373_),
    .B1(_02360_),
    .B2(_02374_),
    .Y(_01716_));
 AND2x2_ASAP7_75t_R _17633_ (.A(_09878_),
    .B(_02358_),
    .Y(_02375_));
 INVx1_ASAP7_75t_R _17634_ (.A(_00324_),
    .Y(_02376_));
 AO32x1_ASAP7_75t_R _17635_ (.A1(_02370_),
    .A2(_09794_),
    .A3(_02375_),
    .B1(_02360_),
    .B2(_02376_),
    .Y(_01717_));
 AND2x2_ASAP7_75t_R _17636_ (.A(_09881_),
    .B(_02352_),
    .Y(_02377_));
 INVx1_ASAP7_75t_R _17637_ (.A(_00291_),
    .Y(_02378_));
 AO32x1_ASAP7_75t_R _17638_ (.A1(_02370_),
    .A2(_09797_),
    .A3(_02377_),
    .B1(_02354_),
    .B2(_02378_),
    .Y(_01718_));
 AND2x2_ASAP7_75t_R _17639_ (.A(_09884_),
    .B(_02352_),
    .Y(_02379_));
 INVx1_ASAP7_75t_R _17640_ (.A(_00258_),
    .Y(_02380_));
 AO32x1_ASAP7_75t_R _17641_ (.A1(_02370_),
    .A2(_09800_),
    .A3(_02379_),
    .B1(_02354_),
    .B2(_02380_),
    .Y(_01719_));
 NOR2x1_ASAP7_75t_R _17642_ (.A(_09804_),
    .B(_02354_),
    .Y(_02381_));
 INVx1_ASAP7_75t_R _17643_ (.A(_00225_),
    .Y(_02382_));
 AO32x1_ASAP7_75t_R _17644_ (.A1(_02370_),
    .A2(_09803_),
    .A3(_02381_),
    .B1(_02354_),
    .B2(_02382_),
    .Y(_01720_));
 INVx1_ASAP7_75t_R _17645_ (.A(_00191_),
    .Y(_02383_));
 AND2x2_ASAP7_75t_R _17646_ (.A(_09890_),
    .B(_02353_),
    .Y(_02384_));
 AO22x1_ASAP7_75t_R _17647_ (.A1(_02383_),
    .A2(_02347_),
    .B1(_02384_),
    .B2(_09808_),
    .Y(_01721_));
 AND4x1_ASAP7_75t_R _17648_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02352_),
    .Y(_02385_));
 AO32x1_ASAP7_75t_R _17649_ (.A1(_02370_),
    .A2(_09811_),
    .A3(_02385_),
    .B1(_02354_),
    .B2(_04487_),
    .Y(_01722_));
 AND3x1_ASAP7_75t_R _17650_ (.A(_09897_),
    .B(_09898_),
    .C(_02358_),
    .Y(_02386_));
 INVx1_ASAP7_75t_R _17651_ (.A(_00124_),
    .Y(_02387_));
 AO32x1_ASAP7_75t_R _17652_ (.A1(_02370_),
    .A2(_09813_),
    .A3(_02386_),
    .B1(_02354_),
    .B2(_02387_),
    .Y(_01723_));
 NAND2x1_ASAP7_75t_R _17653_ (.A(_01021_),
    .B(_02347_),
    .Y(_02388_));
 OA21x2_ASAP7_75t_R _17654_ (.A1(_09901_),
    .A2(_02346_),
    .B(_02388_),
    .Y(_01724_));
 AND4x1_ASAP7_75t_R _17655_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02352_),
    .Y(_02389_));
 INVx1_ASAP7_75t_R _17656_ (.A(_00090_),
    .Y(_02390_));
 AO32x1_ASAP7_75t_R _17657_ (.A1(_02370_),
    .A2(_09816_),
    .A3(_02389_),
    .B1(_02354_),
    .B2(_02390_),
    .Y(_01725_));
 AND3x1_ASAP7_75t_R _17658_ (.A(_09908_),
    .B(_09909_),
    .C(_02358_),
    .Y(_02391_));
 INVx1_ASAP7_75t_R _17659_ (.A(_00058_),
    .Y(_02392_));
 AO32x1_ASAP7_75t_R _17660_ (.A1(_02370_),
    .A2(_09818_),
    .A3(_02391_),
    .B1(_02354_),
    .B2(_02392_),
    .Y(_01726_));
 NAND2x1_ASAP7_75t_R _17661_ (.A(_00988_),
    .B(_02347_),
    .Y(_02393_));
 OA21x2_ASAP7_75t_R _17662_ (.A1(_09912_),
    .A2(_02346_),
    .B(_02393_),
    .Y(_01727_));
 NAND2x1_ASAP7_75t_R _17663_ (.A(_00955_),
    .B(_02360_),
    .Y(_02394_));
 OA21x2_ASAP7_75t_R _17664_ (.A1(_09914_),
    .A2(_02346_),
    .B(_02394_),
    .Y(_01728_));
 AND2x2_ASAP7_75t_R _17665_ (.A(_00921_),
    .B(_02354_),
    .Y(_02395_));
 AOI21x1_ASAP7_75t_R _17666_ (.A1(_09822_),
    .A2(_02353_),
    .B(_02395_),
    .Y(_01729_));
 NOR2x1_ASAP7_75t_R _17667_ (.A(_00888_),
    .B(_02353_),
    .Y(_02396_));
 AO21x1_ASAP7_75t_R _17668_ (.A1(_09917_),
    .A2(_02353_),
    .B(_02396_),
    .Y(_01730_));
 NOR2x1_ASAP7_75t_R _17669_ (.A(_00854_),
    .B(_02353_),
    .Y(_02397_));
 AO21x1_ASAP7_75t_R _17670_ (.A1(_09919_),
    .A2(_02353_),
    .B(_02397_),
    .Y(_01731_));
 NOR2x1_ASAP7_75t_R _17671_ (.A(_00821_),
    .B(_02353_),
    .Y(_02398_));
 AO21x1_ASAP7_75t_R _17672_ (.A1(_09921_),
    .A2(_02353_),
    .B(_02398_),
    .Y(_01732_));
 NAND2x1_ASAP7_75t_R _17673_ (.A(_00787_),
    .B(_02360_),
    .Y(_02399_));
 OA21x2_ASAP7_75t_R _17674_ (.A1(_09923_),
    .A2(_02347_),
    .B(_02399_),
    .Y(_01733_));
 AND3x2_ASAP7_75t_R _17675_ (.A(net2),
    .B(_06807_),
    .C(_09530_),
    .Y(_02400_));
 BUFx12f_ASAP7_75t_R _17676_ (.A(_02400_),
    .Y(_02401_));
 NAND2x2_ASAP7_75t_R _17677_ (.A(_09528_),
    .B(_02401_),
    .Y(_02402_));
 BUFx6f_ASAP7_75t_R _17678_ (.A(_02402_),
    .Y(_02403_));
 BUFx6f_ASAP7_75t_R _17679_ (.A(_02401_),
    .Y(_02404_));
 AO21x1_ASAP7_75t_R _17680_ (.A1(_09543_),
    .A2(_02404_),
    .B(_03751_),
    .Y(_02405_));
 OA21x2_ASAP7_75t_R _17681_ (.A1(_09755_),
    .A2(_02403_),
    .B(_02405_),
    .Y(_01734_));
 AO21x1_ASAP7_75t_R _17682_ (.A1(_09543_),
    .A2(_02404_),
    .B(_06295_),
    .Y(_02406_));
 OA21x2_ASAP7_75t_R _17683_ (.A1(_09835_),
    .A2(_02403_),
    .B(_02406_),
    .Y(_01735_));
 AO21x1_ASAP7_75t_R _17684_ (.A1(_09543_),
    .A2(_02404_),
    .B(_06213_),
    .Y(_02407_));
 OA21x2_ASAP7_75t_R _17685_ (.A1(_09837_),
    .A2(_02403_),
    .B(_02407_),
    .Y(_01736_));
 BUFx12_ASAP7_75t_R _17686_ (.A(_02402_),
    .Y(_02408_));
 NAND2x1_ASAP7_75t_R _17687_ (.A(_00690_),
    .B(_02408_),
    .Y(_02409_));
 OA21x2_ASAP7_75t_R _17688_ (.A1(_09839_),
    .A2(_02403_),
    .B(_02409_),
    .Y(_01737_));
 AND2x2_ASAP7_75t_R _17689_ (.A(_09528_),
    .B(_02401_),
    .Y(_02410_));
 BUFx6f_ASAP7_75t_R _17690_ (.A(_02410_),
    .Y(_02411_));
 AND2x2_ASAP7_75t_R _17691_ (.A(_00657_),
    .B(_02402_),
    .Y(_02412_));
 AOI21x1_ASAP7_75t_R _17692_ (.A1(_09763_),
    .A2(_02411_),
    .B(_02412_),
    .Y(_01738_));
 AO21x1_ASAP7_75t_R _17693_ (.A1(_09543_),
    .A2(_02404_),
    .B(_05895_),
    .Y(_02413_));
 OA21x2_ASAP7_75t_R _17694_ (.A1(_09845_),
    .A2(_02403_),
    .B(_02413_),
    .Y(_01739_));
 AND2x2_ASAP7_75t_R _17695_ (.A(_00590_),
    .B(_02402_),
    .Y(_02414_));
 AOI21x1_ASAP7_75t_R _17696_ (.A1(_09769_),
    .A2(_02411_),
    .B(_02414_),
    .Y(_01740_));
 AND3x1_ASAP7_75t_R _17697_ (.A(_09848_),
    .B(_09849_),
    .C(_02411_),
    .Y(_02415_));
 AO32x1_ASAP7_75t_R _17698_ (.A1(_09771_),
    .A2(_09548_),
    .A3(_02415_),
    .B1(_02408_),
    .B2(_05652_),
    .Y(_01741_));
 BUFx4f_ASAP7_75t_R _17699_ (.A(_09809_),
    .Y(_02416_));
 BUFx4f_ASAP7_75t_R _17700_ (.A(_02410_),
    .Y(_02417_));
 AND2x2_ASAP7_75t_R _17701_ (.A(_09854_),
    .B(_02417_),
    .Y(_02418_));
 AO32x1_ASAP7_75t_R _17702_ (.A1(_02416_),
    .A2(_09776_),
    .A3(_02418_),
    .B1(_02408_),
    .B2(_05624_),
    .Y(_01742_));
 AND3x1_ASAP7_75t_R _17703_ (.A(_09857_),
    .B(_09858_),
    .C(_02411_),
    .Y(_02419_));
 AO32x1_ASAP7_75t_R _17704_ (.A1(_02416_),
    .A2(_09779_),
    .A3(_02419_),
    .B1(_02408_),
    .B2(_05516_),
    .Y(_01743_));
 AND3x1_ASAP7_75t_R _17705_ (.A(_09861_),
    .B(_09862_),
    .C(_02411_),
    .Y(_02420_));
 AO32x1_ASAP7_75t_R _17706_ (.A1(_02416_),
    .A2(_09782_),
    .A3(_02420_),
    .B1(_02408_),
    .B2(_05416_),
    .Y(_01744_));
 NAND2x1_ASAP7_75t_R _17707_ (.A(_01055_),
    .B(_02408_),
    .Y(_02421_));
 OA21x2_ASAP7_75t_R _17708_ (.A1(_09865_),
    .A2(_02403_),
    .B(_02421_),
    .Y(_01745_));
 AND2x2_ASAP7_75t_R _17709_ (.A(_09867_),
    .B(_02417_),
    .Y(_02422_));
 INVx1_ASAP7_75t_R _17710_ (.A(_00425_),
    .Y(_02423_));
 AO32x1_ASAP7_75t_R _17711_ (.A1(_02416_),
    .A2(_09786_),
    .A3(_02422_),
    .B1(_02408_),
    .B2(_02423_),
    .Y(_01746_));
 AND3x1_ASAP7_75t_R _17712_ (.A(_09870_),
    .B(_09871_),
    .C(_02417_),
    .Y(_02424_));
 BUFx3_ASAP7_75t_R _17713_ (.A(_02402_),
    .Y(_02425_));
 AO32x1_ASAP7_75t_R _17714_ (.A1(_02416_),
    .A2(_09789_),
    .A3(_02424_),
    .B1(_02425_),
    .B2(_05167_),
    .Y(_01747_));
 AND2x2_ASAP7_75t_R _17715_ (.A(_09874_),
    .B(_02417_),
    .Y(_02426_));
 AO32x1_ASAP7_75t_R _17716_ (.A1(_02416_),
    .A2(_09792_),
    .A3(_02426_),
    .B1(_02425_),
    .B2(_05107_),
    .Y(_01748_));
 AND2x2_ASAP7_75t_R _17717_ (.A(_09878_),
    .B(_02417_),
    .Y(_02427_));
 AO32x1_ASAP7_75t_R _17718_ (.A1(_02416_),
    .A2(_09794_),
    .A3(_02427_),
    .B1(_02425_),
    .B2(_05017_),
    .Y(_01749_));
 AND2x2_ASAP7_75t_R _17719_ (.A(_09881_),
    .B(_02417_),
    .Y(_02428_));
 AO32x1_ASAP7_75t_R _17720_ (.A1(_02416_),
    .A2(_09797_),
    .A3(_02428_),
    .B1(_02425_),
    .B2(_04908_),
    .Y(_01750_));
 AND2x2_ASAP7_75t_R _17721_ (.A(_09884_),
    .B(_02417_),
    .Y(_02429_));
 AO32x1_ASAP7_75t_R _17722_ (.A1(_02416_),
    .A2(_09800_),
    .A3(_02429_),
    .B1(_02425_),
    .B2(_04798_),
    .Y(_01751_));
 NOR2x1_ASAP7_75t_R _17723_ (.A(_09804_),
    .B(_02402_),
    .Y(_02430_));
 AO32x1_ASAP7_75t_R _17724_ (.A1(_02416_),
    .A2(_09803_),
    .A3(_02430_),
    .B1(_02425_),
    .B2(_04686_),
    .Y(_01752_));
 AND2x2_ASAP7_75t_R _17725_ (.A(_09890_),
    .B(_02411_),
    .Y(_02431_));
 AO22x1_ASAP7_75t_R _17726_ (.A1(_04574_),
    .A2(_02408_),
    .B1(_02431_),
    .B2(_09808_),
    .Y(_01753_));
 BUFx4f_ASAP7_75t_R _17727_ (.A(_09809_),
    .Y(_02432_));
 AND4x1_ASAP7_75t_R _17728_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02417_),
    .Y(_02433_));
 INVx1_ASAP7_75t_R _17729_ (.A(_00159_),
    .Y(_02434_));
 AO32x1_ASAP7_75t_R _17730_ (.A1(_02432_),
    .A2(_09811_),
    .A3(_02433_),
    .B1(_02425_),
    .B2(_02434_),
    .Y(_01754_));
 AND3x1_ASAP7_75t_R _17731_ (.A(_09897_),
    .B(_09898_),
    .C(_02417_),
    .Y(_02435_));
 AO32x1_ASAP7_75t_R _17732_ (.A1(_02432_),
    .A2(_09813_),
    .A3(_02435_),
    .B1(_02425_),
    .B2(_04323_),
    .Y(_01755_));
 NAND2x1_ASAP7_75t_R _17733_ (.A(_01022_),
    .B(_02408_),
    .Y(_02436_));
 OA21x2_ASAP7_75t_R _17734_ (.A1(_09901_),
    .A2(_02403_),
    .B(_02436_),
    .Y(_01756_));
 AND4x1_ASAP7_75t_R _17735_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02410_),
    .Y(_02437_));
 AO32x1_ASAP7_75t_R _17736_ (.A1(_02432_),
    .A2(_09816_),
    .A3(_02437_),
    .B1(_02425_),
    .B2(_04217_),
    .Y(_01757_));
 AND3x1_ASAP7_75t_R _17737_ (.A(_09908_),
    .B(_09909_),
    .C(_02417_),
    .Y(_02438_));
 INVx1_ASAP7_75t_R _17738_ (.A(_00059_),
    .Y(_02439_));
 AO32x1_ASAP7_75t_R _17739_ (.A1(_02432_),
    .A2(_09818_),
    .A3(_02438_),
    .B1(_02425_),
    .B2(_02439_),
    .Y(_01758_));
 NAND2x1_ASAP7_75t_R _17740_ (.A(_00989_),
    .B(_02408_),
    .Y(_02440_));
 OA21x2_ASAP7_75t_R _17741_ (.A1(_09912_),
    .A2(_02403_),
    .B(_02440_),
    .Y(_01759_));
 AO21x1_ASAP7_75t_R _17742_ (.A1(_09543_),
    .A2(_02404_),
    .B(_06848_),
    .Y(_02441_));
 OA21x2_ASAP7_75t_R _17743_ (.A1(_09914_),
    .A2(_02403_),
    .B(_02441_),
    .Y(_01760_));
 AND2x2_ASAP7_75t_R _17744_ (.A(_00922_),
    .B(_02402_),
    .Y(_02442_));
 AOI21x1_ASAP7_75t_R _17745_ (.A1(_09822_),
    .A2(_02411_),
    .B(_02442_),
    .Y(_01761_));
 AND2x2_ASAP7_75t_R _17746_ (.A(_06696_),
    .B(_02402_),
    .Y(_02443_));
 AO21x1_ASAP7_75t_R _17747_ (.A1(_09917_),
    .A2(_02411_),
    .B(_02443_),
    .Y(_01762_));
 AND2x2_ASAP7_75t_R _17748_ (.A(_06525_),
    .B(_02402_),
    .Y(_02444_));
 AO21x1_ASAP7_75t_R _17749_ (.A1(_09919_),
    .A2(_02411_),
    .B(_02444_),
    .Y(_01763_));
 AND2x2_ASAP7_75t_R _17750_ (.A(_06500_),
    .B(_02402_),
    .Y(_02445_));
 AO21x1_ASAP7_75t_R _17751_ (.A1(_09921_),
    .A2(_02411_),
    .B(_02445_),
    .Y(_01764_));
 AO21x1_ASAP7_75t_R _17752_ (.A1(_09529_),
    .A2(_02404_),
    .B(_06405_),
    .Y(_02446_));
 OA21x2_ASAP7_75t_R _17753_ (.A1(_09923_),
    .A2(_02403_),
    .B(_02446_),
    .Y(_01765_));
 NAND2x2_ASAP7_75t_R _17754_ (.A(_09590_),
    .B(_02401_),
    .Y(_02447_));
 BUFx6f_ASAP7_75t_R _17755_ (.A(_02447_),
    .Y(_02448_));
 AO21x1_ASAP7_75t_R _17756_ (.A1(_09597_),
    .A2(_02404_),
    .B(_03743_),
    .Y(_02449_));
 OA21x2_ASAP7_75t_R _17757_ (.A1(_09755_),
    .A2(_02448_),
    .B(_02449_),
    .Y(_01766_));
 BUFx10_ASAP7_75t_R _17758_ (.A(_02447_),
    .Y(_02450_));
 NAND2x1_ASAP7_75t_R _17759_ (.A(_00757_),
    .B(_02450_),
    .Y(_02451_));
 OA21x2_ASAP7_75t_R _17760_ (.A1(_09835_),
    .A2(_02448_),
    .B(_02451_),
    .Y(_01767_));
 NAND2x1_ASAP7_75t_R _17761_ (.A(_00724_),
    .B(_02450_),
    .Y(_02452_));
 OA21x2_ASAP7_75t_R _17762_ (.A1(_09837_),
    .A2(_02448_),
    .B(_02452_),
    .Y(_01768_));
 NAND2x1_ASAP7_75t_R _17763_ (.A(_00691_),
    .B(_02450_),
    .Y(_02453_));
 OA21x2_ASAP7_75t_R _17764_ (.A1(_09839_),
    .A2(_02448_),
    .B(_02453_),
    .Y(_01769_));
 AND2x4_ASAP7_75t_R _17765_ (.A(_09589_),
    .B(_02401_),
    .Y(_02454_));
 BUFx6f_ASAP7_75t_R _17766_ (.A(_02454_),
    .Y(_02455_));
 BUFx6f_ASAP7_75t_R _17767_ (.A(_02447_),
    .Y(_02456_));
 AND2x2_ASAP7_75t_R _17768_ (.A(_00658_),
    .B(_02456_),
    .Y(_02457_));
 AOI21x1_ASAP7_75t_R _17769_ (.A1(_09763_),
    .A2(_02455_),
    .B(_02457_),
    .Y(_01770_));
 NAND2x1_ASAP7_75t_R _17770_ (.A(_00625_),
    .B(_02450_),
    .Y(_02458_));
 OA21x2_ASAP7_75t_R _17771_ (.A1(_09845_),
    .A2(_02448_),
    .B(_02458_),
    .Y(_01771_));
 AO21x1_ASAP7_75t_R _17772_ (.A1(_09597_),
    .A2(_02404_),
    .B(_00591_),
    .Y(_02459_));
 OAI21x1_ASAP7_75t_R _17773_ (.A1(_09937_),
    .A2(_02448_),
    .B(_02459_),
    .Y(_01772_));
 BUFx6f_ASAP7_75t_R _17774_ (.A(_09547_),
    .Y(_02460_));
 AND3x1_ASAP7_75t_R _17775_ (.A(_09848_),
    .B(_09849_),
    .C(_02455_),
    .Y(_02461_));
 BUFx6f_ASAP7_75t_R _17776_ (.A(_02447_),
    .Y(_02462_));
 AO32x1_ASAP7_75t_R _17777_ (.A1(_09771_),
    .A2(_02460_),
    .A3(_02461_),
    .B1(_02462_),
    .B2(_05657_),
    .Y(_01773_));
 BUFx4f_ASAP7_75t_R _17778_ (.A(_02454_),
    .Y(_02463_));
 AND2x2_ASAP7_75t_R _17779_ (.A(_09854_),
    .B(_02463_),
    .Y(_02464_));
 INVx1_ASAP7_75t_R _17780_ (.A(_00525_),
    .Y(_02465_));
 AO32x1_ASAP7_75t_R _17781_ (.A1(_02432_),
    .A2(_09776_),
    .A3(_02464_),
    .B1(_02462_),
    .B2(_02465_),
    .Y(_01774_));
 AND3x1_ASAP7_75t_R _17782_ (.A(_09857_),
    .B(_09858_),
    .C(_02455_),
    .Y(_02466_));
 INVx1_ASAP7_75t_R _17783_ (.A(_00492_),
    .Y(_02467_));
 AO32x1_ASAP7_75t_R _17784_ (.A1(_02432_),
    .A2(_09779_),
    .A3(_02466_),
    .B1(_02462_),
    .B2(_02467_),
    .Y(_01775_));
 AND3x1_ASAP7_75t_R _17785_ (.A(_09861_),
    .B(_09862_),
    .C(_02463_),
    .Y(_02468_));
 INVx1_ASAP7_75t_R _17786_ (.A(_00459_),
    .Y(_02469_));
 AO32x1_ASAP7_75t_R _17787_ (.A1(_02432_),
    .A2(_09782_),
    .A3(_02468_),
    .B1(_02462_),
    .B2(_02469_),
    .Y(_01776_));
 NAND2x1_ASAP7_75t_R _17788_ (.A(_01056_),
    .B(_02450_),
    .Y(_02470_));
 OA21x2_ASAP7_75t_R _17789_ (.A1(_09865_),
    .A2(_02448_),
    .B(_02470_),
    .Y(_01777_));
 AND2x2_ASAP7_75t_R _17790_ (.A(_09867_),
    .B(_02463_),
    .Y(_02471_));
 INVx1_ASAP7_75t_R _17791_ (.A(_00426_),
    .Y(_02472_));
 AO32x1_ASAP7_75t_R _17792_ (.A1(_02432_),
    .A2(_09786_),
    .A3(_02471_),
    .B1(_02462_),
    .B2(_02472_),
    .Y(_01778_));
 AND3x1_ASAP7_75t_R _17793_ (.A(_09870_),
    .B(_09871_),
    .C(_02463_),
    .Y(_02473_));
 AO32x1_ASAP7_75t_R _17794_ (.A1(_02432_),
    .A2(_09789_),
    .A3(_02473_),
    .B1(_02462_),
    .B2(_05172_),
    .Y(_01779_));
 AND2x2_ASAP7_75t_R _17795_ (.A(_09874_),
    .B(_02463_),
    .Y(_02474_));
 INVx1_ASAP7_75t_R _17796_ (.A(_00360_),
    .Y(_02475_));
 AO32x1_ASAP7_75t_R _17797_ (.A1(_02432_),
    .A2(_09792_),
    .A3(_02474_),
    .B1(_02462_),
    .B2(_02475_),
    .Y(_01780_));
 BUFx4f_ASAP7_75t_R _17798_ (.A(_09809_),
    .Y(_02476_));
 AND2x2_ASAP7_75t_R _17799_ (.A(_09878_),
    .B(_02463_),
    .Y(_02477_));
 INVx1_ASAP7_75t_R _17800_ (.A(_00326_),
    .Y(_02478_));
 AO32x1_ASAP7_75t_R _17801_ (.A1(_02476_),
    .A2(_09794_),
    .A3(_02477_),
    .B1(_02462_),
    .B2(_02478_),
    .Y(_01781_));
 AND2x2_ASAP7_75t_R _17802_ (.A(_09881_),
    .B(_02463_),
    .Y(_02479_));
 INVx1_ASAP7_75t_R _17803_ (.A(_00293_),
    .Y(_02480_));
 AO32x1_ASAP7_75t_R _17804_ (.A1(_02476_),
    .A2(_09797_),
    .A3(_02479_),
    .B1(_02462_),
    .B2(_02480_),
    .Y(_01782_));
 AND2x2_ASAP7_75t_R _17805_ (.A(_09884_),
    .B(_02463_),
    .Y(_02481_));
 INVx1_ASAP7_75t_R _17806_ (.A(_00260_),
    .Y(_02482_));
 AO32x1_ASAP7_75t_R _17807_ (.A1(_02476_),
    .A2(_09800_),
    .A3(_02481_),
    .B1(_02456_),
    .B2(_02482_),
    .Y(_01783_));
 NOR2x1_ASAP7_75t_R _17808_ (.A(_09804_),
    .B(_02456_),
    .Y(_02483_));
 INVx1_ASAP7_75t_R _17809_ (.A(_00227_),
    .Y(_02484_));
 AO32x1_ASAP7_75t_R _17810_ (.A1(_02476_),
    .A2(_09803_),
    .A3(_02483_),
    .B1(_02456_),
    .B2(_02484_),
    .Y(_01784_));
 INVx1_ASAP7_75t_R _17811_ (.A(_00193_),
    .Y(_02485_));
 AND2x2_ASAP7_75t_R _17812_ (.A(_09890_),
    .B(_02455_),
    .Y(_02486_));
 AO22x1_ASAP7_75t_R _17813_ (.A1(_02485_),
    .A2(_02450_),
    .B1(_02486_),
    .B2(_09808_),
    .Y(_01785_));
 AND4x1_ASAP7_75t_R _17814_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02454_),
    .Y(_02487_));
 INVx1_ASAP7_75t_R _17815_ (.A(_00160_),
    .Y(_02488_));
 AO32x1_ASAP7_75t_R _17816_ (.A1(_02476_),
    .A2(_09811_),
    .A3(_02487_),
    .B1(_02456_),
    .B2(_02488_),
    .Y(_01786_));
 AND3x1_ASAP7_75t_R _17817_ (.A(_09897_),
    .B(_09898_),
    .C(_02463_),
    .Y(_02489_));
 INVx1_ASAP7_75t_R _17818_ (.A(_00126_),
    .Y(_02490_));
 AO32x1_ASAP7_75t_R _17819_ (.A1(_02476_),
    .A2(_09813_),
    .A3(_02489_),
    .B1(_02456_),
    .B2(_02490_),
    .Y(_01787_));
 NAND2x1_ASAP7_75t_R _17820_ (.A(_01023_),
    .B(_02450_),
    .Y(_02491_));
 OA21x2_ASAP7_75t_R _17821_ (.A1(_09901_),
    .A2(_02448_),
    .B(_02491_),
    .Y(_01788_));
 AND4x1_ASAP7_75t_R _17822_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02454_),
    .Y(_02492_));
 INVx1_ASAP7_75t_R _17823_ (.A(_00092_),
    .Y(_02493_));
 AO32x1_ASAP7_75t_R _17824_ (.A1(_02476_),
    .A2(_09816_),
    .A3(_02492_),
    .B1(_02456_),
    .B2(_02493_),
    .Y(_01789_));
 AND3x1_ASAP7_75t_R _17825_ (.A(_09908_),
    .B(_09909_),
    .C(_02463_),
    .Y(_02494_));
 AO32x1_ASAP7_75t_R _17826_ (.A1(_02476_),
    .A2(_09818_),
    .A3(_02494_),
    .B1(_02456_),
    .B2(_04044_),
    .Y(_01790_));
 NAND2x1_ASAP7_75t_R _17827_ (.A(_00990_),
    .B(_02450_),
    .Y(_02495_));
 OA21x2_ASAP7_75t_R _17828_ (.A1(_09912_),
    .A2(_02448_),
    .B(_02495_),
    .Y(_01791_));
 NAND2x1_ASAP7_75t_R _17829_ (.A(_00957_),
    .B(_02450_),
    .Y(_02496_));
 OA21x2_ASAP7_75t_R _17830_ (.A1(_09914_),
    .A2(_02448_),
    .B(_02496_),
    .Y(_01792_));
 AND2x2_ASAP7_75t_R _17831_ (.A(_00923_),
    .B(_02456_),
    .Y(_02497_));
 AOI21x1_ASAP7_75t_R _17832_ (.A1(_09822_),
    .A2(_02455_),
    .B(_02497_),
    .Y(_01793_));
 NOR2x1_ASAP7_75t_R _17833_ (.A(_00890_),
    .B(_02455_),
    .Y(_02498_));
 AO21x1_ASAP7_75t_R _17834_ (.A1(_09917_),
    .A2(_02455_),
    .B(_02498_),
    .Y(_01794_));
 AND2x2_ASAP7_75t_R _17835_ (.A(_06528_),
    .B(_02456_),
    .Y(_02499_));
 AO21x1_ASAP7_75t_R _17836_ (.A1(_09919_),
    .A2(_02455_),
    .B(_02499_),
    .Y(_01795_));
 NOR2x1_ASAP7_75t_R _17837_ (.A(_00823_),
    .B(_02455_),
    .Y(_02500_));
 AO21x1_ASAP7_75t_R _17838_ (.A1(_09921_),
    .A2(_02455_),
    .B(_02500_),
    .Y(_01796_));
 NAND2x1_ASAP7_75t_R _17839_ (.A(_00789_),
    .B(_02462_),
    .Y(_02501_));
 OA21x2_ASAP7_75t_R _17840_ (.A1(_09923_),
    .A2(_02450_),
    .B(_02501_),
    .Y(_01797_));
 NAND2x2_ASAP7_75t_R _17841_ (.A(_08871_),
    .B(_02404_),
    .Y(_02502_));
 BUFx4f_ASAP7_75t_R _17842_ (.A(_02502_),
    .Y(_02503_));
 BUFx6f_ASAP7_75t_R _17843_ (.A(_02502_),
    .Y(_02504_));
 NAND2x1_ASAP7_75t_R _17844_ (.A(_00026_),
    .B(_02504_),
    .Y(_02505_));
 OA21x2_ASAP7_75t_R _17845_ (.A1(_09755_),
    .A2(_02503_),
    .B(_02505_),
    .Y(_01798_));
 NAND2x1_ASAP7_75t_R _17846_ (.A(_00758_),
    .B(_02504_),
    .Y(_02506_));
 OA21x2_ASAP7_75t_R _17847_ (.A1(_09835_),
    .A2(_02503_),
    .B(_02506_),
    .Y(_01799_));
 NAND2x1_ASAP7_75t_R _17848_ (.A(_00725_),
    .B(_02504_),
    .Y(_02507_));
 OA21x2_ASAP7_75t_R _17849_ (.A1(_09837_),
    .A2(_02503_),
    .B(_02507_),
    .Y(_01800_));
 NAND2x1_ASAP7_75t_R _17850_ (.A(_00692_),
    .B(_02504_),
    .Y(_02508_));
 OA21x2_ASAP7_75t_R _17851_ (.A1(_09839_),
    .A2(_02503_),
    .B(_02508_),
    .Y(_01801_));
 AND2x4_ASAP7_75t_R _17852_ (.A(_08602_),
    .B(_02401_),
    .Y(_02509_));
 BUFx6f_ASAP7_75t_R _17853_ (.A(_02509_),
    .Y(_02510_));
 BUFx6f_ASAP7_75t_R _17854_ (.A(_02502_),
    .Y(_02511_));
 AND2x2_ASAP7_75t_R _17855_ (.A(_00659_),
    .B(_02511_),
    .Y(_02512_));
 AOI21x1_ASAP7_75t_R _17856_ (.A1(_09763_),
    .A2(_02510_),
    .B(_02512_),
    .Y(_01802_));
 NAND2x1_ASAP7_75t_R _17857_ (.A(_00626_),
    .B(_02504_),
    .Y(_02513_));
 OA21x2_ASAP7_75t_R _17858_ (.A1(_09845_),
    .A2(_02503_),
    .B(_02513_),
    .Y(_01803_));
 AO21x1_ASAP7_75t_R _17859_ (.A1(_08871_),
    .A2(_02404_),
    .B(_00592_),
    .Y(_02514_));
 OAI21x1_ASAP7_75t_R _17860_ (.A1(_09937_),
    .A2(_02503_),
    .B(_02514_),
    .Y(_01804_));
 AND3x1_ASAP7_75t_R _17861_ (.A(_09848_),
    .B(_09849_),
    .C(_02510_),
    .Y(_02515_));
 BUFx10_ASAP7_75t_R _17862_ (.A(_02502_),
    .Y(_02516_));
 AO32x1_ASAP7_75t_R _17863_ (.A1(_09771_),
    .A2(_02460_),
    .A3(_02515_),
    .B1(_02516_),
    .B2(_05732_),
    .Y(_01805_));
 BUFx4f_ASAP7_75t_R _17864_ (.A(_02509_),
    .Y(_02517_));
 AND2x2_ASAP7_75t_R _17865_ (.A(_09854_),
    .B(_02517_),
    .Y(_02518_));
 INVx1_ASAP7_75t_R _17866_ (.A(_00526_),
    .Y(_02519_));
 AO32x1_ASAP7_75t_R _17867_ (.A1(_02476_),
    .A2(_09776_),
    .A3(_02518_),
    .B1(_02516_),
    .B2(_02519_),
    .Y(_01806_));
 AND3x1_ASAP7_75t_R _17868_ (.A(_09857_),
    .B(_09858_),
    .C(_02517_),
    .Y(_02520_));
 INVx1_ASAP7_75t_R _17869_ (.A(_00493_),
    .Y(_02521_));
 AO32x1_ASAP7_75t_R _17870_ (.A1(_02476_),
    .A2(_09779_),
    .A3(_02520_),
    .B1(_02516_),
    .B2(_02521_),
    .Y(_01807_));
 BUFx4f_ASAP7_75t_R _17871_ (.A(_09809_),
    .Y(_02522_));
 AND3x1_ASAP7_75t_R _17872_ (.A(_09861_),
    .B(_09862_),
    .C(_02517_),
    .Y(_02523_));
 INVx1_ASAP7_75t_R _17873_ (.A(_00460_),
    .Y(_02524_));
 AO32x1_ASAP7_75t_R _17874_ (.A1(_02522_),
    .A2(_09782_),
    .A3(_02523_),
    .B1(_02516_),
    .B2(_02524_),
    .Y(_01808_));
 NAND2x1_ASAP7_75t_R _17875_ (.A(_01057_),
    .B(_02504_),
    .Y(_02525_));
 OA21x2_ASAP7_75t_R _17876_ (.A1(_09865_),
    .A2(_02503_),
    .B(_02525_),
    .Y(_01809_));
 AND2x2_ASAP7_75t_R _17877_ (.A(_09867_),
    .B(_02517_),
    .Y(_02526_));
 INVx1_ASAP7_75t_R _17878_ (.A(_00427_),
    .Y(_02527_));
 AO32x1_ASAP7_75t_R _17879_ (.A1(_02522_),
    .A2(_09786_),
    .A3(_02526_),
    .B1(_02516_),
    .B2(_02527_),
    .Y(_01810_));
 AND3x1_ASAP7_75t_R _17880_ (.A(_09870_),
    .B(_09871_),
    .C(_02517_),
    .Y(_02528_));
 INVx1_ASAP7_75t_R _17881_ (.A(_00394_),
    .Y(_02529_));
 AO32x1_ASAP7_75t_R _17882_ (.A1(_02522_),
    .A2(_09789_),
    .A3(_02528_),
    .B1(_02516_),
    .B2(_02529_),
    .Y(_01811_));
 AND2x2_ASAP7_75t_R _17883_ (.A(_09874_),
    .B(_02517_),
    .Y(_02530_));
 INVx1_ASAP7_75t_R _17884_ (.A(_00361_),
    .Y(_02531_));
 AO32x1_ASAP7_75t_R _17885_ (.A1(_02522_),
    .A2(_09792_),
    .A3(_02530_),
    .B1(_02516_),
    .B2(_02531_),
    .Y(_01812_));
 AND2x2_ASAP7_75t_R _17886_ (.A(_09878_),
    .B(_02517_),
    .Y(_02532_));
 INVx1_ASAP7_75t_R _17887_ (.A(_00327_),
    .Y(_02533_));
 AO32x1_ASAP7_75t_R _17888_ (.A1(_02522_),
    .A2(_09794_),
    .A3(_02532_),
    .B1(_02516_),
    .B2(_02533_),
    .Y(_01813_));
 AND2x2_ASAP7_75t_R _17889_ (.A(_09881_),
    .B(_02517_),
    .Y(_02534_));
 AO32x1_ASAP7_75t_R _17890_ (.A1(_02522_),
    .A2(_09797_),
    .A3(_02534_),
    .B1(_02511_),
    .B2(_04890_),
    .Y(_01814_));
 AND2x2_ASAP7_75t_R _17891_ (.A(_09884_),
    .B(_02509_),
    .Y(_02535_));
 INVx1_ASAP7_75t_R _17892_ (.A(_00261_),
    .Y(_02536_));
 AO32x1_ASAP7_75t_R _17893_ (.A1(_02522_),
    .A2(_09800_),
    .A3(_02535_),
    .B1(_02511_),
    .B2(_02536_),
    .Y(_01815_));
 NOR2x1_ASAP7_75t_R _17894_ (.A(_09804_),
    .B(_02511_),
    .Y(_02537_));
 INVx1_ASAP7_75t_R _17895_ (.A(_00228_),
    .Y(_02538_));
 AO32x1_ASAP7_75t_R _17896_ (.A1(_02522_),
    .A2(_09803_),
    .A3(_02537_),
    .B1(_02511_),
    .B2(_02538_),
    .Y(_01816_));
 INVx1_ASAP7_75t_R _17897_ (.A(_00194_),
    .Y(_02539_));
 AND2x2_ASAP7_75t_R _17898_ (.A(_09890_),
    .B(_02510_),
    .Y(_02540_));
 AO22x1_ASAP7_75t_R _17899_ (.A1(_02539_),
    .A2(_02504_),
    .B1(_02540_),
    .B2(_09808_),
    .Y(_01817_));
 AND4x1_ASAP7_75t_R _17900_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02509_),
    .Y(_02541_));
 INVx1_ASAP7_75t_R _17901_ (.A(_00161_),
    .Y(_02542_));
 AO32x1_ASAP7_75t_R _17902_ (.A1(_02522_),
    .A2(_09811_),
    .A3(_02541_),
    .B1(_02511_),
    .B2(_02542_),
    .Y(_01818_));
 AND3x1_ASAP7_75t_R _17903_ (.A(_09897_),
    .B(_09898_),
    .C(_02517_),
    .Y(_02543_));
 INVx1_ASAP7_75t_R _17904_ (.A(_00127_),
    .Y(_02544_));
 AO32x1_ASAP7_75t_R _17905_ (.A1(_02522_),
    .A2(_09813_),
    .A3(_02543_),
    .B1(_02511_),
    .B2(_02544_),
    .Y(_01819_));
 NAND2x1_ASAP7_75t_R _17906_ (.A(_01024_),
    .B(_02504_),
    .Y(_02545_));
 OA21x2_ASAP7_75t_R _17907_ (.A1(_09901_),
    .A2(_02503_),
    .B(_02545_),
    .Y(_01820_));
 BUFx10_ASAP7_75t_R _17908_ (.A(_08784_),
    .Y(_02546_));
 BUFx4f_ASAP7_75t_R _17909_ (.A(_02546_),
    .Y(_02547_));
 AND4x1_ASAP7_75t_R _17910_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02509_),
    .Y(_02548_));
 INVx1_ASAP7_75t_R _17911_ (.A(_00093_),
    .Y(_02549_));
 AO32x1_ASAP7_75t_R _17912_ (.A1(_02547_),
    .A2(_09816_),
    .A3(_02548_),
    .B1(_02511_),
    .B2(_02549_),
    .Y(_01821_));
 AND3x1_ASAP7_75t_R _17913_ (.A(_09908_),
    .B(_09909_),
    .C(_02517_),
    .Y(_02550_));
 INVx1_ASAP7_75t_R _17914_ (.A(_00061_),
    .Y(_02551_));
 AO32x1_ASAP7_75t_R _17915_ (.A1(_02547_),
    .A2(_09818_),
    .A3(_02550_),
    .B1(_02511_),
    .B2(_02551_),
    .Y(_01822_));
 NAND2x1_ASAP7_75t_R _17916_ (.A(_00991_),
    .B(_02504_),
    .Y(_02552_));
 OA21x2_ASAP7_75t_R _17917_ (.A1(_09912_),
    .A2(_02503_),
    .B(_02552_),
    .Y(_01823_));
 NAND2x1_ASAP7_75t_R _17918_ (.A(_00958_),
    .B(_02516_),
    .Y(_02553_));
 OA21x2_ASAP7_75t_R _17919_ (.A1(_09914_),
    .A2(_02503_),
    .B(_02553_),
    .Y(_01824_));
 AND2x2_ASAP7_75t_R _17920_ (.A(_00924_),
    .B(_02511_),
    .Y(_02554_));
 AOI21x1_ASAP7_75t_R _17921_ (.A1(_09822_),
    .A2(_02510_),
    .B(_02554_),
    .Y(_01825_));
 NOR2x1_ASAP7_75t_R _17922_ (.A(_00891_),
    .B(_02510_),
    .Y(_02555_));
 AO21x1_ASAP7_75t_R _17923_ (.A1(_09917_),
    .A2(_02510_),
    .B(_02555_),
    .Y(_01826_));
 NOR2x1_ASAP7_75t_R _17924_ (.A(_00857_),
    .B(_02510_),
    .Y(_02556_));
 AO21x1_ASAP7_75t_R _17925_ (.A1(_09919_),
    .A2(_02510_),
    .B(_02556_),
    .Y(_01827_));
 NOR2x1_ASAP7_75t_R _17926_ (.A(_00824_),
    .B(_02510_),
    .Y(_02557_));
 AO21x1_ASAP7_75t_R _17927_ (.A1(_09921_),
    .A2(_02510_),
    .B(_02557_),
    .Y(_01828_));
 NAND2x1_ASAP7_75t_R _17928_ (.A(_00790_),
    .B(_02516_),
    .Y(_02558_));
 OA21x2_ASAP7_75t_R _17929_ (.A1(_09923_),
    .A2(_02504_),
    .B(_02558_),
    .Y(_01829_));
 NAND2x2_ASAP7_75t_R _17930_ (.A(_09191_),
    .B(_02401_),
    .Y(_02559_));
 BUFx4f_ASAP7_75t_R _17931_ (.A(_02559_),
    .Y(_02560_));
 BUFx6f_ASAP7_75t_R _17932_ (.A(_02559_),
    .Y(_02561_));
 NAND2x1_ASAP7_75t_R _17933_ (.A(_00027_),
    .B(_02561_),
    .Y(_02562_));
 OA21x2_ASAP7_75t_R _17934_ (.A1(_09755_),
    .A2(_02560_),
    .B(_02562_),
    .Y(_01830_));
 NAND2x1_ASAP7_75t_R _17935_ (.A(_00759_),
    .B(_02561_),
    .Y(_02563_));
 OA21x2_ASAP7_75t_R _17936_ (.A1(_09835_),
    .A2(_02560_),
    .B(_02563_),
    .Y(_01831_));
 NAND2x1_ASAP7_75t_R _17937_ (.A(_00726_),
    .B(_02561_),
    .Y(_02564_));
 OA21x2_ASAP7_75t_R _17938_ (.A1(_09837_),
    .A2(_02560_),
    .B(_02564_),
    .Y(_01832_));
 NAND2x1_ASAP7_75t_R _17939_ (.A(_00693_),
    .B(_02561_),
    .Y(_02565_));
 OA21x2_ASAP7_75t_R _17940_ (.A1(_09839_),
    .A2(_02560_),
    .B(_02565_),
    .Y(_01833_));
 AND2x6_ASAP7_75t_R _17941_ (.A(_09190_),
    .B(_02401_),
    .Y(_02566_));
 BUFx6f_ASAP7_75t_R _17942_ (.A(_02566_),
    .Y(_02567_));
 BUFx6f_ASAP7_75t_R _17943_ (.A(_02559_),
    .Y(_02568_));
 AND2x2_ASAP7_75t_R _17944_ (.A(_00660_),
    .B(_02568_),
    .Y(_02569_));
 AOI21x1_ASAP7_75t_R _17945_ (.A1(_09763_),
    .A2(_02567_),
    .B(_02569_),
    .Y(_01834_));
 NAND2x1_ASAP7_75t_R _17946_ (.A(_00627_),
    .B(_02561_),
    .Y(_02570_));
 OA21x2_ASAP7_75t_R _17947_ (.A1(_09845_),
    .A2(_02560_),
    .B(_02570_),
    .Y(_01835_));
 AND2x2_ASAP7_75t_R _17948_ (.A(_00593_),
    .B(_02568_),
    .Y(_02571_));
 AOI21x1_ASAP7_75t_R _17949_ (.A1(_09769_),
    .A2(_02567_),
    .B(_02571_),
    .Y(_01836_));
 BUFx4f_ASAP7_75t_R _17950_ (.A(_02566_),
    .Y(_02572_));
 AND3x1_ASAP7_75t_R _17951_ (.A(_09848_),
    .B(_09849_),
    .C(_02572_),
    .Y(_02573_));
 BUFx6f_ASAP7_75t_R _17952_ (.A(_02559_),
    .Y(_02574_));
 AO32x1_ASAP7_75t_R _17953_ (.A1(_09771_),
    .A2(_02460_),
    .A3(_02573_),
    .B1(_02574_),
    .B2(_05655_),
    .Y(_01837_));
 AND2x2_ASAP7_75t_R _17954_ (.A(_09854_),
    .B(_02572_),
    .Y(_02575_));
 INVx1_ASAP7_75t_R _17955_ (.A(_00527_),
    .Y(_02576_));
 AO32x1_ASAP7_75t_R _17956_ (.A1(_02547_),
    .A2(_09776_),
    .A3(_02575_),
    .B1(_02574_),
    .B2(_02576_),
    .Y(_01838_));
 AND3x1_ASAP7_75t_R _17957_ (.A(_09857_),
    .B(_09858_),
    .C(_02572_),
    .Y(_02577_));
 INVx1_ASAP7_75t_R _17958_ (.A(_00494_),
    .Y(_02578_));
 AO32x1_ASAP7_75t_R _17959_ (.A1(_02547_),
    .A2(_09779_),
    .A3(_02577_),
    .B1(_02574_),
    .B2(_02578_),
    .Y(_01839_));
 AND3x1_ASAP7_75t_R _17960_ (.A(_09861_),
    .B(_09862_),
    .C(_02572_),
    .Y(_02579_));
 INVx1_ASAP7_75t_R _17961_ (.A(_00461_),
    .Y(_02580_));
 AO32x1_ASAP7_75t_R _17962_ (.A1(_02547_),
    .A2(_09782_),
    .A3(_02579_),
    .B1(_02574_),
    .B2(_02580_),
    .Y(_01840_));
 NAND2x1_ASAP7_75t_R _17963_ (.A(_01058_),
    .B(_02561_),
    .Y(_02581_));
 OA21x2_ASAP7_75t_R _17964_ (.A1(_09865_),
    .A2(_02560_),
    .B(_02581_),
    .Y(_01841_));
 AND2x2_ASAP7_75t_R _17965_ (.A(_09867_),
    .B(_02572_),
    .Y(_02582_));
 INVx1_ASAP7_75t_R _17966_ (.A(_00428_),
    .Y(_02583_));
 AO32x1_ASAP7_75t_R _17967_ (.A1(_02547_),
    .A2(_09786_),
    .A3(_02582_),
    .B1(_02574_),
    .B2(_02583_),
    .Y(_01842_));
 AND3x1_ASAP7_75t_R _17968_ (.A(_09870_),
    .B(_09871_),
    .C(_02572_),
    .Y(_02584_));
 AO32x1_ASAP7_75t_R _17969_ (.A1(_02547_),
    .A2(_09789_),
    .A3(_02584_),
    .B1(_02574_),
    .B2(_05170_),
    .Y(_01843_));
 AND2x2_ASAP7_75t_R _17970_ (.A(_09874_),
    .B(_02572_),
    .Y(_02585_));
 INVx1_ASAP7_75t_R _17971_ (.A(_00362_),
    .Y(_02586_));
 AO32x1_ASAP7_75t_R _17972_ (.A1(_02547_),
    .A2(_09792_),
    .A3(_02585_),
    .B1(_02574_),
    .B2(_02586_),
    .Y(_01844_));
 AND2x2_ASAP7_75t_R _17973_ (.A(_09878_),
    .B(_02572_),
    .Y(_02587_));
 INVx1_ASAP7_75t_R _17974_ (.A(_00328_),
    .Y(_02588_));
 AO32x1_ASAP7_75t_R _17975_ (.A1(_02547_),
    .A2(_09794_),
    .A3(_02587_),
    .B1(_02574_),
    .B2(_02588_),
    .Y(_01845_));
 AND2x2_ASAP7_75t_R _17976_ (.A(_09881_),
    .B(_02566_),
    .Y(_02589_));
 AO32x1_ASAP7_75t_R _17977_ (.A1(_02547_),
    .A2(_09797_),
    .A3(_02589_),
    .B1(_02574_),
    .B2(_04898_),
    .Y(_01846_));
 BUFx4f_ASAP7_75t_R _17978_ (.A(_02546_),
    .Y(_02590_));
 AND2x2_ASAP7_75t_R _17979_ (.A(_09884_),
    .B(_02566_),
    .Y(_02591_));
 INVx1_ASAP7_75t_R _17980_ (.A(_00262_),
    .Y(_02592_));
 AO32x1_ASAP7_75t_R _17981_ (.A1(_02590_),
    .A2(_09800_),
    .A3(_02591_),
    .B1(_02568_),
    .B2(_02592_),
    .Y(_01847_));
 NOR2x1_ASAP7_75t_R _17982_ (.A(_09804_),
    .B(_02568_),
    .Y(_02593_));
 INVx1_ASAP7_75t_R _17983_ (.A(_00229_),
    .Y(_02594_));
 AO32x1_ASAP7_75t_R _17984_ (.A1(_02590_),
    .A2(_09803_),
    .A3(_02593_),
    .B1(_02568_),
    .B2(_02594_),
    .Y(_01848_));
 INVx1_ASAP7_75t_R _17985_ (.A(_00195_),
    .Y(_02595_));
 AND2x2_ASAP7_75t_R _17986_ (.A(_09890_),
    .B(_02567_),
    .Y(_02596_));
 AO22x1_ASAP7_75t_R _17987_ (.A1(_02595_),
    .A2(_02561_),
    .B1(_02596_),
    .B2(_09808_),
    .Y(_01849_));
 AND4x1_ASAP7_75t_R _17988_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02566_),
    .Y(_02597_));
 INVx1_ASAP7_75t_R _17989_ (.A(_00162_),
    .Y(_02598_));
 AO32x1_ASAP7_75t_R _17990_ (.A1(_02590_),
    .A2(_09811_),
    .A3(_02597_),
    .B1(_02568_),
    .B2(_02598_),
    .Y(_01850_));
 AND3x1_ASAP7_75t_R _17991_ (.A(_09897_),
    .B(_09898_),
    .C(_02572_),
    .Y(_02599_));
 INVx1_ASAP7_75t_R _17992_ (.A(_00128_),
    .Y(_02600_));
 AO32x1_ASAP7_75t_R _17993_ (.A1(_02590_),
    .A2(_09813_),
    .A3(_02599_),
    .B1(_02568_),
    .B2(_02600_),
    .Y(_01851_));
 NAND2x1_ASAP7_75t_R _17994_ (.A(_01025_),
    .B(_02561_),
    .Y(_02601_));
 OA21x2_ASAP7_75t_R _17995_ (.A1(_09901_),
    .A2(_02560_),
    .B(_02601_),
    .Y(_01852_));
 AND4x1_ASAP7_75t_R _17996_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02566_),
    .Y(_02602_));
 INVx1_ASAP7_75t_R _17997_ (.A(_00094_),
    .Y(_02603_));
 AO32x1_ASAP7_75t_R _17998_ (.A1(_02590_),
    .A2(_09816_),
    .A3(_02602_),
    .B1(_02568_),
    .B2(_02603_),
    .Y(_01853_));
 AND3x1_ASAP7_75t_R _17999_ (.A(_09908_),
    .B(_09909_),
    .C(_02572_),
    .Y(_02604_));
 INVx1_ASAP7_75t_R _18000_ (.A(_00062_),
    .Y(_02605_));
 AO32x1_ASAP7_75t_R _18001_ (.A1(_02590_),
    .A2(_09818_),
    .A3(_02604_),
    .B1(_02568_),
    .B2(_02605_),
    .Y(_01854_));
 NAND2x1_ASAP7_75t_R _18002_ (.A(_00992_),
    .B(_02561_),
    .Y(_02606_));
 OA21x2_ASAP7_75t_R _18003_ (.A1(_09912_),
    .A2(_02560_),
    .B(_02606_),
    .Y(_01855_));
 NAND2x1_ASAP7_75t_R _18004_ (.A(_00959_),
    .B(_02561_),
    .Y(_02607_));
 OA21x2_ASAP7_75t_R _18005_ (.A1(_09914_),
    .A2(_02560_),
    .B(_02607_),
    .Y(_01856_));
 AND2x2_ASAP7_75t_R _18006_ (.A(_00925_),
    .B(_02568_),
    .Y(_02608_));
 AOI21x1_ASAP7_75t_R _18007_ (.A1(_09822_),
    .A2(_02567_),
    .B(_02608_),
    .Y(_01857_));
 NOR2x1_ASAP7_75t_R _18008_ (.A(_00892_),
    .B(_02567_),
    .Y(_02609_));
 AO21x1_ASAP7_75t_R _18009_ (.A1(_09917_),
    .A2(_02567_),
    .B(_02609_),
    .Y(_01858_));
 NOR2x1_ASAP7_75t_R _18010_ (.A(_00858_),
    .B(_02567_),
    .Y(_02610_));
 AO21x1_ASAP7_75t_R _18011_ (.A1(_09919_),
    .A2(_02567_),
    .B(_02610_),
    .Y(_01859_));
 NOR2x1_ASAP7_75t_R _18012_ (.A(_00825_),
    .B(_02567_),
    .Y(_02611_));
 AO21x1_ASAP7_75t_R _18013_ (.A1(_09921_),
    .A2(_02567_),
    .B(_02611_),
    .Y(_01860_));
 NAND2x1_ASAP7_75t_R _18014_ (.A(_00791_),
    .B(_02574_),
    .Y(_02612_));
 OA21x2_ASAP7_75t_R _18015_ (.A1(_09923_),
    .A2(_02560_),
    .B(_02612_),
    .Y(_01861_));
 AND3x4_ASAP7_75t_R _18016_ (.A(net2),
    .B(_06807_),
    .C(_08603_),
    .Y(_02613_));
 BUFx12f_ASAP7_75t_R _18017_ (.A(_02613_),
    .Y(_02614_));
 NAND2x2_ASAP7_75t_R _18018_ (.A(_09528_),
    .B(_02614_),
    .Y(_02615_));
 BUFx10_ASAP7_75t_R _18019_ (.A(_02615_),
    .Y(_02616_));
 BUFx4f_ASAP7_75t_R _18020_ (.A(_02616_),
    .Y(_02617_));
 AO21x1_ASAP7_75t_R _18021_ (.A1(_09529_),
    .A2(_02614_),
    .B(_03436_),
    .Y(_02618_));
 OA21x2_ASAP7_75t_R _18022_ (.A1(_09755_),
    .A2(_02617_),
    .B(_02618_),
    .Y(_01862_));
 BUFx10_ASAP7_75t_R _18023_ (.A(_02615_),
    .Y(_02619_));
 NAND2x1_ASAP7_75t_R _18024_ (.A(_00760_),
    .B(_02619_),
    .Y(_02620_));
 OA21x2_ASAP7_75t_R _18025_ (.A1(_09835_),
    .A2(_02617_),
    .B(_02620_),
    .Y(_01863_));
 NAND2x1_ASAP7_75t_R _18026_ (.A(_00727_),
    .B(_02619_),
    .Y(_02621_));
 OA21x2_ASAP7_75t_R _18027_ (.A1(_09837_),
    .A2(_02617_),
    .B(_02621_),
    .Y(_01864_));
 NAND2x1_ASAP7_75t_R _18028_ (.A(_00694_),
    .B(_02619_),
    .Y(_02622_));
 OA21x2_ASAP7_75t_R _18029_ (.A1(_09839_),
    .A2(_02617_),
    .B(_02622_),
    .Y(_01865_));
 AND2x6_ASAP7_75t_R _18030_ (.A(_09528_),
    .B(_02613_),
    .Y(_02623_));
 BUFx6f_ASAP7_75t_R _18031_ (.A(_02623_),
    .Y(_02624_));
 AND2x2_ASAP7_75t_R _18032_ (.A(_00661_),
    .B(_02616_),
    .Y(_02625_));
 AOI21x1_ASAP7_75t_R _18033_ (.A1(_09763_),
    .A2(_02624_),
    .B(_02625_),
    .Y(_01866_));
 NAND2x1_ASAP7_75t_R _18034_ (.A(_00628_),
    .B(_02619_),
    .Y(_02626_));
 OA21x2_ASAP7_75t_R _18035_ (.A1(_09845_),
    .A2(_02617_),
    .B(_02626_),
    .Y(_01867_));
 AND2x2_ASAP7_75t_R _18036_ (.A(_00594_),
    .B(_02616_),
    .Y(_02627_));
 AOI21x1_ASAP7_75t_R _18037_ (.A1(_09769_),
    .A2(_02624_),
    .B(_02627_),
    .Y(_01868_));
 BUFx4f_ASAP7_75t_R _18038_ (.A(_02623_),
    .Y(_02628_));
 AND3x1_ASAP7_75t_R _18039_ (.A(_09848_),
    .B(_09849_),
    .C(_02628_),
    .Y(_02629_));
 BUFx6f_ASAP7_75t_R _18040_ (.A(_02615_),
    .Y(_02630_));
 INVx1_ASAP7_75t_R _18041_ (.A(_00561_),
    .Y(_02631_));
 AO32x1_ASAP7_75t_R _18042_ (.A1(_09771_),
    .A2(_02460_),
    .A3(_02629_),
    .B1(_02630_),
    .B2(_02631_),
    .Y(_01869_));
 AND2x2_ASAP7_75t_R _18043_ (.A(_09854_),
    .B(_02628_),
    .Y(_02632_));
 INVx1_ASAP7_75t_R _18044_ (.A(_00528_),
    .Y(_02633_));
 AO32x1_ASAP7_75t_R _18045_ (.A1(_02590_),
    .A2(_09776_),
    .A3(_02632_),
    .B1(_02630_),
    .B2(_02633_),
    .Y(_01870_));
 AND3x1_ASAP7_75t_R _18046_ (.A(_09857_),
    .B(_09858_),
    .C(_02628_),
    .Y(_02634_));
 INVx1_ASAP7_75t_R _18047_ (.A(_00495_),
    .Y(_02635_));
 AO32x1_ASAP7_75t_R _18048_ (.A1(_02590_),
    .A2(_09779_),
    .A3(_02634_),
    .B1(_02630_),
    .B2(_02635_),
    .Y(_01871_));
 AND3x1_ASAP7_75t_R _18049_ (.A(_09861_),
    .B(_09862_),
    .C(_02628_),
    .Y(_02636_));
 INVx1_ASAP7_75t_R _18050_ (.A(_00462_),
    .Y(_02637_));
 AO32x1_ASAP7_75t_R _18051_ (.A1(_02590_),
    .A2(_09782_),
    .A3(_02636_),
    .B1(_02630_),
    .B2(_02637_),
    .Y(_01872_));
 NAND2x1_ASAP7_75t_R _18052_ (.A(_01059_),
    .B(_02619_),
    .Y(_02638_));
 OA21x2_ASAP7_75t_R _18053_ (.A1(_09865_),
    .A2(_02617_),
    .B(_02638_),
    .Y(_01873_));
 AND2x2_ASAP7_75t_R _18054_ (.A(_09867_),
    .B(_02628_),
    .Y(_02639_));
 INVx1_ASAP7_75t_R _18055_ (.A(_00429_),
    .Y(_02640_));
 AO32x1_ASAP7_75t_R _18056_ (.A1(_02590_),
    .A2(_09786_),
    .A3(_02639_),
    .B1(_02630_),
    .B2(_02640_),
    .Y(_01874_));
 BUFx4f_ASAP7_75t_R _18057_ (.A(_02546_),
    .Y(_02641_));
 AND3x1_ASAP7_75t_R _18058_ (.A(_09870_),
    .B(_09871_),
    .C(_02628_),
    .Y(_02642_));
 INVx1_ASAP7_75t_R _18059_ (.A(_00396_),
    .Y(_02643_));
 AO32x1_ASAP7_75t_R _18060_ (.A1(_02641_),
    .A2(_09789_),
    .A3(_02642_),
    .B1(_02630_),
    .B2(_02643_),
    .Y(_01875_));
 AND2x2_ASAP7_75t_R _18061_ (.A(_09874_),
    .B(_02628_),
    .Y(_02644_));
 INVx1_ASAP7_75t_R _18062_ (.A(_00363_),
    .Y(_02645_));
 AO32x1_ASAP7_75t_R _18063_ (.A1(_02641_),
    .A2(_09792_),
    .A3(_02644_),
    .B1(_02630_),
    .B2(_02645_),
    .Y(_01876_));
 AND2x2_ASAP7_75t_R _18064_ (.A(_09878_),
    .B(_02628_),
    .Y(_02646_));
 INVx1_ASAP7_75t_R _18065_ (.A(_00329_),
    .Y(_02647_));
 AO32x1_ASAP7_75t_R _18066_ (.A1(_02641_),
    .A2(_09794_),
    .A3(_02646_),
    .B1(_02630_),
    .B2(_02647_),
    .Y(_01877_));
 AND2x2_ASAP7_75t_R _18067_ (.A(_09881_),
    .B(_02623_),
    .Y(_02648_));
 INVx1_ASAP7_75t_R _18068_ (.A(_00296_),
    .Y(_02649_));
 AO32x1_ASAP7_75t_R _18069_ (.A1(_02641_),
    .A2(_09797_),
    .A3(_02648_),
    .B1(_02630_),
    .B2(_02649_),
    .Y(_01878_));
 AND2x2_ASAP7_75t_R _18070_ (.A(_09884_),
    .B(_02623_),
    .Y(_02650_));
 INVx1_ASAP7_75t_R _18071_ (.A(_00263_),
    .Y(_02651_));
 AO32x1_ASAP7_75t_R _18072_ (.A1(_02641_),
    .A2(_09800_),
    .A3(_02650_),
    .B1(_02630_),
    .B2(_02651_),
    .Y(_01879_));
 NOR2x1_ASAP7_75t_R _18073_ (.A(_09804_),
    .B(_02616_),
    .Y(_02652_));
 INVx1_ASAP7_75t_R _18074_ (.A(_00230_),
    .Y(_02653_));
 AO32x1_ASAP7_75t_R _18075_ (.A1(_02641_),
    .A2(_09803_),
    .A3(_02652_),
    .B1(_02616_),
    .B2(_02653_),
    .Y(_01880_));
 INVx1_ASAP7_75t_R _18076_ (.A(_00196_),
    .Y(_02654_));
 AND2x2_ASAP7_75t_R _18077_ (.A(_09890_),
    .B(_02624_),
    .Y(_02655_));
 AO22x1_ASAP7_75t_R _18078_ (.A1(_02654_),
    .A2(_02619_),
    .B1(_02655_),
    .B2(_09808_),
    .Y(_01881_));
 AND4x1_ASAP7_75t_R _18079_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02623_),
    .Y(_02656_));
 INVx1_ASAP7_75t_R _18080_ (.A(_00163_),
    .Y(_02657_));
 AO32x1_ASAP7_75t_R _18081_ (.A1(_02641_),
    .A2(_09811_),
    .A3(_02656_),
    .B1(_02616_),
    .B2(_02657_),
    .Y(_01882_));
 AND3x1_ASAP7_75t_R _18082_ (.A(_09897_),
    .B(_09898_),
    .C(_02628_),
    .Y(_02658_));
 INVx1_ASAP7_75t_R _18083_ (.A(_00129_),
    .Y(_02659_));
 AO32x1_ASAP7_75t_R _18084_ (.A1(_02641_),
    .A2(_09813_),
    .A3(_02658_),
    .B1(_02616_),
    .B2(_02659_),
    .Y(_01883_));
 NAND2x1_ASAP7_75t_R _18085_ (.A(_01026_),
    .B(_02619_),
    .Y(_02660_));
 OA21x2_ASAP7_75t_R _18086_ (.A1(_09901_),
    .A2(_02617_),
    .B(_02660_),
    .Y(_01884_));
 AND4x1_ASAP7_75t_R _18087_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02623_),
    .Y(_02661_));
 INVx1_ASAP7_75t_R _18088_ (.A(_00095_),
    .Y(_02662_));
 AO32x1_ASAP7_75t_R _18089_ (.A1(_02641_),
    .A2(_09816_),
    .A3(_02661_),
    .B1(_02616_),
    .B2(_02662_),
    .Y(_01885_));
 AND3x1_ASAP7_75t_R _18090_ (.A(_09908_),
    .B(_09909_),
    .C(_02628_),
    .Y(_02663_));
 INVx1_ASAP7_75t_R _18091_ (.A(_00063_),
    .Y(_02664_));
 AO32x1_ASAP7_75t_R _18092_ (.A1(_02641_),
    .A2(_09818_),
    .A3(_02663_),
    .B1(_02616_),
    .B2(_02664_),
    .Y(_01886_));
 NAND2x1_ASAP7_75t_R _18093_ (.A(_00993_),
    .B(_02619_),
    .Y(_02665_));
 OA21x2_ASAP7_75t_R _18094_ (.A1(_09912_),
    .A2(_02617_),
    .B(_02665_),
    .Y(_01887_));
 NAND2x1_ASAP7_75t_R _18095_ (.A(_00960_),
    .B(_02619_),
    .Y(_02666_));
 OA21x2_ASAP7_75t_R _18096_ (.A1(_09914_),
    .A2(_02617_),
    .B(_02666_),
    .Y(_01888_));
 AND2x2_ASAP7_75t_R _18097_ (.A(_00926_),
    .B(_02616_),
    .Y(_02667_));
 AOI21x1_ASAP7_75t_R _18098_ (.A1(_09822_),
    .A2(_02624_),
    .B(_02667_),
    .Y(_01889_));
 NOR2x1_ASAP7_75t_R _18099_ (.A(_00893_),
    .B(_02624_),
    .Y(_02668_));
 AO21x1_ASAP7_75t_R _18100_ (.A1(_09917_),
    .A2(_02624_),
    .B(_02668_),
    .Y(_01890_));
 NOR2x1_ASAP7_75t_R _18101_ (.A(_00859_),
    .B(_02624_),
    .Y(_02669_));
 AO21x1_ASAP7_75t_R _18102_ (.A1(_09919_),
    .A2(_02624_),
    .B(_02669_),
    .Y(_01891_));
 NOR2x1_ASAP7_75t_R _18103_ (.A(_00826_),
    .B(_02624_),
    .Y(_02670_));
 AO21x1_ASAP7_75t_R _18104_ (.A1(_09921_),
    .A2(_02624_),
    .B(_02670_),
    .Y(_01892_));
 NAND2x1_ASAP7_75t_R _18105_ (.A(_00792_),
    .B(_02619_),
    .Y(_02671_));
 OA21x2_ASAP7_75t_R _18106_ (.A1(_09923_),
    .A2(_02617_),
    .B(_02671_),
    .Y(_01893_));
 BUFx6f_ASAP7_75t_R _18107_ (.A(_08596_),
    .Y(_02672_));
 NAND2x2_ASAP7_75t_R _18108_ (.A(_09590_),
    .B(_02614_),
    .Y(_02673_));
 BUFx6f_ASAP7_75t_R _18109_ (.A(_02673_),
    .Y(_02674_));
 BUFx10_ASAP7_75t_R _18110_ (.A(_02674_),
    .Y(_02675_));
 INVx1_ASAP7_75t_R _18111_ (.A(_00029_),
    .Y(_02676_));
 AO21x1_ASAP7_75t_R _18112_ (.A1(_09597_),
    .A2(_02614_),
    .B(_02676_),
    .Y(_02677_));
 OA21x2_ASAP7_75t_R _18113_ (.A1(_02672_),
    .A2(_02675_),
    .B(_02677_),
    .Y(_01894_));
 BUFx12_ASAP7_75t_R _18114_ (.A(_02673_),
    .Y(_02678_));
 NAND2x1_ASAP7_75t_R _18115_ (.A(_00761_),
    .B(_02678_),
    .Y(_02679_));
 OA21x2_ASAP7_75t_R _18116_ (.A1(_09835_),
    .A2(_02675_),
    .B(_02679_),
    .Y(_01895_));
 NAND2x1_ASAP7_75t_R _18117_ (.A(_00728_),
    .B(_02678_),
    .Y(_02680_));
 OA21x2_ASAP7_75t_R _18118_ (.A1(_09837_),
    .A2(_02675_),
    .B(_02680_),
    .Y(_01896_));
 NAND2x1_ASAP7_75t_R _18119_ (.A(_00695_),
    .B(_02678_),
    .Y(_02681_));
 OA21x2_ASAP7_75t_R _18120_ (.A1(_09839_),
    .A2(_02675_),
    .B(_02681_),
    .Y(_01897_));
 BUFx12f_ASAP7_75t_R _18121_ (.A(_08724_),
    .Y(_02682_));
 AND2x4_ASAP7_75t_R _18122_ (.A(_09589_),
    .B(_02613_),
    .Y(_02683_));
 BUFx10_ASAP7_75t_R _18123_ (.A(_02683_),
    .Y(_02684_));
 AND2x2_ASAP7_75t_R _18124_ (.A(_00662_),
    .B(_02674_),
    .Y(_02685_));
 AOI21x1_ASAP7_75t_R _18125_ (.A1(_02682_),
    .A2(_02684_),
    .B(_02685_),
    .Y(_01898_));
 NAND2x1_ASAP7_75t_R _18126_ (.A(_00629_),
    .B(_02678_),
    .Y(_02686_));
 OA21x2_ASAP7_75t_R _18127_ (.A1(_09845_),
    .A2(_02675_),
    .B(_02686_),
    .Y(_01899_));
 AO21x1_ASAP7_75t_R _18128_ (.A1(_09597_),
    .A2(_02614_),
    .B(_00595_),
    .Y(_02687_));
 OAI21x1_ASAP7_75t_R _18129_ (.A1(_09937_),
    .A2(_02675_),
    .B(_02687_),
    .Y(_01900_));
 BUFx6f_ASAP7_75t_R _18130_ (.A(_08782_),
    .Y(_02688_));
 AND3x1_ASAP7_75t_R _18131_ (.A(_09848_),
    .B(_09849_),
    .C(_02684_),
    .Y(_02689_));
 BUFx10_ASAP7_75t_R _18132_ (.A(_02673_),
    .Y(_02690_));
 INVx1_ASAP7_75t_R _18133_ (.A(_00562_),
    .Y(_02691_));
 AO32x1_ASAP7_75t_R _18134_ (.A1(_02688_),
    .A2(_02460_),
    .A3(_02689_),
    .B1(_02690_),
    .B2(_02691_),
    .Y(_01901_));
 BUFx4f_ASAP7_75t_R _18135_ (.A(_02546_),
    .Y(_02692_));
 BUFx6f_ASAP7_75t_R _18136_ (.A(_08804_),
    .Y(_02693_));
 BUFx3_ASAP7_75t_R _18137_ (.A(_02683_),
    .Y(_02694_));
 AND2x2_ASAP7_75t_R _18138_ (.A(_09854_),
    .B(_02694_),
    .Y(_02695_));
 INVx1_ASAP7_75t_R _18139_ (.A(_00529_),
    .Y(_02696_));
 AO32x1_ASAP7_75t_R _18140_ (.A1(_02692_),
    .A2(_02693_),
    .A3(_02695_),
    .B1(_02690_),
    .B2(_02696_),
    .Y(_01902_));
 BUFx4f_ASAP7_75t_R _18141_ (.A(_08829_),
    .Y(_02697_));
 AND3x1_ASAP7_75t_R _18142_ (.A(_09857_),
    .B(_09858_),
    .C(_02694_),
    .Y(_02698_));
 INVx1_ASAP7_75t_R _18143_ (.A(_00496_),
    .Y(_02699_));
 AO32x1_ASAP7_75t_R _18144_ (.A1(_02692_),
    .A2(_02697_),
    .A3(_02698_),
    .B1(_02690_),
    .B2(_02699_),
    .Y(_01903_));
 BUFx4f_ASAP7_75t_R _18145_ (.A(_08849_),
    .Y(_02700_));
 AND3x1_ASAP7_75t_R _18146_ (.A(_09861_),
    .B(_09862_),
    .C(_02694_),
    .Y(_02701_));
 INVx1_ASAP7_75t_R _18147_ (.A(_00463_),
    .Y(_02702_));
 AO32x1_ASAP7_75t_R _18148_ (.A1(_02692_),
    .A2(_02700_),
    .A3(_02701_),
    .B1(_02690_),
    .B2(_02702_),
    .Y(_01904_));
 NAND2x1_ASAP7_75t_R _18149_ (.A(_01060_),
    .B(_02678_),
    .Y(_02703_));
 OA21x2_ASAP7_75t_R _18150_ (.A1(_09865_),
    .A2(_02675_),
    .B(_02703_),
    .Y(_01905_));
 BUFx6f_ASAP7_75t_R _18151_ (.A(_08878_),
    .Y(_02704_));
 AND2x2_ASAP7_75t_R _18152_ (.A(_09867_),
    .B(_02694_),
    .Y(_02705_));
 INVx1_ASAP7_75t_R _18153_ (.A(_00430_),
    .Y(_02706_));
 AO32x1_ASAP7_75t_R _18154_ (.A1(_02692_),
    .A2(_02704_),
    .A3(_02705_),
    .B1(_02690_),
    .B2(_02706_),
    .Y(_01906_));
 BUFx6f_ASAP7_75t_R _18155_ (.A(_08900_),
    .Y(_02707_));
 AND3x1_ASAP7_75t_R _18156_ (.A(_09870_),
    .B(_09871_),
    .C(_02694_),
    .Y(_02708_));
 INVx1_ASAP7_75t_R _18157_ (.A(_00397_),
    .Y(_02709_));
 AO32x1_ASAP7_75t_R _18158_ (.A1(_02692_),
    .A2(_02707_),
    .A3(_02708_),
    .B1(_02690_),
    .B2(_02709_),
    .Y(_01907_));
 BUFx4f_ASAP7_75t_R _18159_ (.A(_08917_),
    .Y(_02710_));
 AND2x2_ASAP7_75t_R _18160_ (.A(_09874_),
    .B(_02694_),
    .Y(_02711_));
 INVx1_ASAP7_75t_R _18161_ (.A(_00364_),
    .Y(_02712_));
 AO32x1_ASAP7_75t_R _18162_ (.A1(_02692_),
    .A2(_02710_),
    .A3(_02711_),
    .B1(_02690_),
    .B2(_02712_),
    .Y(_01908_));
 BUFx6f_ASAP7_75t_R _18163_ (.A(_08936_),
    .Y(_02713_));
 AND2x2_ASAP7_75t_R _18164_ (.A(_09878_),
    .B(_02694_),
    .Y(_02714_));
 INVx1_ASAP7_75t_R _18165_ (.A(_00330_),
    .Y(_02715_));
 AO32x1_ASAP7_75t_R _18166_ (.A1(_02692_),
    .A2(_02713_),
    .A3(_02714_),
    .B1(_02690_),
    .B2(_02715_),
    .Y(_01909_));
 BUFx6f_ASAP7_75t_R _18167_ (.A(_08950_),
    .Y(_02716_));
 AND2x2_ASAP7_75t_R _18168_ (.A(_09881_),
    .B(_02694_),
    .Y(_02717_));
 INVx1_ASAP7_75t_R _18169_ (.A(_00297_),
    .Y(_02718_));
 AO32x1_ASAP7_75t_R _18170_ (.A1(_02692_),
    .A2(_02716_),
    .A3(_02717_),
    .B1(_02690_),
    .B2(_02718_),
    .Y(_01910_));
 BUFx6f_ASAP7_75t_R _18171_ (.A(_08969_),
    .Y(_02719_));
 AND2x2_ASAP7_75t_R _18172_ (.A(_09884_),
    .B(_02683_),
    .Y(_02720_));
 INVx1_ASAP7_75t_R _18173_ (.A(_00264_),
    .Y(_02721_));
 AO32x1_ASAP7_75t_R _18174_ (.A1(_02692_),
    .A2(_02719_),
    .A3(_02720_),
    .B1(_02674_),
    .B2(_02721_),
    .Y(_01911_));
 BUFx6f_ASAP7_75t_R _18175_ (.A(_08986_),
    .Y(_02722_));
 BUFx10_ASAP7_75t_R _18176_ (.A(_08996_),
    .Y(_02723_));
 NOR2x1_ASAP7_75t_R _18177_ (.A(_02723_),
    .B(_02674_),
    .Y(_02724_));
 INVx1_ASAP7_75t_R _18178_ (.A(_00231_),
    .Y(_02725_));
 AO32x1_ASAP7_75t_R _18179_ (.A1(_02692_),
    .A2(_02722_),
    .A3(_02724_),
    .B1(_02674_),
    .B2(_02725_),
    .Y(_01912_));
 INVx1_ASAP7_75t_R _18180_ (.A(_00197_),
    .Y(_02726_));
 AND2x2_ASAP7_75t_R _18181_ (.A(_09890_),
    .B(_02684_),
    .Y(_02727_));
 BUFx6f_ASAP7_75t_R _18182_ (.A(_09005_),
    .Y(_02728_));
 AO22x1_ASAP7_75t_R _18183_ (.A1(_02726_),
    .A2(_02678_),
    .B1(_02727_),
    .B2(_02728_),
    .Y(_01913_));
 BUFx6f_ASAP7_75t_R _18184_ (.A(_02546_),
    .Y(_02729_));
 BUFx4f_ASAP7_75t_R _18185_ (.A(_09024_),
    .Y(_02730_));
 AND4x1_ASAP7_75t_R _18186_ (.A(_09892_),
    .B(_09893_),
    .C(_09894_),
    .D(_02683_),
    .Y(_02731_));
 INVx1_ASAP7_75t_R _18187_ (.A(_00164_),
    .Y(_02732_));
 AO32x1_ASAP7_75t_R _18188_ (.A1(_02729_),
    .A2(_02730_),
    .A3(_02731_),
    .B1(_02674_),
    .B2(_02732_),
    .Y(_01914_));
 BUFx6f_ASAP7_75t_R _18189_ (.A(_09042_),
    .Y(_02733_));
 AND3x1_ASAP7_75t_R _18190_ (.A(_09897_),
    .B(_09898_),
    .C(_02694_),
    .Y(_02734_));
 INVx1_ASAP7_75t_R _18191_ (.A(_00130_),
    .Y(_02735_));
 AO32x1_ASAP7_75t_R _18192_ (.A1(_02729_),
    .A2(_02733_),
    .A3(_02734_),
    .B1(_02674_),
    .B2(_02735_),
    .Y(_01915_));
 NAND2x1_ASAP7_75t_R _18193_ (.A(_01027_),
    .B(_02678_),
    .Y(_02736_));
 OA21x2_ASAP7_75t_R _18194_ (.A1(_09901_),
    .A2(_02675_),
    .B(_02736_),
    .Y(_01916_));
 BUFx6f_ASAP7_75t_R _18195_ (.A(_09069_),
    .Y(_02737_));
 AND4x1_ASAP7_75t_R _18196_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .D(_02683_),
    .Y(_02738_));
 INVx1_ASAP7_75t_R _18197_ (.A(_00096_),
    .Y(_02739_));
 AO32x1_ASAP7_75t_R _18198_ (.A1(_02729_),
    .A2(_02737_),
    .A3(_02738_),
    .B1(_02674_),
    .B2(_02739_),
    .Y(_01917_));
 BUFx4f_ASAP7_75t_R _18199_ (.A(_09085_),
    .Y(_02740_));
 AND3x1_ASAP7_75t_R _18200_ (.A(_09908_),
    .B(_09909_),
    .C(_02694_),
    .Y(_02741_));
 INVx1_ASAP7_75t_R _18201_ (.A(_00064_),
    .Y(_02742_));
 AO32x1_ASAP7_75t_R _18202_ (.A1(_02729_),
    .A2(_02740_),
    .A3(_02741_),
    .B1(_02674_),
    .B2(_02742_),
    .Y(_01918_));
 NAND2x1_ASAP7_75t_R _18203_ (.A(_00994_),
    .B(_02678_),
    .Y(_02743_));
 OA21x2_ASAP7_75t_R _18204_ (.A1(_09912_),
    .A2(_02675_),
    .B(_02743_),
    .Y(_01919_));
 NAND2x1_ASAP7_75t_R _18205_ (.A(_00961_),
    .B(_02678_),
    .Y(_02744_));
 OA21x2_ASAP7_75t_R _18206_ (.A1(_09914_),
    .A2(_02675_),
    .B(_02744_),
    .Y(_01920_));
 BUFx10_ASAP7_75t_R _18207_ (.A(_09136_),
    .Y(_02745_));
 AND2x2_ASAP7_75t_R _18208_ (.A(_00927_),
    .B(_02674_),
    .Y(_02746_));
 AOI21x1_ASAP7_75t_R _18209_ (.A1(_02745_),
    .A2(_02684_),
    .B(_02746_),
    .Y(_01921_));
 NOR2x1_ASAP7_75t_R _18210_ (.A(_00894_),
    .B(_02684_),
    .Y(_02747_));
 AO21x1_ASAP7_75t_R _18211_ (.A1(_09917_),
    .A2(_02684_),
    .B(_02747_),
    .Y(_01922_));
 NOR2x1_ASAP7_75t_R _18212_ (.A(_00860_),
    .B(_02684_),
    .Y(_02748_));
 AO21x1_ASAP7_75t_R _18213_ (.A1(_09919_),
    .A2(_02684_),
    .B(_02748_),
    .Y(_01923_));
 NOR2x1_ASAP7_75t_R _18214_ (.A(_00827_),
    .B(_02684_),
    .Y(_02749_));
 AO21x1_ASAP7_75t_R _18215_ (.A1(_09921_),
    .A2(_02684_),
    .B(_02749_),
    .Y(_01924_));
 NAND2x1_ASAP7_75t_R _18216_ (.A(_00793_),
    .B(_02690_),
    .Y(_02750_));
 OA21x2_ASAP7_75t_R _18217_ (.A1(_09923_),
    .A2(_02678_),
    .B(_02750_),
    .Y(_01925_));
 OR3x4_ASAP7_75t_R _18218_ (.A(_09408_),
    .B(_08601_),
    .C(_09526_),
    .Y(_02751_));
 BUFx4f_ASAP7_75t_R _18219_ (.A(_02751_),
    .Y(_02752_));
 BUFx6f_ASAP7_75t_R _18220_ (.A(_02751_),
    .Y(_02753_));
 NAND2x1_ASAP7_75t_R _18221_ (.A(_00002_),
    .B(_02753_),
    .Y(_02754_));
 OA21x2_ASAP7_75t_R _18222_ (.A1(_02672_),
    .A2(_02752_),
    .B(_02754_),
    .Y(_01926_));
 BUFx6f_ASAP7_75t_R _18223_ (.A(_08654_),
    .Y(_02755_));
 NAND2x1_ASAP7_75t_R _18224_ (.A(_00734_),
    .B(_02753_),
    .Y(_02756_));
 OA21x2_ASAP7_75t_R _18225_ (.A1(_02755_),
    .A2(_02752_),
    .B(_02756_),
    .Y(_01927_));
 BUFx6f_ASAP7_75t_R _18226_ (.A(_08681_),
    .Y(_02757_));
 NAND2x1_ASAP7_75t_R _18227_ (.A(_00701_),
    .B(_02753_),
    .Y(_02758_));
 OA21x2_ASAP7_75t_R _18228_ (.A1(_02757_),
    .A2(_02752_),
    .B(_02758_),
    .Y(_01928_));
 BUFx6f_ASAP7_75t_R _18229_ (.A(_08697_),
    .Y(_02759_));
 NAND2x1_ASAP7_75t_R _18230_ (.A(_00668_),
    .B(_02753_),
    .Y(_02760_));
 OA21x2_ASAP7_75t_R _18231_ (.A1(_02759_),
    .A2(_02752_),
    .B(_02760_),
    .Y(_01929_));
 AND2x4_ASAP7_75t_R _18232_ (.A(_08602_),
    .B(_09288_),
    .Y(_02761_));
 BUFx6f_ASAP7_75t_R _18233_ (.A(_02761_),
    .Y(_02762_));
 BUFx4f_ASAP7_75t_R _18234_ (.A(_02751_),
    .Y(_02763_));
 AND2x2_ASAP7_75t_R _18235_ (.A(_00635_),
    .B(_02763_),
    .Y(_02764_));
 AOI21x1_ASAP7_75t_R _18236_ (.A1(_02682_),
    .A2(_02762_),
    .B(_02764_),
    .Y(_01930_));
 BUFx6f_ASAP7_75t_R _18237_ (.A(_08744_),
    .Y(_02765_));
 NAND2x1_ASAP7_75t_R _18238_ (.A(_00602_),
    .B(_02753_),
    .Y(_02766_));
 OA21x2_ASAP7_75t_R _18239_ (.A1(_02765_),
    .A2(_02752_),
    .B(_02766_),
    .Y(_01931_));
 AND2x2_ASAP7_75t_R _18240_ (.A(_00568_),
    .B(_02763_),
    .Y(_02767_));
 AOI21x1_ASAP7_75t_R _18241_ (.A1(_09769_),
    .A2(_02762_),
    .B(_02767_),
    .Y(_01932_));
 BUFx3_ASAP7_75t_R _18242_ (.A(_08786_),
    .Y(_02768_));
 BUFx3_ASAP7_75t_R _18243_ (.A(_08794_),
    .Y(_02769_));
 BUFx4f_ASAP7_75t_R _18244_ (.A(_02761_),
    .Y(_02770_));
 AND3x1_ASAP7_75t_R _18245_ (.A(_02768_),
    .B(_02769_),
    .C(_02770_),
    .Y(_02771_));
 BUFx6f_ASAP7_75t_R _18246_ (.A(_02751_),
    .Y(_02772_));
 AO32x1_ASAP7_75t_R _18247_ (.A1(_02688_),
    .A2(_02460_),
    .A3(_02771_),
    .B1(_02772_),
    .B2(_05708_),
    .Y(_01933_));
 BUFx4f_ASAP7_75t_R _18248_ (.A(_08821_),
    .Y(_02773_));
 AND2x2_ASAP7_75t_R _18249_ (.A(_02773_),
    .B(_02770_),
    .Y(_02774_));
 INVx1_ASAP7_75t_R _18250_ (.A(_00502_),
    .Y(_02775_));
 AO32x1_ASAP7_75t_R _18251_ (.A1(_02729_),
    .A2(_02693_),
    .A3(_02774_),
    .B1(_02772_),
    .B2(_02775_),
    .Y(_01934_));
 BUFx4f_ASAP7_75t_R _18252_ (.A(_08834_),
    .Y(_02776_));
 BUFx4f_ASAP7_75t_R _18253_ (.A(_08841_),
    .Y(_02777_));
 AND3x1_ASAP7_75t_R _18254_ (.A(_02776_),
    .B(_02777_),
    .C(_02770_),
    .Y(_02778_));
 INVx1_ASAP7_75t_R _18255_ (.A(_00469_),
    .Y(_02779_));
 AO32x1_ASAP7_75t_R _18256_ (.A1(_02729_),
    .A2(_02697_),
    .A3(_02778_),
    .B1(_02772_),
    .B2(_02779_),
    .Y(_01935_));
 BUFx4f_ASAP7_75t_R _18257_ (.A(_08851_),
    .Y(_02780_));
 BUFx4f_ASAP7_75t_R _18258_ (.A(_08860_),
    .Y(_02781_));
 AND3x1_ASAP7_75t_R _18259_ (.A(_02780_),
    .B(_02781_),
    .C(_02770_),
    .Y(_02782_));
 INVx1_ASAP7_75t_R _18260_ (.A(_00436_),
    .Y(_02783_));
 AO32x1_ASAP7_75t_R _18261_ (.A1(_02729_),
    .A2(_02700_),
    .A3(_02782_),
    .B1(_02772_),
    .B2(_02783_),
    .Y(_01936_));
 BUFx4f_ASAP7_75t_R _18262_ (.A(_08870_),
    .Y(_02784_));
 NAND2x1_ASAP7_75t_R _18263_ (.A(_01033_),
    .B(_02753_),
    .Y(_02785_));
 OA21x2_ASAP7_75t_R _18264_ (.A1(_02784_),
    .A2(_02752_),
    .B(_02785_),
    .Y(_01937_));
 BUFx4f_ASAP7_75t_R _18265_ (.A(_08892_),
    .Y(_02786_));
 AND2x2_ASAP7_75t_R _18266_ (.A(_02786_),
    .B(_02770_),
    .Y(_02787_));
 INVx1_ASAP7_75t_R _18267_ (.A(_00403_),
    .Y(_02788_));
 AO32x1_ASAP7_75t_R _18268_ (.A1(_02729_),
    .A2(_02704_),
    .A3(_02787_),
    .B1(_02772_),
    .B2(_02788_),
    .Y(_01938_));
 BUFx4f_ASAP7_75t_R _18269_ (.A(_08902_),
    .Y(_02789_));
 BUFx4f_ASAP7_75t_R _18270_ (.A(_08910_),
    .Y(_02790_));
 AND3x1_ASAP7_75t_R _18271_ (.A(_02789_),
    .B(_02790_),
    .C(_02770_),
    .Y(_02791_));
 INVx1_ASAP7_75t_R _18272_ (.A(_00370_),
    .Y(_02792_));
 AO32x1_ASAP7_75t_R _18273_ (.A1(_02729_),
    .A2(_02707_),
    .A3(_02791_),
    .B1(_02772_),
    .B2(_02792_),
    .Y(_01939_));
 BUFx4f_ASAP7_75t_R _18274_ (.A(_08929_),
    .Y(_02793_));
 AND2x2_ASAP7_75t_R _18275_ (.A(_02793_),
    .B(_02770_),
    .Y(_02794_));
 AO32x1_ASAP7_75t_R _18276_ (.A1(_02729_),
    .A2(_02710_),
    .A3(_02794_),
    .B1(_02772_),
    .B2(_05148_),
    .Y(_01940_));
 BUFx4f_ASAP7_75t_R _18277_ (.A(_02546_),
    .Y(_02795_));
 BUFx4f_ASAP7_75t_R _18278_ (.A(_08943_),
    .Y(_02796_));
 AND2x2_ASAP7_75t_R _18279_ (.A(_02796_),
    .B(_02770_),
    .Y(_02797_));
 INVx1_ASAP7_75t_R _18280_ (.A(_00303_),
    .Y(_02798_));
 AO32x1_ASAP7_75t_R _18281_ (.A1(_02795_),
    .A2(_02713_),
    .A3(_02797_),
    .B1(_02772_),
    .B2(_02798_),
    .Y(_01941_));
 BUFx4f_ASAP7_75t_R _18282_ (.A(_08962_),
    .Y(_02799_));
 AND2x2_ASAP7_75t_R _18283_ (.A(_02799_),
    .B(_02761_),
    .Y(_02800_));
 INVx1_ASAP7_75t_R _18284_ (.A(_00270_),
    .Y(_02801_));
 AO32x1_ASAP7_75t_R _18285_ (.A1(_02795_),
    .A2(_02716_),
    .A3(_02800_),
    .B1(_02772_),
    .B2(_02801_),
    .Y(_01942_));
 BUFx4f_ASAP7_75t_R _18286_ (.A(_08979_),
    .Y(_02802_));
 AND2x2_ASAP7_75t_R _18287_ (.A(_02802_),
    .B(_02761_),
    .Y(_02803_));
 INVx1_ASAP7_75t_R _18288_ (.A(_00237_),
    .Y(_02804_));
 AO32x1_ASAP7_75t_R _18289_ (.A1(_02795_),
    .A2(_02719_),
    .A3(_02803_),
    .B1(_02763_),
    .B2(_02804_),
    .Y(_01943_));
 NOR2x1_ASAP7_75t_R _18290_ (.A(_02723_),
    .B(_02763_),
    .Y(_02805_));
 AO32x1_ASAP7_75t_R _18291_ (.A1(_02795_),
    .A2(_02722_),
    .A3(_02805_),
    .B1(_02763_),
    .B2(_04731_),
    .Y(_01944_));
 INVx1_ASAP7_75t_R _18292_ (.A(_00170_),
    .Y(_02806_));
 BUFx6f_ASAP7_75t_R _18293_ (.A(_09017_),
    .Y(_02807_));
 AND2x2_ASAP7_75t_R _18294_ (.A(_02807_),
    .B(_02762_),
    .Y(_02808_));
 AO22x1_ASAP7_75t_R _18295_ (.A1(_02806_),
    .A2(_02753_),
    .B1(_02808_),
    .B2(_02728_),
    .Y(_01945_));
 BUFx4f_ASAP7_75t_R _18296_ (.A(_09030_),
    .Y(_02809_));
 BUFx4f_ASAP7_75t_R _18297_ (.A(_09031_),
    .Y(_02810_));
 BUFx4f_ASAP7_75t_R _18298_ (.A(_09035_),
    .Y(_02811_));
 AND4x1_ASAP7_75t_R _18299_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_02761_),
    .Y(_02812_));
 AO32x1_ASAP7_75t_R _18300_ (.A1(_02795_),
    .A2(_02730_),
    .A3(_02812_),
    .B1(_02763_),
    .B2(_04441_),
    .Y(_01946_));
 BUFx4f_ASAP7_75t_R _18301_ (.A(_09048_),
    .Y(_02813_));
 BUFx4f_ASAP7_75t_R _18302_ (.A(_09051_),
    .Y(_02814_));
 AND3x1_ASAP7_75t_R _18303_ (.A(_02813_),
    .B(_02814_),
    .C(_02770_),
    .Y(_02815_));
 AO32x1_ASAP7_75t_R _18304_ (.A1(_02795_),
    .A2(_02733_),
    .A3(_02815_),
    .B1(_02763_),
    .B2(_04367_),
    .Y(_01947_));
 BUFx6f_ASAP7_75t_R _18305_ (.A(_09063_),
    .Y(_02816_));
 NAND2x1_ASAP7_75t_R _18306_ (.A(_01000_),
    .B(_02753_),
    .Y(_02817_));
 OA21x2_ASAP7_75t_R _18307_ (.A1(_02816_),
    .A2(_02752_),
    .B(_02817_),
    .Y(_01948_));
 BUFx4f_ASAP7_75t_R _18308_ (.A(_09074_),
    .Y(_02818_));
 BUFx4f_ASAP7_75t_R _18309_ (.A(_09077_),
    .Y(_02819_));
 BUFx4f_ASAP7_75t_R _18310_ (.A(_09078_),
    .Y(_02820_));
 AND4x1_ASAP7_75t_R _18311_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_02761_),
    .Y(_02821_));
 AO32x1_ASAP7_75t_R _18312_ (.A1(_02795_),
    .A2(_02737_),
    .A3(_02821_),
    .B1(_02763_),
    .B2(_04184_),
    .Y(_01949_));
 BUFx4f_ASAP7_75t_R _18313_ (.A(_09094_),
    .Y(_02822_));
 BUFx3_ASAP7_75t_R _18314_ (.A(_09097_),
    .Y(_02823_));
 AND3x1_ASAP7_75t_R _18315_ (.A(_02822_),
    .B(_02823_),
    .C(_02770_),
    .Y(_02824_));
 INVx1_ASAP7_75t_R _18316_ (.A(_00037_),
    .Y(_02825_));
 AO32x1_ASAP7_75t_R _18317_ (.A1(_02795_),
    .A2(_02740_),
    .A3(_02824_),
    .B1(_02763_),
    .B2(_02825_),
    .Y(_01950_));
 BUFx6f_ASAP7_75t_R _18318_ (.A(_09109_),
    .Y(_02826_));
 NAND2x1_ASAP7_75t_R _18319_ (.A(_00967_),
    .B(_02753_),
    .Y(_02827_));
 OA21x2_ASAP7_75t_R _18320_ (.A1(_02826_),
    .A2(_02752_),
    .B(_02827_),
    .Y(_01951_));
 BUFx6f_ASAP7_75t_R _18321_ (.A(_09122_),
    .Y(_02828_));
 NAND2x1_ASAP7_75t_R _18322_ (.A(_00934_),
    .B(_02753_),
    .Y(_02829_));
 OA21x2_ASAP7_75t_R _18323_ (.A1(_02828_),
    .A2(_02752_),
    .B(_02829_),
    .Y(_01952_));
 AND2x2_ASAP7_75t_R _18324_ (.A(_00900_),
    .B(_02763_),
    .Y(_02830_));
 AOI21x1_ASAP7_75t_R _18325_ (.A1(_02745_),
    .A2(_02762_),
    .B(_02830_),
    .Y(_01953_));
 BUFx6f_ASAP7_75t_R _18326_ (.A(_09148_),
    .Y(_02831_));
 NOR2x1_ASAP7_75t_R _18327_ (.A(_00867_),
    .B(_02762_),
    .Y(_02832_));
 AO21x1_ASAP7_75t_R _18328_ (.A1(_02831_),
    .A2(_02762_),
    .B(_02832_),
    .Y(_01954_));
 BUFx6f_ASAP7_75t_R _18329_ (.A(_09158_),
    .Y(_02833_));
 NOR2x1_ASAP7_75t_R _18330_ (.A(_00833_),
    .B(_02762_),
    .Y(_02834_));
 AO21x1_ASAP7_75t_R _18331_ (.A1(_02833_),
    .A2(_02762_),
    .B(_02834_),
    .Y(_01955_));
 BUFx10_ASAP7_75t_R _18332_ (.A(_09173_),
    .Y(_02835_));
 NOR2x1_ASAP7_75t_R _18333_ (.A(_00800_),
    .B(_02762_),
    .Y(_02836_));
 AO21x1_ASAP7_75t_R _18334_ (.A1(_02835_),
    .A2(_02762_),
    .B(_02836_),
    .Y(_01956_));
 BUFx6f_ASAP7_75t_R _18335_ (.A(_09186_),
    .Y(_02837_));
 NAND2x1_ASAP7_75t_R _18336_ (.A(_00766_),
    .B(_02772_),
    .Y(_02838_));
 OA21x2_ASAP7_75t_R _18337_ (.A1(_02837_),
    .A2(_02752_),
    .B(_02838_),
    .Y(_01957_));
 NAND2x2_ASAP7_75t_R _18338_ (.A(_08871_),
    .B(_02614_),
    .Y(_02839_));
 BUFx4f_ASAP7_75t_R _18339_ (.A(_02839_),
    .Y(_02840_));
 BUFx6f_ASAP7_75t_R _18340_ (.A(_02839_),
    .Y(_02841_));
 NAND2x1_ASAP7_75t_R _18341_ (.A(_00030_),
    .B(_02841_),
    .Y(_02842_));
 OA21x2_ASAP7_75t_R _18342_ (.A1(_02672_),
    .A2(_02840_),
    .B(_02842_),
    .Y(_01958_));
 NAND2x1_ASAP7_75t_R _18343_ (.A(_00762_),
    .B(_02841_),
    .Y(_02843_));
 OA21x2_ASAP7_75t_R _18344_ (.A1(_02755_),
    .A2(_02840_),
    .B(_02843_),
    .Y(_01959_));
 NAND2x1_ASAP7_75t_R _18345_ (.A(_00729_),
    .B(_02841_),
    .Y(_02844_));
 OA21x2_ASAP7_75t_R _18346_ (.A1(_02757_),
    .A2(_02840_),
    .B(_02844_),
    .Y(_01960_));
 NAND2x1_ASAP7_75t_R _18347_ (.A(_00696_),
    .B(_02841_),
    .Y(_02845_));
 OA21x2_ASAP7_75t_R _18348_ (.A1(_02759_),
    .A2(_02840_),
    .B(_02845_),
    .Y(_01961_));
 AND2x4_ASAP7_75t_R _18349_ (.A(_08602_),
    .B(_02613_),
    .Y(_02846_));
 BUFx16f_ASAP7_75t_R _18350_ (.A(_02846_),
    .Y(_02847_));
 BUFx12_ASAP7_75t_R _18351_ (.A(_02839_),
    .Y(_02848_));
 AND2x2_ASAP7_75t_R _18352_ (.A(_00663_),
    .B(_02848_),
    .Y(_02849_));
 AOI21x1_ASAP7_75t_R _18353_ (.A1(_02682_),
    .A2(_02847_),
    .B(_02849_),
    .Y(_01962_));
 NAND2x1_ASAP7_75t_R _18354_ (.A(_00630_),
    .B(_02841_),
    .Y(_02850_));
 OA21x2_ASAP7_75t_R _18355_ (.A1(_02765_),
    .A2(_02840_),
    .B(_02850_),
    .Y(_01963_));
 AO21x1_ASAP7_75t_R _18356_ (.A1(_08871_),
    .A2(_02614_),
    .B(_00596_),
    .Y(_02851_));
 OAI21x1_ASAP7_75t_R _18357_ (.A1(_09937_),
    .A2(_02840_),
    .B(_02851_),
    .Y(_01964_));
 AND3x1_ASAP7_75t_R _18358_ (.A(_02768_),
    .B(_02769_),
    .C(_02847_),
    .Y(_02852_));
 BUFx12_ASAP7_75t_R _18359_ (.A(_02839_),
    .Y(_02853_));
 AO32x1_ASAP7_75t_R _18360_ (.A1(_02688_),
    .A2(_02460_),
    .A3(_02852_),
    .B1(_02853_),
    .B2(_05727_),
    .Y(_01965_));
 BUFx4f_ASAP7_75t_R _18361_ (.A(_02846_),
    .Y(_02854_));
 AND2x2_ASAP7_75t_R _18362_ (.A(_02773_),
    .B(_02854_),
    .Y(_02855_));
 INVx1_ASAP7_75t_R _18363_ (.A(_00530_),
    .Y(_02856_));
 AO32x1_ASAP7_75t_R _18364_ (.A1(_02795_),
    .A2(_02693_),
    .A3(_02855_),
    .B1(_02853_),
    .B2(_02856_),
    .Y(_01966_));
 AND3x1_ASAP7_75t_R _18365_ (.A(_02776_),
    .B(_02777_),
    .C(_02854_),
    .Y(_02857_));
 INVx1_ASAP7_75t_R _18366_ (.A(_00497_),
    .Y(_02858_));
 AO32x1_ASAP7_75t_R _18367_ (.A1(_02795_),
    .A2(_02697_),
    .A3(_02857_),
    .B1(_02853_),
    .B2(_02858_),
    .Y(_01967_));
 BUFx4f_ASAP7_75t_R _18368_ (.A(_02546_),
    .Y(_02859_));
 AND3x1_ASAP7_75t_R _18369_ (.A(_02780_),
    .B(_02781_),
    .C(_02854_),
    .Y(_02860_));
 INVx1_ASAP7_75t_R _18370_ (.A(_00464_),
    .Y(_02861_));
 AO32x1_ASAP7_75t_R _18371_ (.A1(_02859_),
    .A2(_02700_),
    .A3(_02860_),
    .B1(_02853_),
    .B2(_02861_),
    .Y(_01968_));
 NAND2x1_ASAP7_75t_R _18372_ (.A(_01061_),
    .B(_02841_),
    .Y(_02862_));
 OA21x2_ASAP7_75t_R _18373_ (.A1(_02784_),
    .A2(_02840_),
    .B(_02862_),
    .Y(_01969_));
 AND2x2_ASAP7_75t_R _18374_ (.A(_02786_),
    .B(_02854_),
    .Y(_02863_));
 INVx1_ASAP7_75t_R _18375_ (.A(_00431_),
    .Y(_02864_));
 AO32x1_ASAP7_75t_R _18376_ (.A1(_02859_),
    .A2(_02704_),
    .A3(_02863_),
    .B1(_02853_),
    .B2(_02864_),
    .Y(_01970_));
 AND3x1_ASAP7_75t_R _18377_ (.A(_02789_),
    .B(_02790_),
    .C(_02854_),
    .Y(_02865_));
 INVx1_ASAP7_75t_R _18378_ (.A(_00398_),
    .Y(_02866_));
 AO32x1_ASAP7_75t_R _18379_ (.A1(_02859_),
    .A2(_02707_),
    .A3(_02865_),
    .B1(_02853_),
    .B2(_02866_),
    .Y(_01971_));
 AND2x2_ASAP7_75t_R _18380_ (.A(_02793_),
    .B(_02854_),
    .Y(_02867_));
 INVx1_ASAP7_75t_R _18381_ (.A(_00365_),
    .Y(_02868_));
 AO32x1_ASAP7_75t_R _18382_ (.A1(_02859_),
    .A2(_02710_),
    .A3(_02867_),
    .B1(_02853_),
    .B2(_02868_),
    .Y(_01972_));
 AND2x2_ASAP7_75t_R _18383_ (.A(_02796_),
    .B(_02854_),
    .Y(_02869_));
 INVx1_ASAP7_75t_R _18384_ (.A(_00331_),
    .Y(_02870_));
 AO32x1_ASAP7_75t_R _18385_ (.A1(_02859_),
    .A2(_02713_),
    .A3(_02869_),
    .B1(_02853_),
    .B2(_02870_),
    .Y(_01973_));
 AND2x2_ASAP7_75t_R _18386_ (.A(_02799_),
    .B(_02854_),
    .Y(_02871_));
 AO32x1_ASAP7_75t_R _18387_ (.A1(_02859_),
    .A2(_02716_),
    .A3(_02871_),
    .B1(_02848_),
    .B2(_04900_),
    .Y(_01974_));
 AND2x2_ASAP7_75t_R _18388_ (.A(_02802_),
    .B(_02846_),
    .Y(_02872_));
 INVx1_ASAP7_75t_R _18389_ (.A(_00265_),
    .Y(_02873_));
 AO32x1_ASAP7_75t_R _18390_ (.A1(_02859_),
    .A2(_02719_),
    .A3(_02872_),
    .B1(_02848_),
    .B2(_02873_),
    .Y(_01975_));
 NOR2x1_ASAP7_75t_R _18391_ (.A(_02723_),
    .B(_02848_),
    .Y(_02874_));
 INVx1_ASAP7_75t_R _18392_ (.A(_00232_),
    .Y(_02875_));
 AO32x1_ASAP7_75t_R _18393_ (.A1(_02859_),
    .A2(_02722_),
    .A3(_02874_),
    .B1(_02848_),
    .B2(_02875_),
    .Y(_01976_));
 INVx1_ASAP7_75t_R _18394_ (.A(_00198_),
    .Y(_02876_));
 AND2x2_ASAP7_75t_R _18395_ (.A(_02807_),
    .B(_02847_),
    .Y(_02877_));
 AO22x1_ASAP7_75t_R _18396_ (.A1(_02876_),
    .A2(_02841_),
    .B1(_02877_),
    .B2(_02728_),
    .Y(_01977_));
 AND4x1_ASAP7_75t_R _18397_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_02846_),
    .Y(_02878_));
 INVx1_ASAP7_75t_R _18398_ (.A(_00165_),
    .Y(_02879_));
 AO32x1_ASAP7_75t_R _18399_ (.A1(_02859_),
    .A2(_02730_),
    .A3(_02878_),
    .B1(_02848_),
    .B2(_02879_),
    .Y(_01978_));
 AND3x1_ASAP7_75t_R _18400_ (.A(_02813_),
    .B(_02814_),
    .C(_02854_),
    .Y(_02880_));
 INVx1_ASAP7_75t_R _18401_ (.A(_00131_),
    .Y(_02881_));
 AO32x1_ASAP7_75t_R _18402_ (.A1(_02859_),
    .A2(_02733_),
    .A3(_02880_),
    .B1(_02848_),
    .B2(_02881_),
    .Y(_01979_));
 NAND2x1_ASAP7_75t_R _18403_ (.A(_01028_),
    .B(_02841_),
    .Y(_02882_));
 OA21x2_ASAP7_75t_R _18404_ (.A1(_02816_),
    .A2(_02840_),
    .B(_02882_),
    .Y(_01980_));
 BUFx4f_ASAP7_75t_R _18405_ (.A(_02546_),
    .Y(_02883_));
 AND4x1_ASAP7_75t_R _18406_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_02846_),
    .Y(_02884_));
 INVx1_ASAP7_75t_R _18407_ (.A(_00097_),
    .Y(_02885_));
 AO32x1_ASAP7_75t_R _18408_ (.A1(_02883_),
    .A2(_02737_),
    .A3(_02884_),
    .B1(_02848_),
    .B2(_02885_),
    .Y(_01981_));
 AND3x1_ASAP7_75t_R _18409_ (.A(_02822_),
    .B(_02823_),
    .C(_02854_),
    .Y(_02886_));
 AO32x1_ASAP7_75t_R _18410_ (.A1(_02883_),
    .A2(_02740_),
    .A3(_02886_),
    .B1(_02848_),
    .B2(_03846_),
    .Y(_01982_));
 NAND2x1_ASAP7_75t_R _18411_ (.A(_00995_),
    .B(_02841_),
    .Y(_02887_));
 OA21x2_ASAP7_75t_R _18412_ (.A1(_02826_),
    .A2(_02840_),
    .B(_02887_),
    .Y(_01983_));
 NAND2x1_ASAP7_75t_R _18413_ (.A(_00962_),
    .B(_02853_),
    .Y(_02888_));
 OA21x2_ASAP7_75t_R _18414_ (.A1(_02828_),
    .A2(_02840_),
    .B(_02888_),
    .Y(_01984_));
 AND2x2_ASAP7_75t_R _18415_ (.A(_00928_),
    .B(_02848_),
    .Y(_02889_));
 AOI21x1_ASAP7_75t_R _18416_ (.A1(_02745_),
    .A2(_02847_),
    .B(_02889_),
    .Y(_01985_));
 NOR2x1_ASAP7_75t_R _18417_ (.A(_00895_),
    .B(_02847_),
    .Y(_02890_));
 AO21x1_ASAP7_75t_R _18418_ (.A1(_02831_),
    .A2(_02847_),
    .B(_02890_),
    .Y(_01986_));
 NOR2x1_ASAP7_75t_R _18419_ (.A(_00861_),
    .B(_02847_),
    .Y(_02891_));
 AO21x1_ASAP7_75t_R _18420_ (.A1(_02833_),
    .A2(_02847_),
    .B(_02891_),
    .Y(_01987_));
 NOR2x1_ASAP7_75t_R _18421_ (.A(_00828_),
    .B(_02847_),
    .Y(_02892_));
 AO21x1_ASAP7_75t_R _18422_ (.A1(_02835_),
    .A2(_02847_),
    .B(_02892_),
    .Y(_01988_));
 NAND2x1_ASAP7_75t_R _18423_ (.A(_00794_),
    .B(_02853_),
    .Y(_02893_));
 OA21x2_ASAP7_75t_R _18424_ (.A1(_02837_),
    .A2(_02841_),
    .B(_02893_),
    .Y(_01989_));
 NAND2x2_ASAP7_75t_R _18425_ (.A(_09191_),
    .B(_02614_),
    .Y(_02894_));
 BUFx10_ASAP7_75t_R _18426_ (.A(_02894_),
    .Y(_02895_));
 BUFx4f_ASAP7_75t_R _18427_ (.A(_02895_),
    .Y(_02896_));
 BUFx6f_ASAP7_75t_R _18428_ (.A(_02894_),
    .Y(_02897_));
 NAND2x1_ASAP7_75t_R _18429_ (.A(_00031_),
    .B(_02897_),
    .Y(_02898_));
 OA21x2_ASAP7_75t_R _18430_ (.A1(_02672_),
    .A2(_02896_),
    .B(_02898_),
    .Y(_01990_));
 NAND2x1_ASAP7_75t_R _18431_ (.A(_00763_),
    .B(_02897_),
    .Y(_02899_));
 OA21x2_ASAP7_75t_R _18432_ (.A1(_02755_),
    .A2(_02896_),
    .B(_02899_),
    .Y(_01991_));
 NAND2x1_ASAP7_75t_R _18433_ (.A(_00730_),
    .B(_02897_),
    .Y(_02900_));
 OA21x2_ASAP7_75t_R _18434_ (.A1(_02757_),
    .A2(_02896_),
    .B(_02900_),
    .Y(_01992_));
 NAND2x1_ASAP7_75t_R _18435_ (.A(_00697_),
    .B(_02897_),
    .Y(_02901_));
 OA21x2_ASAP7_75t_R _18436_ (.A1(_02759_),
    .A2(_02896_),
    .B(_02901_),
    .Y(_01993_));
 AND2x4_ASAP7_75t_R _18437_ (.A(_09190_),
    .B(_02613_),
    .Y(_02902_));
 BUFx16f_ASAP7_75t_R _18438_ (.A(_02902_),
    .Y(_02903_));
 AND2x2_ASAP7_75t_R _18439_ (.A(_00664_),
    .B(_02895_),
    .Y(_02904_));
 AOI21x1_ASAP7_75t_R _18440_ (.A1(_02682_),
    .A2(_02903_),
    .B(_02904_),
    .Y(_01994_));
 NAND2x1_ASAP7_75t_R _18441_ (.A(_00631_),
    .B(_02897_),
    .Y(_02905_));
 OA21x2_ASAP7_75t_R _18442_ (.A1(_02765_),
    .A2(_02896_),
    .B(_02905_),
    .Y(_01995_));
 AO21x1_ASAP7_75t_R _18443_ (.A1(_09191_),
    .A2(_02614_),
    .B(_00597_),
    .Y(_02906_));
 OAI21x1_ASAP7_75t_R _18444_ (.A1(_09937_),
    .A2(_02896_),
    .B(_02906_),
    .Y(_01996_));
 AND3x1_ASAP7_75t_R _18445_ (.A(_02768_),
    .B(_02769_),
    .C(_02903_),
    .Y(_02907_));
 BUFx10_ASAP7_75t_R _18446_ (.A(_02894_),
    .Y(_02908_));
 AO32x1_ASAP7_75t_R _18447_ (.A1(_02688_),
    .A2(_02460_),
    .A3(_02907_),
    .B1(_02908_),
    .B2(_05729_),
    .Y(_01997_));
 BUFx4f_ASAP7_75t_R _18448_ (.A(_02902_),
    .Y(_02909_));
 AND2x2_ASAP7_75t_R _18449_ (.A(_02773_),
    .B(_02909_),
    .Y(_02910_));
 INVx1_ASAP7_75t_R _18450_ (.A(_00531_),
    .Y(_02911_));
 AO32x1_ASAP7_75t_R _18451_ (.A1(_02883_),
    .A2(_02693_),
    .A3(_02910_),
    .B1(_02908_),
    .B2(_02911_),
    .Y(_01998_));
 AND3x1_ASAP7_75t_R _18452_ (.A(_02776_),
    .B(_02777_),
    .C(_02909_),
    .Y(_02912_));
 INVx1_ASAP7_75t_R _18453_ (.A(_00498_),
    .Y(_02913_));
 AO32x1_ASAP7_75t_R _18454_ (.A1(_02883_),
    .A2(_02697_),
    .A3(_02912_),
    .B1(_02908_),
    .B2(_02913_),
    .Y(_01999_));
 AND3x1_ASAP7_75t_R _18455_ (.A(_02780_),
    .B(_02781_),
    .C(_02909_),
    .Y(_02914_));
 INVx1_ASAP7_75t_R _18456_ (.A(_00465_),
    .Y(_02915_));
 AO32x1_ASAP7_75t_R _18457_ (.A1(_02883_),
    .A2(_02700_),
    .A3(_02914_),
    .B1(_02908_),
    .B2(_02915_),
    .Y(_02000_));
 NAND2x1_ASAP7_75t_R _18458_ (.A(_01062_),
    .B(_02897_),
    .Y(_02916_));
 OA21x2_ASAP7_75t_R _18459_ (.A1(_02784_),
    .A2(_02896_),
    .B(_02916_),
    .Y(_02001_));
 AND2x2_ASAP7_75t_R _18460_ (.A(_02786_),
    .B(_02909_),
    .Y(_02917_));
 INVx1_ASAP7_75t_R _18461_ (.A(_00432_),
    .Y(_02918_));
 AO32x1_ASAP7_75t_R _18462_ (.A1(_02883_),
    .A2(_02704_),
    .A3(_02917_),
    .B1(_02908_),
    .B2(_02918_),
    .Y(_02002_));
 AND3x1_ASAP7_75t_R _18463_ (.A(_02789_),
    .B(_02790_),
    .C(_02909_),
    .Y(_02919_));
 INVx1_ASAP7_75t_R _18464_ (.A(_00399_),
    .Y(_02920_));
 AO32x1_ASAP7_75t_R _18465_ (.A1(_02883_),
    .A2(_02707_),
    .A3(_02919_),
    .B1(_02908_),
    .B2(_02920_),
    .Y(_02003_));
 AND2x2_ASAP7_75t_R _18466_ (.A(_02793_),
    .B(_02909_),
    .Y(_02921_));
 INVx1_ASAP7_75t_R _18467_ (.A(_00366_),
    .Y(_02922_));
 AO32x1_ASAP7_75t_R _18468_ (.A1(_02883_),
    .A2(_02710_),
    .A3(_02921_),
    .B1(_02908_),
    .B2(_02922_),
    .Y(_02004_));
 AND2x2_ASAP7_75t_R _18469_ (.A(_02796_),
    .B(_02909_),
    .Y(_02923_));
 INVx1_ASAP7_75t_R _18470_ (.A(_00332_),
    .Y(_02924_));
 AO32x1_ASAP7_75t_R _18471_ (.A1(_02883_),
    .A2(_02713_),
    .A3(_02923_),
    .B1(_02908_),
    .B2(_02924_),
    .Y(_02005_));
 AND2x2_ASAP7_75t_R _18472_ (.A(_02799_),
    .B(_02909_),
    .Y(_02925_));
 AO32x1_ASAP7_75t_R _18473_ (.A1(_02883_),
    .A2(_02716_),
    .A3(_02925_),
    .B1(_02908_),
    .B2(_04902_),
    .Y(_02006_));
 BUFx4f_ASAP7_75t_R _18474_ (.A(_02546_),
    .Y(_02926_));
 AND2x2_ASAP7_75t_R _18475_ (.A(_02802_),
    .B(_02902_),
    .Y(_02927_));
 INVx1_ASAP7_75t_R _18476_ (.A(_00266_),
    .Y(_02928_));
 AO32x1_ASAP7_75t_R _18477_ (.A1(_02926_),
    .A2(_02719_),
    .A3(_02927_),
    .B1(_02895_),
    .B2(_02928_),
    .Y(_02007_));
 NOR2x1_ASAP7_75t_R _18478_ (.A(_02723_),
    .B(_02895_),
    .Y(_02929_));
 INVx1_ASAP7_75t_R _18479_ (.A(_00233_),
    .Y(_02930_));
 AO32x1_ASAP7_75t_R _18480_ (.A1(_02926_),
    .A2(_02722_),
    .A3(_02929_),
    .B1(_02895_),
    .B2(_02930_),
    .Y(_02008_));
 INVx1_ASAP7_75t_R _18481_ (.A(_00199_),
    .Y(_02931_));
 AND2x2_ASAP7_75t_R _18482_ (.A(_02807_),
    .B(_02903_),
    .Y(_02932_));
 AO22x1_ASAP7_75t_R _18483_ (.A1(_02931_),
    .A2(_02897_),
    .B1(_02932_),
    .B2(_02728_),
    .Y(_02009_));
 AND4x1_ASAP7_75t_R _18484_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_02902_),
    .Y(_02933_));
 INVx1_ASAP7_75t_R _18485_ (.A(_00166_),
    .Y(_02934_));
 AO32x1_ASAP7_75t_R _18486_ (.A1(_02926_),
    .A2(_02730_),
    .A3(_02933_),
    .B1(_02895_),
    .B2(_02934_),
    .Y(_02010_));
 AND3x1_ASAP7_75t_R _18487_ (.A(_02813_),
    .B(_02814_),
    .C(_02909_),
    .Y(_02935_));
 INVx1_ASAP7_75t_R _18488_ (.A(_00132_),
    .Y(_02936_));
 AO32x1_ASAP7_75t_R _18489_ (.A1(_02926_),
    .A2(_02733_),
    .A3(_02935_),
    .B1(_02895_),
    .B2(_02936_),
    .Y(_02011_));
 NAND2x1_ASAP7_75t_R _18490_ (.A(_01029_),
    .B(_02897_),
    .Y(_02937_));
 OA21x2_ASAP7_75t_R _18491_ (.A1(_02816_),
    .A2(_02896_),
    .B(_02937_),
    .Y(_02012_));
 AND4x1_ASAP7_75t_R _18492_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_02902_),
    .Y(_02938_));
 INVx1_ASAP7_75t_R _18493_ (.A(_00098_),
    .Y(_02939_));
 AO32x1_ASAP7_75t_R _18494_ (.A1(_02926_),
    .A2(_02737_),
    .A3(_02938_),
    .B1(_02895_),
    .B2(_02939_),
    .Y(_02013_));
 AND3x1_ASAP7_75t_R _18495_ (.A(_02822_),
    .B(_02823_),
    .C(_02909_),
    .Y(_02940_));
 AO32x1_ASAP7_75t_R _18496_ (.A1(_02926_),
    .A2(_02740_),
    .A3(_02940_),
    .B1(_02895_),
    .B2(_03841_),
    .Y(_02014_));
 AO21x1_ASAP7_75t_R _18497_ (.A1(_09191_),
    .A2(_02614_),
    .B(_06915_),
    .Y(_02941_));
 OA21x2_ASAP7_75t_R _18498_ (.A1(_02826_),
    .A2(_02896_),
    .B(_02941_),
    .Y(_02015_));
 NAND2x1_ASAP7_75t_R _18499_ (.A(_00963_),
    .B(_02897_),
    .Y(_02942_));
 OA21x2_ASAP7_75t_R _18500_ (.A1(_02828_),
    .A2(_02896_),
    .B(_02942_),
    .Y(_02016_));
 AND2x2_ASAP7_75t_R _18501_ (.A(_00929_),
    .B(_02895_),
    .Y(_02943_));
 AOI21x1_ASAP7_75t_R _18502_ (.A1(_02745_),
    .A2(_02903_),
    .B(_02943_),
    .Y(_02017_));
 NOR2x1_ASAP7_75t_R _18503_ (.A(_00896_),
    .B(_02903_),
    .Y(_02944_));
 AO21x1_ASAP7_75t_R _18504_ (.A1(_02831_),
    .A2(_02903_),
    .B(_02944_),
    .Y(_02018_));
 NOR2x1_ASAP7_75t_R _18505_ (.A(_00862_),
    .B(_02903_),
    .Y(_02945_));
 AO21x1_ASAP7_75t_R _18506_ (.A1(_02833_),
    .A2(_02903_),
    .B(_02945_),
    .Y(_02019_));
 NOR2x1_ASAP7_75t_R _18507_ (.A(_00829_),
    .B(_02903_),
    .Y(_02946_));
 AO21x1_ASAP7_75t_R _18508_ (.A1(_02835_),
    .A2(_02903_),
    .B(_02946_),
    .Y(_02020_));
 NAND2x1_ASAP7_75t_R _18509_ (.A(_00795_),
    .B(_02908_),
    .Y(_02947_));
 OA21x2_ASAP7_75t_R _18510_ (.A1(_02837_),
    .A2(_02897_),
    .B(_02947_),
    .Y(_02021_));
 OR3x4_ASAP7_75t_R _18511_ (.A(_09408_),
    .B(_09349_),
    .C(_09526_),
    .Y(_02948_));
 BUFx4f_ASAP7_75t_R _18512_ (.A(_02948_),
    .Y(_02949_));
 BUFx6f_ASAP7_75t_R _18513_ (.A(_02948_),
    .Y(_02950_));
 NAND2x1_ASAP7_75t_R _18514_ (.A(_00003_),
    .B(_02950_),
    .Y(_02951_));
 OA21x2_ASAP7_75t_R _18515_ (.A1(_02672_),
    .A2(_02949_),
    .B(_02951_),
    .Y(_02022_));
 NAND2x1_ASAP7_75t_R _18516_ (.A(_00735_),
    .B(_02950_),
    .Y(_02952_));
 OA21x2_ASAP7_75t_R _18517_ (.A1(_02755_),
    .A2(_02949_),
    .B(_02952_),
    .Y(_02023_));
 NAND2x1_ASAP7_75t_R _18518_ (.A(_00702_),
    .B(_02950_),
    .Y(_02953_));
 OA21x2_ASAP7_75t_R _18519_ (.A1(_02757_),
    .A2(_02949_),
    .B(_02953_),
    .Y(_02024_));
 NAND2x1_ASAP7_75t_R _18520_ (.A(_00669_),
    .B(_02950_),
    .Y(_02954_));
 OA21x2_ASAP7_75t_R _18521_ (.A1(_02759_),
    .A2(_02949_),
    .B(_02954_),
    .Y(_02025_));
 AND2x4_ASAP7_75t_R _18522_ (.A(_09190_),
    .B(_09288_),
    .Y(_02955_));
 BUFx10_ASAP7_75t_R _18523_ (.A(_02955_),
    .Y(_02956_));
 BUFx4f_ASAP7_75t_R _18524_ (.A(_02948_),
    .Y(_02957_));
 AND2x2_ASAP7_75t_R _18525_ (.A(_00636_),
    .B(_02957_),
    .Y(_02958_));
 AOI21x1_ASAP7_75t_R _18526_ (.A1(_02682_),
    .A2(_02956_),
    .B(_02958_),
    .Y(_02026_));
 NAND2x1_ASAP7_75t_R _18527_ (.A(_00603_),
    .B(_02950_),
    .Y(_02959_));
 OA21x2_ASAP7_75t_R _18528_ (.A1(_02765_),
    .A2(_02949_),
    .B(_02959_),
    .Y(_02027_));
 AND2x2_ASAP7_75t_R _18529_ (.A(_00569_),
    .B(_02957_),
    .Y(_02960_));
 AOI21x1_ASAP7_75t_R _18530_ (.A1(_09769_),
    .A2(_02956_),
    .B(_02960_),
    .Y(_02028_));
 BUFx4f_ASAP7_75t_R _18531_ (.A(_02955_),
    .Y(_02961_));
 AND3x1_ASAP7_75t_R _18532_ (.A(_02768_),
    .B(_02769_),
    .C(_02961_),
    .Y(_02962_));
 BUFx6f_ASAP7_75t_R _18533_ (.A(_02948_),
    .Y(_02963_));
 INVx1_ASAP7_75t_R _18534_ (.A(_00536_),
    .Y(_02964_));
 AO32x1_ASAP7_75t_R _18535_ (.A1(_02688_),
    .A2(_02460_),
    .A3(_02962_),
    .B1(_02963_),
    .B2(_02964_),
    .Y(_02029_));
 AND2x2_ASAP7_75t_R _18536_ (.A(_02773_),
    .B(_02961_),
    .Y(_02965_));
 INVx1_ASAP7_75t_R _18537_ (.A(_00503_),
    .Y(_02966_));
 AO32x1_ASAP7_75t_R _18538_ (.A1(_02926_),
    .A2(_02693_),
    .A3(_02965_),
    .B1(_02963_),
    .B2(_02966_),
    .Y(_02030_));
 AND3x1_ASAP7_75t_R _18539_ (.A(_02776_),
    .B(_02777_),
    .C(_02961_),
    .Y(_02967_));
 INVx1_ASAP7_75t_R _18540_ (.A(_00470_),
    .Y(_02968_));
 AO32x1_ASAP7_75t_R _18541_ (.A1(_02926_),
    .A2(_02697_),
    .A3(_02967_),
    .B1(_02963_),
    .B2(_02968_),
    .Y(_02031_));
 AND3x1_ASAP7_75t_R _18542_ (.A(_02780_),
    .B(_02781_),
    .C(_02961_),
    .Y(_02969_));
 INVx1_ASAP7_75t_R _18543_ (.A(_00437_),
    .Y(_02970_));
 AO32x1_ASAP7_75t_R _18544_ (.A1(_02926_),
    .A2(_02700_),
    .A3(_02969_),
    .B1(_02963_),
    .B2(_02970_),
    .Y(_02032_));
 NAND2x1_ASAP7_75t_R _18545_ (.A(_01034_),
    .B(_02950_),
    .Y(_02971_));
 OA21x2_ASAP7_75t_R _18546_ (.A1(_02784_),
    .A2(_02949_),
    .B(_02971_),
    .Y(_02033_));
 AND2x2_ASAP7_75t_R _18547_ (.A(_02786_),
    .B(_02961_),
    .Y(_02972_));
 INVx1_ASAP7_75t_R _18548_ (.A(_00404_),
    .Y(_02973_));
 AO32x1_ASAP7_75t_R _18549_ (.A1(_02926_),
    .A2(_02704_),
    .A3(_02972_),
    .B1(_02963_),
    .B2(_02973_),
    .Y(_02034_));
 BUFx4f_ASAP7_75t_R _18550_ (.A(_02546_),
    .Y(_02974_));
 AND3x1_ASAP7_75t_R _18551_ (.A(_02789_),
    .B(_02790_),
    .C(_02961_),
    .Y(_02975_));
 INVx1_ASAP7_75t_R _18552_ (.A(_00371_),
    .Y(_02976_));
 AO32x1_ASAP7_75t_R _18553_ (.A1(_02974_),
    .A2(_02707_),
    .A3(_02975_),
    .B1(_02963_),
    .B2(_02976_),
    .Y(_02035_));
 AND2x2_ASAP7_75t_R _18554_ (.A(_02793_),
    .B(_02961_),
    .Y(_02977_));
 INVx1_ASAP7_75t_R _18555_ (.A(_00338_),
    .Y(_02978_));
 AO32x1_ASAP7_75t_R _18556_ (.A1(_02974_),
    .A2(_02710_),
    .A3(_02977_),
    .B1(_02963_),
    .B2(_02978_),
    .Y(_02036_));
 AND2x2_ASAP7_75t_R _18557_ (.A(_02796_),
    .B(_02961_),
    .Y(_02979_));
 INVx1_ASAP7_75t_R _18558_ (.A(_00304_),
    .Y(_02980_));
 AO32x1_ASAP7_75t_R _18559_ (.A1(_02974_),
    .A2(_02713_),
    .A3(_02979_),
    .B1(_02963_),
    .B2(_02980_),
    .Y(_02037_));
 AND2x2_ASAP7_75t_R _18560_ (.A(_02799_),
    .B(_02955_),
    .Y(_02981_));
 INVx1_ASAP7_75t_R _18561_ (.A(_00271_),
    .Y(_02982_));
 AO32x1_ASAP7_75t_R _18562_ (.A1(_02974_),
    .A2(_02716_),
    .A3(_02981_),
    .B1(_02963_),
    .B2(_02982_),
    .Y(_02038_));
 AND2x2_ASAP7_75t_R _18563_ (.A(_02802_),
    .B(_02955_),
    .Y(_02983_));
 INVx1_ASAP7_75t_R _18564_ (.A(_00238_),
    .Y(_02984_));
 AO32x1_ASAP7_75t_R _18565_ (.A1(_02974_),
    .A2(_02719_),
    .A3(_02983_),
    .B1(_02957_),
    .B2(_02984_),
    .Y(_02039_));
 NOR2x1_ASAP7_75t_R _18566_ (.A(_02723_),
    .B(_02957_),
    .Y(_02985_));
 INVx1_ASAP7_75t_R _18567_ (.A(_00205_),
    .Y(_02986_));
 AO32x1_ASAP7_75t_R _18568_ (.A1(_02974_),
    .A2(_02722_),
    .A3(_02985_),
    .B1(_02957_),
    .B2(_02986_),
    .Y(_02040_));
 INVx1_ASAP7_75t_R _18569_ (.A(_00171_),
    .Y(_02987_));
 AND2x2_ASAP7_75t_R _18570_ (.A(_02807_),
    .B(_02956_),
    .Y(_02988_));
 AO22x1_ASAP7_75t_R _18571_ (.A1(_02987_),
    .A2(_02950_),
    .B1(_02988_),
    .B2(_02728_),
    .Y(_02041_));
 AND4x1_ASAP7_75t_R _18572_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_02955_),
    .Y(_02989_));
 INVx1_ASAP7_75t_R _18573_ (.A(_00138_),
    .Y(_02990_));
 AO32x1_ASAP7_75t_R _18574_ (.A1(_02974_),
    .A2(_02730_),
    .A3(_02989_),
    .B1(_02957_),
    .B2(_02990_),
    .Y(_02042_));
 AND3x1_ASAP7_75t_R _18575_ (.A(_02813_),
    .B(_02814_),
    .C(_02961_),
    .Y(_02991_));
 INVx1_ASAP7_75t_R _18576_ (.A(_00104_),
    .Y(_02992_));
 AO32x1_ASAP7_75t_R _18577_ (.A1(_02974_),
    .A2(_02733_),
    .A3(_02991_),
    .B1(_02957_),
    .B2(_02992_),
    .Y(_02043_));
 NAND2x1_ASAP7_75t_R _18578_ (.A(_01001_),
    .B(_02950_),
    .Y(_02993_));
 OA21x2_ASAP7_75t_R _18579_ (.A1(_02816_),
    .A2(_02949_),
    .B(_02993_),
    .Y(_02044_));
 AND4x1_ASAP7_75t_R _18580_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_02955_),
    .Y(_02994_));
 INVx1_ASAP7_75t_R _18581_ (.A(_00070_),
    .Y(_02995_));
 AO32x1_ASAP7_75t_R _18582_ (.A1(_02974_),
    .A2(_02737_),
    .A3(_02994_),
    .B1(_02957_),
    .B2(_02995_),
    .Y(_02045_));
 AND3x1_ASAP7_75t_R _18583_ (.A(_02822_),
    .B(_02823_),
    .C(_02961_),
    .Y(_02996_));
 AO32x1_ASAP7_75t_R _18584_ (.A1(_02974_),
    .A2(_02740_),
    .A3(_02996_),
    .B1(_02957_),
    .B2(_03895_),
    .Y(_02046_));
 NAND2x1_ASAP7_75t_R _18585_ (.A(_00968_),
    .B(_02950_),
    .Y(_02997_));
 OA21x2_ASAP7_75t_R _18586_ (.A1(_02826_),
    .A2(_02949_),
    .B(_02997_),
    .Y(_02047_));
 NAND2x1_ASAP7_75t_R _18587_ (.A(_00935_),
    .B(_02950_),
    .Y(_02998_));
 OA21x2_ASAP7_75t_R _18588_ (.A1(_02828_),
    .A2(_02949_),
    .B(_02998_),
    .Y(_02048_));
 AND2x2_ASAP7_75t_R _18589_ (.A(_00901_),
    .B(_02957_),
    .Y(_02999_));
 AOI21x1_ASAP7_75t_R _18590_ (.A1(_02745_),
    .A2(_02956_),
    .B(_02999_),
    .Y(_02049_));
 NOR2x1_ASAP7_75t_R _18591_ (.A(_00868_),
    .B(_02956_),
    .Y(_03000_));
 AO21x1_ASAP7_75t_R _18592_ (.A1(_02831_),
    .A2(_02956_),
    .B(_03000_),
    .Y(_02050_));
 NOR2x1_ASAP7_75t_R _18593_ (.A(_00834_),
    .B(_02956_),
    .Y(_03001_));
 AO21x1_ASAP7_75t_R _18594_ (.A1(_02833_),
    .A2(_02956_),
    .B(_03001_),
    .Y(_02051_));
 NOR2x1_ASAP7_75t_R _18595_ (.A(_00801_),
    .B(_02956_),
    .Y(_03002_));
 AO21x1_ASAP7_75t_R _18596_ (.A1(_02835_),
    .A2(_02956_),
    .B(_03002_),
    .Y(_02052_));
 NAND2x1_ASAP7_75t_R _18597_ (.A(_00767_),
    .B(_02963_),
    .Y(_03003_));
 OA21x2_ASAP7_75t_R _18598_ (.A1(_02837_),
    .A2(_02949_),
    .B(_03003_),
    .Y(_02053_));
 AO21x1_ASAP7_75t_R _18599_ (.A1(_03566_),
    .A2(_07020_),
    .B(_09287_),
    .Y(_03004_));
 BUFx6f_ASAP7_75t_R _18600_ (.A(_03004_),
    .Y(_03005_));
 OR2x4_ASAP7_75t_R _18601_ (.A(_09289_),
    .B(_03005_),
    .Y(_03006_));
 BUFx4f_ASAP7_75t_R _18602_ (.A(_03006_),
    .Y(_03007_));
 BUFx6f_ASAP7_75t_R _18603_ (.A(_03006_),
    .Y(_03008_));
 NAND2x1_ASAP7_75t_R _18604_ (.A(_00004_),
    .B(_03008_),
    .Y(_03009_));
 OA21x2_ASAP7_75t_R _18605_ (.A1(_02672_),
    .A2(_03007_),
    .B(_03009_),
    .Y(_02054_));
 NAND2x1_ASAP7_75t_R _18606_ (.A(_00736_),
    .B(_03008_),
    .Y(_03010_));
 OA21x2_ASAP7_75t_R _18607_ (.A1(_02755_),
    .A2(_03007_),
    .B(_03010_),
    .Y(_02055_));
 NAND2x1_ASAP7_75t_R _18608_ (.A(_00703_),
    .B(_03008_),
    .Y(_03011_));
 OA21x2_ASAP7_75t_R _18609_ (.A1(_02757_),
    .A2(_03007_),
    .B(_03011_),
    .Y(_02056_));
 NAND2x1_ASAP7_75t_R _18610_ (.A(_00670_),
    .B(_03008_),
    .Y(_03012_));
 OA21x2_ASAP7_75t_R _18611_ (.A1(_02759_),
    .A2(_03007_),
    .B(_03012_),
    .Y(_02057_));
 NOR2x2_ASAP7_75t_R _18612_ (.A(_09289_),
    .B(_03005_),
    .Y(_03013_));
 BUFx4f_ASAP7_75t_R _18613_ (.A(_03013_),
    .Y(_03014_));
 BUFx4f_ASAP7_75t_R _18614_ (.A(_03006_),
    .Y(_03015_));
 AND2x2_ASAP7_75t_R _18615_ (.A(_00637_),
    .B(_03015_),
    .Y(_03016_));
 AOI21x1_ASAP7_75t_R _18616_ (.A1(_02682_),
    .A2(_03014_),
    .B(_03016_),
    .Y(_02058_));
 NAND2x1_ASAP7_75t_R _18617_ (.A(_00604_),
    .B(_03008_),
    .Y(_03017_));
 OA21x2_ASAP7_75t_R _18618_ (.A1(_02765_),
    .A2(_03007_),
    .B(_03017_),
    .Y(_02059_));
 AND2x2_ASAP7_75t_R _18619_ (.A(_00570_),
    .B(_03015_),
    .Y(_03018_));
 AOI21x1_ASAP7_75t_R _18620_ (.A1(_09769_),
    .A2(_03014_),
    .B(_03018_),
    .Y(_02060_));
 BUFx4f_ASAP7_75t_R _18621_ (.A(_03013_),
    .Y(_03019_));
 AND3x1_ASAP7_75t_R _18622_ (.A(_02768_),
    .B(_02769_),
    .C(_03019_),
    .Y(_03020_));
 BUFx4f_ASAP7_75t_R _18623_ (.A(_03006_),
    .Y(_03021_));
 INVx1_ASAP7_75t_R _18624_ (.A(_00537_),
    .Y(_03022_));
 AO32x1_ASAP7_75t_R _18625_ (.A1(_02688_),
    .A2(_02460_),
    .A3(_03020_),
    .B1(_03021_),
    .B2(_03022_),
    .Y(_02061_));
 BUFx4f_ASAP7_75t_R _18626_ (.A(_09547_),
    .Y(_03023_));
 AND2x2_ASAP7_75t_R _18627_ (.A(_02773_),
    .B(_03019_),
    .Y(_03024_));
 INVx1_ASAP7_75t_R _18628_ (.A(_00504_),
    .Y(_03025_));
 AO32x1_ASAP7_75t_R _18629_ (.A1(_03023_),
    .A2(_02693_),
    .A3(_03024_),
    .B1(_03021_),
    .B2(_03025_),
    .Y(_02062_));
 AND3x1_ASAP7_75t_R _18630_ (.A(_02776_),
    .B(_02777_),
    .C(_03019_),
    .Y(_03026_));
 INVx1_ASAP7_75t_R _18631_ (.A(_00471_),
    .Y(_03027_));
 AO32x1_ASAP7_75t_R _18632_ (.A1(_03023_),
    .A2(_02697_),
    .A3(_03026_),
    .B1(_03021_),
    .B2(_03027_),
    .Y(_02063_));
 AND3x1_ASAP7_75t_R _18633_ (.A(_02780_),
    .B(_02781_),
    .C(_03019_),
    .Y(_03028_));
 INVx1_ASAP7_75t_R _18634_ (.A(_00438_),
    .Y(_03029_));
 AO32x1_ASAP7_75t_R _18635_ (.A1(_03023_),
    .A2(_02700_),
    .A3(_03028_),
    .B1(_03021_),
    .B2(_03029_),
    .Y(_02064_));
 NAND2x1_ASAP7_75t_R _18636_ (.A(_01035_),
    .B(_03008_),
    .Y(_03030_));
 OA21x2_ASAP7_75t_R _18637_ (.A1(_02784_),
    .A2(_03007_),
    .B(_03030_),
    .Y(_02065_));
 AND2x2_ASAP7_75t_R _18638_ (.A(_02786_),
    .B(_03019_),
    .Y(_03031_));
 INVx1_ASAP7_75t_R _18639_ (.A(_00405_),
    .Y(_03032_));
 AO32x1_ASAP7_75t_R _18640_ (.A1(_03023_),
    .A2(_02704_),
    .A3(_03031_),
    .B1(_03021_),
    .B2(_03032_),
    .Y(_02066_));
 AND3x1_ASAP7_75t_R _18641_ (.A(_02789_),
    .B(_02790_),
    .C(_03019_),
    .Y(_03033_));
 INVx1_ASAP7_75t_R _18642_ (.A(_00372_),
    .Y(_03034_));
 AO32x1_ASAP7_75t_R _18643_ (.A1(_03023_),
    .A2(_02707_),
    .A3(_03033_),
    .B1(_03021_),
    .B2(_03034_),
    .Y(_02067_));
 AND2x2_ASAP7_75t_R _18644_ (.A(_02793_),
    .B(_03019_),
    .Y(_03035_));
 INVx1_ASAP7_75t_R _18645_ (.A(_00339_),
    .Y(_03036_));
 AO32x1_ASAP7_75t_R _18646_ (.A1(_03023_),
    .A2(_02710_),
    .A3(_03035_),
    .B1(_03021_),
    .B2(_03036_),
    .Y(_02068_));
 AND2x2_ASAP7_75t_R _18647_ (.A(_02796_),
    .B(_03019_),
    .Y(_03037_));
 INVx1_ASAP7_75t_R _18648_ (.A(_00305_),
    .Y(_03038_));
 AO32x1_ASAP7_75t_R _18649_ (.A1(_03023_),
    .A2(_02713_),
    .A3(_03037_),
    .B1(_03021_),
    .B2(_03038_),
    .Y(_02069_));
 AND2x2_ASAP7_75t_R _18650_ (.A(_02799_),
    .B(_03013_),
    .Y(_03039_));
 INVx1_ASAP7_75t_R _18651_ (.A(_00272_),
    .Y(_03040_));
 AO32x1_ASAP7_75t_R _18652_ (.A1(_03023_),
    .A2(_02716_),
    .A3(_03039_),
    .B1(_03021_),
    .B2(_03040_),
    .Y(_02070_));
 AND2x2_ASAP7_75t_R _18653_ (.A(_02802_),
    .B(_03013_),
    .Y(_03041_));
 INVx1_ASAP7_75t_R _18654_ (.A(_00239_),
    .Y(_03042_));
 AO32x1_ASAP7_75t_R _18655_ (.A1(_03023_),
    .A2(_02719_),
    .A3(_03041_),
    .B1(_03015_),
    .B2(_03042_),
    .Y(_02071_));
 NOR2x1_ASAP7_75t_R _18656_ (.A(_02723_),
    .B(_03015_),
    .Y(_03043_));
 INVx1_ASAP7_75t_R _18657_ (.A(_00206_),
    .Y(_03044_));
 AO32x1_ASAP7_75t_R _18658_ (.A1(_03023_),
    .A2(_02722_),
    .A3(_03043_),
    .B1(_03015_),
    .B2(_03044_),
    .Y(_02072_));
 INVx1_ASAP7_75t_R _18659_ (.A(_00172_),
    .Y(_03045_));
 AND2x2_ASAP7_75t_R _18660_ (.A(_02807_),
    .B(_03014_),
    .Y(_03046_));
 AO22x1_ASAP7_75t_R _18661_ (.A1(_03045_),
    .A2(_03008_),
    .B1(_03046_),
    .B2(_02728_),
    .Y(_02073_));
 BUFx4f_ASAP7_75t_R _18662_ (.A(_09547_),
    .Y(_03047_));
 AND4x1_ASAP7_75t_R _18663_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_03013_),
    .Y(_03048_));
 INVx1_ASAP7_75t_R _18664_ (.A(_00139_),
    .Y(_03049_));
 AO32x1_ASAP7_75t_R _18665_ (.A1(_03047_),
    .A2(_02730_),
    .A3(_03048_),
    .B1(_03015_),
    .B2(_03049_),
    .Y(_02074_));
 AND3x1_ASAP7_75t_R _18666_ (.A(_02813_),
    .B(_02814_),
    .C(_03019_),
    .Y(_03050_));
 INVx1_ASAP7_75t_R _18667_ (.A(_00105_),
    .Y(_03051_));
 AO32x1_ASAP7_75t_R _18668_ (.A1(_03047_),
    .A2(_02733_),
    .A3(_03050_),
    .B1(_03015_),
    .B2(_03051_),
    .Y(_02075_));
 NAND2x1_ASAP7_75t_R _18669_ (.A(_01002_),
    .B(_03008_),
    .Y(_03052_));
 OA21x2_ASAP7_75t_R _18670_ (.A1(_02816_),
    .A2(_03007_),
    .B(_03052_),
    .Y(_02076_));
 AND4x1_ASAP7_75t_R _18671_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_03013_),
    .Y(_03053_));
 INVx1_ASAP7_75t_R _18672_ (.A(_00071_),
    .Y(_03054_));
 AO32x1_ASAP7_75t_R _18673_ (.A1(_03047_),
    .A2(_02737_),
    .A3(_03053_),
    .B1(_03015_),
    .B2(_03054_),
    .Y(_02077_));
 AND3x1_ASAP7_75t_R _18674_ (.A(_02822_),
    .B(_02823_),
    .C(_03019_),
    .Y(_03055_));
 INVx1_ASAP7_75t_R _18675_ (.A(_00039_),
    .Y(_03056_));
 AO32x1_ASAP7_75t_R _18676_ (.A1(_03047_),
    .A2(_02740_),
    .A3(_03055_),
    .B1(_03015_),
    .B2(_03056_),
    .Y(_02078_));
 NAND2x1_ASAP7_75t_R _18677_ (.A(_00969_),
    .B(_03008_),
    .Y(_03057_));
 OA21x2_ASAP7_75t_R _18678_ (.A1(_02826_),
    .A2(_03007_),
    .B(_03057_),
    .Y(_02079_));
 NAND2x1_ASAP7_75t_R _18679_ (.A(_00936_),
    .B(_03008_),
    .Y(_03058_));
 OA21x2_ASAP7_75t_R _18680_ (.A1(_02828_),
    .A2(_03007_),
    .B(_03058_),
    .Y(_02080_));
 AND2x2_ASAP7_75t_R _18681_ (.A(_00902_),
    .B(_03015_),
    .Y(_03059_));
 AOI21x1_ASAP7_75t_R _18682_ (.A1(_02745_),
    .A2(_03014_),
    .B(_03059_),
    .Y(_02081_));
 NOR2x1_ASAP7_75t_R _18683_ (.A(_00869_),
    .B(_03014_),
    .Y(_03060_));
 AO21x1_ASAP7_75t_R _18684_ (.A1(_02831_),
    .A2(_03014_),
    .B(_03060_),
    .Y(_02082_));
 NOR2x1_ASAP7_75t_R _18685_ (.A(_00835_),
    .B(_03014_),
    .Y(_03061_));
 AO21x1_ASAP7_75t_R _18686_ (.A1(_02833_),
    .A2(_03014_),
    .B(_03061_),
    .Y(_02083_));
 NOR2x1_ASAP7_75t_R _18687_ (.A(_00802_),
    .B(_03014_),
    .Y(_03062_));
 AO21x1_ASAP7_75t_R _18688_ (.A1(_02835_),
    .A2(_03014_),
    .B(_03062_),
    .Y(_02084_));
 NAND2x1_ASAP7_75t_R _18689_ (.A(_00768_),
    .B(_03021_),
    .Y(_03063_));
 OA21x2_ASAP7_75t_R _18690_ (.A1(_02837_),
    .A2(_03007_),
    .B(_03063_),
    .Y(_02085_));
 OR3x4_ASAP7_75t_R _18691_ (.A(_07131_),
    .B(_09349_),
    .C(_03005_),
    .Y(_03064_));
 BUFx4f_ASAP7_75t_R _18692_ (.A(_03064_),
    .Y(_03065_));
 BUFx6f_ASAP7_75t_R _18693_ (.A(_03064_),
    .Y(_03066_));
 NAND2x1_ASAP7_75t_R _18694_ (.A(_00005_),
    .B(_03066_),
    .Y(_03067_));
 OA21x2_ASAP7_75t_R _18695_ (.A1(_02672_),
    .A2(_03065_),
    .B(_03067_),
    .Y(_02086_));
 NAND2x1_ASAP7_75t_R _18696_ (.A(_00737_),
    .B(_03066_),
    .Y(_03068_));
 OA21x2_ASAP7_75t_R _18697_ (.A1(_02755_),
    .A2(_03065_),
    .B(_03068_),
    .Y(_02087_));
 NAND2x1_ASAP7_75t_R _18698_ (.A(_00704_),
    .B(_03066_),
    .Y(_03069_));
 OA21x2_ASAP7_75t_R _18699_ (.A1(_02757_),
    .A2(_03065_),
    .B(_03069_),
    .Y(_02088_));
 NAND2x1_ASAP7_75t_R _18700_ (.A(_00671_),
    .B(_03066_),
    .Y(_03070_));
 OA21x2_ASAP7_75t_R _18701_ (.A1(_02759_),
    .A2(_03065_),
    .B(_03070_),
    .Y(_02089_));
 NOR2x2_ASAP7_75t_R _18702_ (.A(_09357_),
    .B(_03005_),
    .Y(_03071_));
 BUFx6f_ASAP7_75t_R _18703_ (.A(_03071_),
    .Y(_03072_));
 BUFx4f_ASAP7_75t_R _18704_ (.A(_03064_),
    .Y(_03073_));
 AND2x2_ASAP7_75t_R _18705_ (.A(_00638_),
    .B(_03073_),
    .Y(_03074_));
 AOI21x1_ASAP7_75t_R _18706_ (.A1(_02682_),
    .A2(_03072_),
    .B(_03074_),
    .Y(_02090_));
 NAND2x1_ASAP7_75t_R _18707_ (.A(_00605_),
    .B(_03066_),
    .Y(_03075_));
 OA21x2_ASAP7_75t_R _18708_ (.A1(_02765_),
    .A2(_03065_),
    .B(_03075_),
    .Y(_02091_));
 AND2x2_ASAP7_75t_R _18709_ (.A(_00571_),
    .B(_03073_),
    .Y(_03076_));
 AOI21x1_ASAP7_75t_R _18710_ (.A1(_09769_),
    .A2(_03072_),
    .B(_03076_),
    .Y(_02092_));
 BUFx4f_ASAP7_75t_R _18711_ (.A(_03071_),
    .Y(_03077_));
 AND3x1_ASAP7_75t_R _18712_ (.A(_02768_),
    .B(_02769_),
    .C(_03077_),
    .Y(_03078_));
 BUFx6f_ASAP7_75t_R _18713_ (.A(_03064_),
    .Y(_03079_));
 INVx1_ASAP7_75t_R _18714_ (.A(_00538_),
    .Y(_03080_));
 AO32x1_ASAP7_75t_R _18715_ (.A1(_02688_),
    .A2(_08798_),
    .A3(_03078_),
    .B1(_03079_),
    .B2(_03080_),
    .Y(_02093_));
 AND2x2_ASAP7_75t_R _18716_ (.A(_02773_),
    .B(_03077_),
    .Y(_03081_));
 INVx1_ASAP7_75t_R _18717_ (.A(_00505_),
    .Y(_03082_));
 AO32x1_ASAP7_75t_R _18718_ (.A1(_03047_),
    .A2(_02693_),
    .A3(_03081_),
    .B1(_03079_),
    .B2(_03082_),
    .Y(_02094_));
 AND3x1_ASAP7_75t_R _18719_ (.A(_02776_),
    .B(_02777_),
    .C(_03077_),
    .Y(_03083_));
 INVx1_ASAP7_75t_R _18720_ (.A(_00472_),
    .Y(_03084_));
 AO32x1_ASAP7_75t_R _18721_ (.A1(_03047_),
    .A2(_02697_),
    .A3(_03083_),
    .B1(_03079_),
    .B2(_03084_),
    .Y(_02095_));
 AND3x1_ASAP7_75t_R _18722_ (.A(_02780_),
    .B(_02781_),
    .C(_03077_),
    .Y(_03085_));
 INVx1_ASAP7_75t_R _18723_ (.A(_00439_),
    .Y(_03086_));
 AO32x1_ASAP7_75t_R _18724_ (.A1(_03047_),
    .A2(_02700_),
    .A3(_03085_),
    .B1(_03079_),
    .B2(_03086_),
    .Y(_02096_));
 NAND2x1_ASAP7_75t_R _18725_ (.A(_01036_),
    .B(_03066_),
    .Y(_03087_));
 OA21x2_ASAP7_75t_R _18726_ (.A1(_02784_),
    .A2(_03065_),
    .B(_03087_),
    .Y(_02097_));
 AND2x2_ASAP7_75t_R _18727_ (.A(_02786_),
    .B(_03077_),
    .Y(_03088_));
 INVx1_ASAP7_75t_R _18728_ (.A(_00406_),
    .Y(_03089_));
 AO32x1_ASAP7_75t_R _18729_ (.A1(_03047_),
    .A2(_02704_),
    .A3(_03088_),
    .B1(_03079_),
    .B2(_03089_),
    .Y(_02098_));
 AND3x1_ASAP7_75t_R _18730_ (.A(_02789_),
    .B(_02790_),
    .C(_03077_),
    .Y(_03090_));
 INVx1_ASAP7_75t_R _18731_ (.A(_00373_),
    .Y(_03091_));
 AO32x1_ASAP7_75t_R _18732_ (.A1(_03047_),
    .A2(_02707_),
    .A3(_03090_),
    .B1(_03079_),
    .B2(_03091_),
    .Y(_02099_));
 AND2x2_ASAP7_75t_R _18733_ (.A(_02793_),
    .B(_03077_),
    .Y(_03092_));
 INVx1_ASAP7_75t_R _18734_ (.A(_00340_),
    .Y(_03093_));
 AO32x1_ASAP7_75t_R _18735_ (.A1(_03047_),
    .A2(_02710_),
    .A3(_03092_),
    .B1(_03079_),
    .B2(_03093_),
    .Y(_02100_));
 BUFx4f_ASAP7_75t_R _18736_ (.A(_09547_),
    .Y(_03094_));
 AND2x2_ASAP7_75t_R _18737_ (.A(_02796_),
    .B(_03077_),
    .Y(_03095_));
 INVx1_ASAP7_75t_R _18738_ (.A(_00306_),
    .Y(_03096_));
 AO32x1_ASAP7_75t_R _18739_ (.A1(_03094_),
    .A2(_02713_),
    .A3(_03095_),
    .B1(_03079_),
    .B2(_03096_),
    .Y(_02101_));
 AND2x2_ASAP7_75t_R _18740_ (.A(_02799_),
    .B(_03071_),
    .Y(_03097_));
 INVx1_ASAP7_75t_R _18741_ (.A(_00273_),
    .Y(_03098_));
 AO32x1_ASAP7_75t_R _18742_ (.A1(_03094_),
    .A2(_02716_),
    .A3(_03097_),
    .B1(_03079_),
    .B2(_03098_),
    .Y(_02102_));
 AND2x2_ASAP7_75t_R _18743_ (.A(_02802_),
    .B(_03071_),
    .Y(_03099_));
 INVx1_ASAP7_75t_R _18744_ (.A(_00240_),
    .Y(_03100_));
 AO32x1_ASAP7_75t_R _18745_ (.A1(_03094_),
    .A2(_02719_),
    .A3(_03099_),
    .B1(_03073_),
    .B2(_03100_),
    .Y(_02103_));
 NOR2x1_ASAP7_75t_R _18746_ (.A(_02723_),
    .B(_03073_),
    .Y(_03101_));
 INVx1_ASAP7_75t_R _18747_ (.A(_00207_),
    .Y(_03102_));
 AO32x1_ASAP7_75t_R _18748_ (.A1(_03094_),
    .A2(_02722_),
    .A3(_03101_),
    .B1(_03073_),
    .B2(_03102_),
    .Y(_02104_));
 INVx1_ASAP7_75t_R _18749_ (.A(_00173_),
    .Y(_03103_));
 AND2x2_ASAP7_75t_R _18750_ (.A(_02807_),
    .B(_03072_),
    .Y(_03104_));
 AO22x1_ASAP7_75t_R _18751_ (.A1(_03103_),
    .A2(_03066_),
    .B1(_03104_),
    .B2(_02728_),
    .Y(_02105_));
 AND4x1_ASAP7_75t_R _18752_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_03071_),
    .Y(_03105_));
 INVx1_ASAP7_75t_R _18753_ (.A(_00140_),
    .Y(_03106_));
 AO32x1_ASAP7_75t_R _18754_ (.A1(_03094_),
    .A2(_02730_),
    .A3(_03105_),
    .B1(_03073_),
    .B2(_03106_),
    .Y(_02106_));
 AND3x1_ASAP7_75t_R _18755_ (.A(_02813_),
    .B(_02814_),
    .C(_03077_),
    .Y(_03107_));
 INVx1_ASAP7_75t_R _18756_ (.A(_00106_),
    .Y(_03108_));
 AO32x1_ASAP7_75t_R _18757_ (.A1(_03094_),
    .A2(_02733_),
    .A3(_03107_),
    .B1(_03073_),
    .B2(_03108_),
    .Y(_02107_));
 NAND2x1_ASAP7_75t_R _18758_ (.A(_01003_),
    .B(_03066_),
    .Y(_03109_));
 OA21x2_ASAP7_75t_R _18759_ (.A1(_02816_),
    .A2(_03065_),
    .B(_03109_),
    .Y(_02108_));
 AND4x1_ASAP7_75t_R _18760_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_03071_),
    .Y(_03110_));
 INVx1_ASAP7_75t_R _18761_ (.A(_00072_),
    .Y(_03111_));
 AO32x1_ASAP7_75t_R _18762_ (.A1(_03094_),
    .A2(_02737_),
    .A3(_03110_),
    .B1(_03073_),
    .B2(_03111_),
    .Y(_02109_));
 AND3x1_ASAP7_75t_R _18763_ (.A(_02822_),
    .B(_02823_),
    .C(_03077_),
    .Y(_03112_));
 INVx1_ASAP7_75t_R _18764_ (.A(_00040_),
    .Y(_03113_));
 AO32x1_ASAP7_75t_R _18765_ (.A1(_03094_),
    .A2(_02740_),
    .A3(_03112_),
    .B1(_03073_),
    .B2(_03113_),
    .Y(_02110_));
 NAND2x1_ASAP7_75t_R _18766_ (.A(_00970_),
    .B(_03066_),
    .Y(_03114_));
 OA21x2_ASAP7_75t_R _18767_ (.A1(_02826_),
    .A2(_03065_),
    .B(_03114_),
    .Y(_02111_));
 NAND2x1_ASAP7_75t_R _18768_ (.A(_00937_),
    .B(_03066_),
    .Y(_03115_));
 OA21x2_ASAP7_75t_R _18769_ (.A1(_02828_),
    .A2(_03065_),
    .B(_03115_),
    .Y(_02112_));
 AND2x2_ASAP7_75t_R _18770_ (.A(_00903_),
    .B(_03073_),
    .Y(_03116_));
 AOI21x1_ASAP7_75t_R _18771_ (.A1(_02745_),
    .A2(_03072_),
    .B(_03116_),
    .Y(_02113_));
 NOR2x1_ASAP7_75t_R _18772_ (.A(_00870_),
    .B(_03072_),
    .Y(_03117_));
 AO21x1_ASAP7_75t_R _18773_ (.A1(_02831_),
    .A2(_03072_),
    .B(_03117_),
    .Y(_02114_));
 NOR2x1_ASAP7_75t_R _18774_ (.A(_00836_),
    .B(_03072_),
    .Y(_03118_));
 AO21x1_ASAP7_75t_R _18775_ (.A1(_02833_),
    .A2(_03072_),
    .B(_03118_),
    .Y(_02115_));
 NOR2x1_ASAP7_75t_R _18776_ (.A(_00803_),
    .B(_03072_),
    .Y(_03119_));
 AO21x1_ASAP7_75t_R _18777_ (.A1(_02835_),
    .A2(_03072_),
    .B(_03119_),
    .Y(_02116_));
 NAND2x1_ASAP7_75t_R _18778_ (.A(_00769_),
    .B(_03079_),
    .Y(_03120_));
 OA21x2_ASAP7_75t_R _18779_ (.A1(_02837_),
    .A2(_03065_),
    .B(_03120_),
    .Y(_02117_));
 OR3x4_ASAP7_75t_R _18780_ (.A(_09408_),
    .B(_08601_),
    .C(_03005_),
    .Y(_03121_));
 BUFx4f_ASAP7_75t_R _18781_ (.A(_03121_),
    .Y(_03122_));
 BUFx6f_ASAP7_75t_R _18782_ (.A(_03121_),
    .Y(_03123_));
 NAND2x1_ASAP7_75t_R _18783_ (.A(_00006_),
    .B(_03123_),
    .Y(_03124_));
 OA21x2_ASAP7_75t_R _18784_ (.A1(_02672_),
    .A2(_03122_),
    .B(_03124_),
    .Y(_02118_));
 NAND2x1_ASAP7_75t_R _18785_ (.A(_00738_),
    .B(_03123_),
    .Y(_03125_));
 OA21x2_ASAP7_75t_R _18786_ (.A1(_02755_),
    .A2(_03122_),
    .B(_03125_),
    .Y(_02119_));
 NAND2x1_ASAP7_75t_R _18787_ (.A(_00705_),
    .B(_03123_),
    .Y(_03126_));
 OA21x2_ASAP7_75t_R _18788_ (.A1(_02757_),
    .A2(_03122_),
    .B(_03126_),
    .Y(_02120_));
 NAND2x1_ASAP7_75t_R _18789_ (.A(_00672_),
    .B(_03123_),
    .Y(_03127_));
 OA21x2_ASAP7_75t_R _18790_ (.A1(_02759_),
    .A2(_03122_),
    .B(_03127_),
    .Y(_02121_));
 NOR2x2_ASAP7_75t_R _18791_ (.A(_09416_),
    .B(_03005_),
    .Y(_03128_));
 BUFx6f_ASAP7_75t_R _18792_ (.A(_03128_),
    .Y(_03129_));
 BUFx4f_ASAP7_75t_R _18793_ (.A(_03121_),
    .Y(_03130_));
 AND2x2_ASAP7_75t_R _18794_ (.A(_00639_),
    .B(_03130_),
    .Y(_03131_));
 AOI21x1_ASAP7_75t_R _18795_ (.A1(_02682_),
    .A2(_03129_),
    .B(_03131_),
    .Y(_02122_));
 NAND2x1_ASAP7_75t_R _18796_ (.A(_00606_),
    .B(_03123_),
    .Y(_03132_));
 OA21x2_ASAP7_75t_R _18797_ (.A1(_02765_),
    .A2(_03122_),
    .B(_03132_),
    .Y(_02123_));
 OR2x2_ASAP7_75t_R _18798_ (.A(_00572_),
    .B(_03129_),
    .Y(_03133_));
 OAI21x1_ASAP7_75t_R _18799_ (.A1(_09937_),
    .A2(_03122_),
    .B(_03133_),
    .Y(_02124_));
 BUFx4f_ASAP7_75t_R _18800_ (.A(_03128_),
    .Y(_03134_));
 AND3x1_ASAP7_75t_R _18801_ (.A(_02768_),
    .B(_02769_),
    .C(_03134_),
    .Y(_03135_));
 BUFx6f_ASAP7_75t_R _18802_ (.A(_03121_),
    .Y(_03136_));
 AO32x1_ASAP7_75t_R _18803_ (.A1(_02688_),
    .A2(_08798_),
    .A3(_03135_),
    .B1(_03136_),
    .B2(_05699_),
    .Y(_02125_));
 AND2x2_ASAP7_75t_R _18804_ (.A(_02773_),
    .B(_03134_),
    .Y(_03137_));
 INVx1_ASAP7_75t_R _18805_ (.A(_00506_),
    .Y(_03138_));
 AO32x1_ASAP7_75t_R _18806_ (.A1(_03094_),
    .A2(_02693_),
    .A3(_03137_),
    .B1(_03136_),
    .B2(_03138_),
    .Y(_02126_));
 AND3x1_ASAP7_75t_R _18807_ (.A(_02776_),
    .B(_02777_),
    .C(_03134_),
    .Y(_03139_));
 INVx1_ASAP7_75t_R _18808_ (.A(_00473_),
    .Y(_03140_));
 AO32x1_ASAP7_75t_R _18809_ (.A1(_03094_),
    .A2(_02697_),
    .A3(_03139_),
    .B1(_03136_),
    .B2(_03140_),
    .Y(_02127_));
 BUFx4f_ASAP7_75t_R _18810_ (.A(_09547_),
    .Y(_03141_));
 AND3x1_ASAP7_75t_R _18811_ (.A(_02780_),
    .B(_02781_),
    .C(_03134_),
    .Y(_03142_));
 INVx1_ASAP7_75t_R _18812_ (.A(_00440_),
    .Y(_03143_));
 AO32x1_ASAP7_75t_R _18813_ (.A1(_03141_),
    .A2(_02700_),
    .A3(_03142_),
    .B1(_03136_),
    .B2(_03143_),
    .Y(_02128_));
 NAND2x1_ASAP7_75t_R _18814_ (.A(_01037_),
    .B(_03123_),
    .Y(_03144_));
 OA21x2_ASAP7_75t_R _18815_ (.A1(_02784_),
    .A2(_03122_),
    .B(_03144_),
    .Y(_02129_));
 AND2x2_ASAP7_75t_R _18816_ (.A(_02786_),
    .B(_03134_),
    .Y(_03145_));
 INVx1_ASAP7_75t_R _18817_ (.A(_00407_),
    .Y(_03146_));
 AO32x1_ASAP7_75t_R _18818_ (.A1(_03141_),
    .A2(_02704_),
    .A3(_03145_),
    .B1(_03136_),
    .B2(_03146_),
    .Y(_02130_));
 AND3x1_ASAP7_75t_R _18819_ (.A(_02789_),
    .B(_02790_),
    .C(_03134_),
    .Y(_03147_));
 INVx1_ASAP7_75t_R _18820_ (.A(_00374_),
    .Y(_03148_));
 AO32x1_ASAP7_75t_R _18821_ (.A1(_03141_),
    .A2(_02707_),
    .A3(_03147_),
    .B1(_03136_),
    .B2(_03148_),
    .Y(_02131_));
 AND2x2_ASAP7_75t_R _18822_ (.A(_02793_),
    .B(_03134_),
    .Y(_03149_));
 INVx1_ASAP7_75t_R _18823_ (.A(_00341_),
    .Y(_03150_));
 AO32x1_ASAP7_75t_R _18824_ (.A1(_03141_),
    .A2(_02710_),
    .A3(_03149_),
    .B1(_03136_),
    .B2(_03150_),
    .Y(_02132_));
 AND2x2_ASAP7_75t_R _18825_ (.A(_02796_),
    .B(_03134_),
    .Y(_03151_));
 INVx1_ASAP7_75t_R _18826_ (.A(_00307_),
    .Y(_03152_));
 AO32x1_ASAP7_75t_R _18827_ (.A1(_03141_),
    .A2(_02713_),
    .A3(_03151_),
    .B1(_03136_),
    .B2(_03152_),
    .Y(_02133_));
 AND2x2_ASAP7_75t_R _18828_ (.A(_02799_),
    .B(_03128_),
    .Y(_03153_));
 INVx1_ASAP7_75t_R _18829_ (.A(_00274_),
    .Y(_03154_));
 AO32x1_ASAP7_75t_R _18830_ (.A1(_03141_),
    .A2(_02716_),
    .A3(_03153_),
    .B1(_03130_),
    .B2(_03154_),
    .Y(_02134_));
 AND2x2_ASAP7_75t_R _18831_ (.A(_02802_),
    .B(_03128_),
    .Y(_03155_));
 INVx1_ASAP7_75t_R _18832_ (.A(_00241_),
    .Y(_03156_));
 AO32x1_ASAP7_75t_R _18833_ (.A1(_03141_),
    .A2(_02719_),
    .A3(_03155_),
    .B1(_03130_),
    .B2(_03156_),
    .Y(_02135_));
 NOR2x1_ASAP7_75t_R _18834_ (.A(_02723_),
    .B(_03130_),
    .Y(_03157_));
 AO32x1_ASAP7_75t_R _18835_ (.A1(_03141_),
    .A2(_02722_),
    .A3(_03157_),
    .B1(_03130_),
    .B2(_04723_),
    .Y(_02136_));
 INVx1_ASAP7_75t_R _18836_ (.A(_00174_),
    .Y(_03158_));
 AND2x2_ASAP7_75t_R _18837_ (.A(_02807_),
    .B(_03129_),
    .Y(_03159_));
 AO22x1_ASAP7_75t_R _18838_ (.A1(_03158_),
    .A2(_03123_),
    .B1(_03159_),
    .B2(_02728_),
    .Y(_02137_));
 AND4x1_ASAP7_75t_R _18839_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_03128_),
    .Y(_03160_));
 INVx1_ASAP7_75t_R _18840_ (.A(_00141_),
    .Y(_03161_));
 AO32x1_ASAP7_75t_R _18841_ (.A1(_03141_),
    .A2(_02730_),
    .A3(_03160_),
    .B1(_03130_),
    .B2(_03161_),
    .Y(_02138_));
 AND3x1_ASAP7_75t_R _18842_ (.A(_02813_),
    .B(_02814_),
    .C(_03134_),
    .Y(_03162_));
 INVx1_ASAP7_75t_R _18843_ (.A(_00107_),
    .Y(_03163_));
 AO32x1_ASAP7_75t_R _18844_ (.A1(_03141_),
    .A2(_02733_),
    .A3(_03162_),
    .B1(_03130_),
    .B2(_03163_),
    .Y(_02139_));
 NAND2x1_ASAP7_75t_R _18845_ (.A(_01004_),
    .B(_03123_),
    .Y(_03164_));
 OA21x2_ASAP7_75t_R _18846_ (.A1(_02816_),
    .A2(_03122_),
    .B(_03164_),
    .Y(_02140_));
 BUFx4f_ASAP7_75t_R _18847_ (.A(_09547_),
    .Y(_03165_));
 AND4x1_ASAP7_75t_R _18848_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_03128_),
    .Y(_03166_));
 INVx1_ASAP7_75t_R _18849_ (.A(_00073_),
    .Y(_03167_));
 AO32x1_ASAP7_75t_R _18850_ (.A1(_03165_),
    .A2(_02737_),
    .A3(_03166_),
    .B1(_03130_),
    .B2(_03167_),
    .Y(_02141_));
 AND3x1_ASAP7_75t_R _18851_ (.A(_02822_),
    .B(_02823_),
    .C(_03134_),
    .Y(_03168_));
 INVx1_ASAP7_75t_R _18852_ (.A(_00041_),
    .Y(_03169_));
 AO32x1_ASAP7_75t_R _18853_ (.A1(_03165_),
    .A2(_02740_),
    .A3(_03168_),
    .B1(_03130_),
    .B2(_03169_),
    .Y(_02142_));
 NAND2x1_ASAP7_75t_R _18854_ (.A(_00971_),
    .B(_03123_),
    .Y(_03170_));
 OA21x2_ASAP7_75t_R _18855_ (.A1(_02826_),
    .A2(_03122_),
    .B(_03170_),
    .Y(_02143_));
 NAND2x1_ASAP7_75t_R _18856_ (.A(_00938_),
    .B(_03136_),
    .Y(_03171_));
 OA21x2_ASAP7_75t_R _18857_ (.A1(_02828_),
    .A2(_03122_),
    .B(_03171_),
    .Y(_02144_));
 AND2x2_ASAP7_75t_R _18858_ (.A(_00904_),
    .B(_03130_),
    .Y(_03172_));
 AOI21x1_ASAP7_75t_R _18859_ (.A1(_02745_),
    .A2(_03129_),
    .B(_03172_),
    .Y(_02145_));
 NOR2x1_ASAP7_75t_R _18860_ (.A(_00871_),
    .B(_03129_),
    .Y(_03173_));
 AO21x1_ASAP7_75t_R _18861_ (.A1(_02831_),
    .A2(_03129_),
    .B(_03173_),
    .Y(_02146_));
 NOR2x1_ASAP7_75t_R _18862_ (.A(_00837_),
    .B(_03129_),
    .Y(_03174_));
 AO21x1_ASAP7_75t_R _18863_ (.A1(_02833_),
    .A2(_03129_),
    .B(_03174_),
    .Y(_02147_));
 NOR2x1_ASAP7_75t_R _18864_ (.A(_00804_),
    .B(_03129_),
    .Y(_03175_));
 AO21x1_ASAP7_75t_R _18865_ (.A1(_02835_),
    .A2(_03129_),
    .B(_03175_),
    .Y(_02148_));
 NAND2x1_ASAP7_75t_R _18866_ (.A(_00770_),
    .B(_03136_),
    .Y(_03176_));
 OA21x2_ASAP7_75t_R _18867_ (.A1(_02837_),
    .A2(_03123_),
    .B(_03176_),
    .Y(_02149_));
 OR3x4_ASAP7_75t_R _18868_ (.A(_09408_),
    .B(_09349_),
    .C(_03005_),
    .Y(_03177_));
 BUFx4f_ASAP7_75t_R _18869_ (.A(_03177_),
    .Y(_03178_));
 BUFx6f_ASAP7_75t_R _18870_ (.A(_03177_),
    .Y(_03179_));
 NAND2x1_ASAP7_75t_R _18871_ (.A(_00007_),
    .B(_03179_),
    .Y(_03180_));
 OA21x2_ASAP7_75t_R _18872_ (.A1(_02672_),
    .A2(_03178_),
    .B(_03180_),
    .Y(_02150_));
 NAND2x1_ASAP7_75t_R _18873_ (.A(_00739_),
    .B(_03179_),
    .Y(_03181_));
 OA21x2_ASAP7_75t_R _18874_ (.A1(_02755_),
    .A2(_03178_),
    .B(_03181_),
    .Y(_02151_));
 NAND2x1_ASAP7_75t_R _18875_ (.A(_00706_),
    .B(_03179_),
    .Y(_03182_));
 OA21x2_ASAP7_75t_R _18876_ (.A1(_02757_),
    .A2(_03178_),
    .B(_03182_),
    .Y(_02152_));
 NAND2x1_ASAP7_75t_R _18877_ (.A(_00673_),
    .B(_03179_),
    .Y(_03183_));
 OA21x2_ASAP7_75t_R _18878_ (.A1(_02759_),
    .A2(_03178_),
    .B(_03183_),
    .Y(_02153_));
 NOR2x2_ASAP7_75t_R _18879_ (.A(_09473_),
    .B(_03005_),
    .Y(_03184_));
 BUFx4f_ASAP7_75t_R _18880_ (.A(_03184_),
    .Y(_03185_));
 BUFx4f_ASAP7_75t_R _18881_ (.A(_03177_),
    .Y(_03186_));
 AND2x2_ASAP7_75t_R _18882_ (.A(_00640_),
    .B(_03186_),
    .Y(_03187_));
 AOI21x1_ASAP7_75t_R _18883_ (.A1(_02682_),
    .A2(_03185_),
    .B(_03187_),
    .Y(_02154_));
 NAND2x1_ASAP7_75t_R _18884_ (.A(_00607_),
    .B(_03179_),
    .Y(_03188_));
 OA21x2_ASAP7_75t_R _18885_ (.A1(_02765_),
    .A2(_03178_),
    .B(_03188_),
    .Y(_02155_));
 AND2x2_ASAP7_75t_R _18886_ (.A(_00573_),
    .B(_03186_),
    .Y(_03189_));
 AOI21x1_ASAP7_75t_R _18887_ (.A1(_08765_),
    .A2(_03185_),
    .B(_03189_),
    .Y(_02156_));
 BUFx4f_ASAP7_75t_R _18888_ (.A(_03184_),
    .Y(_03190_));
 AND3x1_ASAP7_75t_R _18889_ (.A(_02768_),
    .B(_02769_),
    .C(_03190_),
    .Y(_03191_));
 BUFx6f_ASAP7_75t_R _18890_ (.A(_03177_),
    .Y(_03192_));
 AO32x1_ASAP7_75t_R _18891_ (.A1(_02688_),
    .A2(_08798_),
    .A3(_03191_),
    .B1(_03192_),
    .B2(_05700_),
    .Y(_02157_));
 AND2x2_ASAP7_75t_R _18892_ (.A(_02773_),
    .B(_03190_),
    .Y(_03193_));
 INVx1_ASAP7_75t_R _18893_ (.A(_00507_),
    .Y(_03194_));
 AO32x1_ASAP7_75t_R _18894_ (.A1(_03165_),
    .A2(_02693_),
    .A3(_03193_),
    .B1(_03192_),
    .B2(_03194_),
    .Y(_02158_));
 AND3x1_ASAP7_75t_R _18895_ (.A(_02776_),
    .B(_02777_),
    .C(_03190_),
    .Y(_03195_));
 INVx1_ASAP7_75t_R _18896_ (.A(_00474_),
    .Y(_03196_));
 AO32x1_ASAP7_75t_R _18897_ (.A1(_03165_),
    .A2(_02697_),
    .A3(_03195_),
    .B1(_03192_),
    .B2(_03196_),
    .Y(_02159_));
 AND3x1_ASAP7_75t_R _18898_ (.A(_02780_),
    .B(_02781_),
    .C(_03190_),
    .Y(_03197_));
 INVx1_ASAP7_75t_R _18899_ (.A(_00441_),
    .Y(_03198_));
 AO32x1_ASAP7_75t_R _18900_ (.A1(_03165_),
    .A2(_02700_),
    .A3(_03197_),
    .B1(_03192_),
    .B2(_03198_),
    .Y(_02160_));
 NAND2x1_ASAP7_75t_R _18901_ (.A(_01038_),
    .B(_03179_),
    .Y(_03199_));
 OA21x2_ASAP7_75t_R _18902_ (.A1(_02784_),
    .A2(_03178_),
    .B(_03199_),
    .Y(_02161_));
 AND2x2_ASAP7_75t_R _18903_ (.A(_02786_),
    .B(_03190_),
    .Y(_03200_));
 INVx1_ASAP7_75t_R _18904_ (.A(_00408_),
    .Y(_03201_));
 AO32x1_ASAP7_75t_R _18905_ (.A1(_03165_),
    .A2(_02704_),
    .A3(_03200_),
    .B1(_03192_),
    .B2(_03201_),
    .Y(_02162_));
 AND3x1_ASAP7_75t_R _18906_ (.A(_02789_),
    .B(_02790_),
    .C(_03190_),
    .Y(_03202_));
 INVx1_ASAP7_75t_R _18907_ (.A(_00375_),
    .Y(_03203_));
 AO32x1_ASAP7_75t_R _18908_ (.A1(_03165_),
    .A2(_02707_),
    .A3(_03202_),
    .B1(_03192_),
    .B2(_03203_),
    .Y(_02163_));
 AND2x2_ASAP7_75t_R _18909_ (.A(_02793_),
    .B(_03190_),
    .Y(_03204_));
 INVx1_ASAP7_75t_R _18910_ (.A(_00342_),
    .Y(_03205_));
 AO32x1_ASAP7_75t_R _18911_ (.A1(_03165_),
    .A2(_02710_),
    .A3(_03204_),
    .B1(_03192_),
    .B2(_03205_),
    .Y(_02164_));
 AND2x2_ASAP7_75t_R _18912_ (.A(_02796_),
    .B(_03190_),
    .Y(_03206_));
 INVx1_ASAP7_75t_R _18913_ (.A(_00308_),
    .Y(_03207_));
 AO32x1_ASAP7_75t_R _18914_ (.A1(_03165_),
    .A2(_02713_),
    .A3(_03206_),
    .B1(_03192_),
    .B2(_03207_),
    .Y(_02165_));
 AND2x2_ASAP7_75t_R _18915_ (.A(_02799_),
    .B(_03184_),
    .Y(_03208_));
 INVx1_ASAP7_75t_R _18916_ (.A(_00275_),
    .Y(_03209_));
 AO32x1_ASAP7_75t_R _18917_ (.A1(_03165_),
    .A2(_02716_),
    .A3(_03208_),
    .B1(_03192_),
    .B2(_03209_),
    .Y(_02166_));
 BUFx4f_ASAP7_75t_R _18918_ (.A(_09547_),
    .Y(_03210_));
 AND2x2_ASAP7_75t_R _18919_ (.A(_02802_),
    .B(_03184_),
    .Y(_03211_));
 INVx1_ASAP7_75t_R _18920_ (.A(_00242_),
    .Y(_03212_));
 AO32x1_ASAP7_75t_R _18921_ (.A1(_03210_),
    .A2(_02719_),
    .A3(_03211_),
    .B1(_03186_),
    .B2(_03212_),
    .Y(_02167_));
 NOR2x1_ASAP7_75t_R _18922_ (.A(_02723_),
    .B(_03186_),
    .Y(_03213_));
 AO32x1_ASAP7_75t_R _18923_ (.A1(_03210_),
    .A2(_02722_),
    .A3(_03213_),
    .B1(_03186_),
    .B2(_04724_),
    .Y(_02168_));
 INVx1_ASAP7_75t_R _18924_ (.A(_00175_),
    .Y(_03214_));
 AND2x2_ASAP7_75t_R _18925_ (.A(_02807_),
    .B(_03185_),
    .Y(_03215_));
 AO22x1_ASAP7_75t_R _18926_ (.A1(_03214_),
    .A2(_03179_),
    .B1(_03215_),
    .B2(_02728_),
    .Y(_02169_));
 AND4x1_ASAP7_75t_R _18927_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_03184_),
    .Y(_03216_));
 INVx1_ASAP7_75t_R _18928_ (.A(_00142_),
    .Y(_03217_));
 AO32x1_ASAP7_75t_R _18929_ (.A1(_03210_),
    .A2(_02730_),
    .A3(_03216_),
    .B1(_03186_),
    .B2(_03217_),
    .Y(_02170_));
 AND3x1_ASAP7_75t_R _18930_ (.A(_02813_),
    .B(_02814_),
    .C(_03190_),
    .Y(_03218_));
 INVx1_ASAP7_75t_R _18931_ (.A(_00108_),
    .Y(_03219_));
 AO32x1_ASAP7_75t_R _18932_ (.A1(_03210_),
    .A2(_02733_),
    .A3(_03218_),
    .B1(_03186_),
    .B2(_03219_),
    .Y(_02171_));
 NAND2x1_ASAP7_75t_R _18933_ (.A(_01005_),
    .B(_03179_),
    .Y(_03220_));
 OA21x2_ASAP7_75t_R _18934_ (.A1(_02816_),
    .A2(_03178_),
    .B(_03220_),
    .Y(_02172_));
 AND4x1_ASAP7_75t_R _18935_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_03184_),
    .Y(_03221_));
 INVx1_ASAP7_75t_R _18936_ (.A(_00074_),
    .Y(_03222_));
 AO32x1_ASAP7_75t_R _18937_ (.A1(_03210_),
    .A2(_02737_),
    .A3(_03221_),
    .B1(_03186_),
    .B2(_03222_),
    .Y(_02173_));
 AND3x1_ASAP7_75t_R _18938_ (.A(_02822_),
    .B(_02823_),
    .C(_03190_),
    .Y(_03223_));
 INVx1_ASAP7_75t_R _18939_ (.A(_00042_),
    .Y(_03224_));
 AO32x1_ASAP7_75t_R _18940_ (.A1(_03210_),
    .A2(_02740_),
    .A3(_03223_),
    .B1(_03186_),
    .B2(_03224_),
    .Y(_02174_));
 NAND2x1_ASAP7_75t_R _18941_ (.A(_00972_),
    .B(_03179_),
    .Y(_03225_));
 OA21x2_ASAP7_75t_R _18942_ (.A1(_02826_),
    .A2(_03178_),
    .B(_03225_),
    .Y(_02175_));
 NAND2x1_ASAP7_75t_R _18943_ (.A(_00939_),
    .B(_03179_),
    .Y(_03226_));
 OA21x2_ASAP7_75t_R _18944_ (.A1(_02828_),
    .A2(_03178_),
    .B(_03226_),
    .Y(_02176_));
 AND2x2_ASAP7_75t_R _18945_ (.A(_00905_),
    .B(_03186_),
    .Y(_03227_));
 AOI21x1_ASAP7_75t_R _18946_ (.A1(_02745_),
    .A2(_03185_),
    .B(_03227_),
    .Y(_02177_));
 NOR2x1_ASAP7_75t_R _18947_ (.A(_00872_),
    .B(_03185_),
    .Y(_03228_));
 AO21x1_ASAP7_75t_R _18948_ (.A1(_02831_),
    .A2(_03185_),
    .B(_03228_),
    .Y(_02178_));
 NOR2x1_ASAP7_75t_R _18949_ (.A(_00838_),
    .B(_03185_),
    .Y(_03229_));
 AO21x1_ASAP7_75t_R _18950_ (.A1(_02833_),
    .A2(_03185_),
    .B(_03229_),
    .Y(_02179_));
 NOR2x1_ASAP7_75t_R _18951_ (.A(_00805_),
    .B(_03185_),
    .Y(_03230_));
 AO21x1_ASAP7_75t_R _18952_ (.A1(_02835_),
    .A2(_03185_),
    .B(_03230_),
    .Y(_02180_));
 NAND2x1_ASAP7_75t_R _18953_ (.A(_00771_),
    .B(_03192_),
    .Y(_03231_));
 OA21x2_ASAP7_75t_R _18954_ (.A1(_02837_),
    .A2(_03178_),
    .B(_03231_),
    .Y(_02181_));
 NAND2x2_ASAP7_75t_R _18955_ (.A(_08607_),
    .B(_09528_),
    .Y(_03232_));
 BUFx6f_ASAP7_75t_R _18956_ (.A(_03232_),
    .Y(_03233_));
 AO21x1_ASAP7_75t_R _18957_ (.A1(_09208_),
    .A2(_09529_),
    .B(_03693_),
    .Y(_03234_));
 OA21x2_ASAP7_75t_R _18958_ (.A1(_02672_),
    .A2(_03233_),
    .B(_03234_),
    .Y(_02182_));
 AO21x1_ASAP7_75t_R _18959_ (.A1(_09208_),
    .A2(_09529_),
    .B(_06320_),
    .Y(_03235_));
 OA21x2_ASAP7_75t_R _18960_ (.A1(_02755_),
    .A2(_03233_),
    .B(_03235_),
    .Y(_02183_));
 AO21x1_ASAP7_75t_R _18961_ (.A1(_09208_),
    .A2(_09529_),
    .B(_06196_),
    .Y(_03236_));
 OA21x2_ASAP7_75t_R _18962_ (.A1(_02757_),
    .A2(_03233_),
    .B(_03236_),
    .Y(_02184_));
 BUFx12f_ASAP7_75t_R _18963_ (.A(_03232_),
    .Y(_03237_));
 NAND2x1_ASAP7_75t_R _18964_ (.A(_00674_),
    .B(_03237_),
    .Y(_03238_));
 OA21x2_ASAP7_75t_R _18965_ (.A1(_02759_),
    .A2(_03233_),
    .B(_03238_),
    .Y(_02185_));
 AND2x2_ASAP7_75t_R _18966_ (.A(_08606_),
    .B(_09528_),
    .Y(_03239_));
 BUFx10_ASAP7_75t_R _18967_ (.A(_03239_),
    .Y(_03240_));
 AND2x2_ASAP7_75t_R _18968_ (.A(_00641_),
    .B(_03232_),
    .Y(_03241_));
 AOI21x1_ASAP7_75t_R _18969_ (.A1(_02682_),
    .A2(_03240_),
    .B(_03241_),
    .Y(_02186_));
 AO21x1_ASAP7_75t_R _18970_ (.A1(_09208_),
    .A2(_09529_),
    .B(_05933_),
    .Y(_03242_));
 OA21x2_ASAP7_75t_R _18971_ (.A1(_02765_),
    .A2(_03233_),
    .B(_03242_),
    .Y(_02187_));
 AO21x1_ASAP7_75t_R _18972_ (.A1(_09208_),
    .A2(_09543_),
    .B(_00574_),
    .Y(_03243_));
 OAI21x1_ASAP7_75t_R _18973_ (.A1(_09937_),
    .A2(_03233_),
    .B(_03243_),
    .Y(_02188_));
 AND3x1_ASAP7_75t_R _18974_ (.A(_02768_),
    .B(_02769_),
    .C(_03240_),
    .Y(_03244_));
 INVx1_ASAP7_75t_R _18975_ (.A(_00541_),
    .Y(_03245_));
 AO32x1_ASAP7_75t_R _18976_ (.A1(_02688_),
    .A2(_08798_),
    .A3(_03244_),
    .B1(_03237_),
    .B2(_03245_),
    .Y(_02189_));
 BUFx4f_ASAP7_75t_R _18977_ (.A(_03239_),
    .Y(_03246_));
 AND2x2_ASAP7_75t_R _18978_ (.A(_02773_),
    .B(_03246_),
    .Y(_03247_));
 AO32x1_ASAP7_75t_R _18979_ (.A1(_03210_),
    .A2(_02693_),
    .A3(_03247_),
    .B1(_03237_),
    .B2(_05604_),
    .Y(_02190_));
 AND3x1_ASAP7_75t_R _18980_ (.A(_02776_),
    .B(_02777_),
    .C(_03240_),
    .Y(_03248_));
 AO32x1_ASAP7_75t_R _18981_ (.A1(_03210_),
    .A2(_02697_),
    .A3(_03248_),
    .B1(_03237_),
    .B2(_05530_),
    .Y(_02191_));
 AND3x1_ASAP7_75t_R _18982_ (.A(_02780_),
    .B(_02781_),
    .C(_03240_),
    .Y(_03249_));
 AO32x1_ASAP7_75t_R _18983_ (.A1(_03210_),
    .A2(_02700_),
    .A3(_03249_),
    .B1(_03237_),
    .B2(_05439_),
    .Y(_02192_));
 NAND2x1_ASAP7_75t_R _18984_ (.A(_01039_),
    .B(_03237_),
    .Y(_03250_));
 OA21x2_ASAP7_75t_R _18985_ (.A1(_02784_),
    .A2(_03233_),
    .B(_03250_),
    .Y(_02193_));
 AND2x2_ASAP7_75t_R _18986_ (.A(_02786_),
    .B(_03246_),
    .Y(_03251_));
 BUFx4f_ASAP7_75t_R _18987_ (.A(_03232_),
    .Y(_03252_));
 AO32x1_ASAP7_75t_R _18988_ (.A1(_03210_),
    .A2(_02704_),
    .A3(_03251_),
    .B1(_03252_),
    .B2(_05330_),
    .Y(_02194_));
 BUFx4f_ASAP7_75t_R _18989_ (.A(_09547_),
    .Y(_03253_));
 AND3x1_ASAP7_75t_R _18990_ (.A(_02789_),
    .B(_02790_),
    .C(_03240_),
    .Y(_03254_));
 AO32x1_ASAP7_75t_R _18991_ (.A1(_03253_),
    .A2(_02707_),
    .A3(_03254_),
    .B1(_03252_),
    .B2(_05239_),
    .Y(_02195_));
 AND2x2_ASAP7_75t_R _18992_ (.A(_02793_),
    .B(_03246_),
    .Y(_03255_));
 AO32x1_ASAP7_75t_R _18993_ (.A1(_03253_),
    .A2(_02710_),
    .A3(_03255_),
    .B1(_03252_),
    .B2(_05132_),
    .Y(_02196_));
 AND2x2_ASAP7_75t_R _18994_ (.A(_02796_),
    .B(_03246_),
    .Y(_03256_));
 AO32x1_ASAP7_75t_R _18995_ (.A1(_03253_),
    .A2(_02713_),
    .A3(_03256_),
    .B1(_03252_),
    .B2(_05042_),
    .Y(_02197_));
 AND2x2_ASAP7_75t_R _18996_ (.A(_02799_),
    .B(_03246_),
    .Y(_03257_));
 AO32x1_ASAP7_75t_R _18997_ (.A1(_03253_),
    .A2(_02716_),
    .A3(_03257_),
    .B1(_03252_),
    .B2(_04933_),
    .Y(_02198_));
 AND2x2_ASAP7_75t_R _18998_ (.A(_02802_),
    .B(_03246_),
    .Y(_03258_));
 AO32x1_ASAP7_75t_R _18999_ (.A1(_03253_),
    .A2(_02719_),
    .A3(_03258_),
    .B1(_03252_),
    .B2(_04840_),
    .Y(_02199_));
 NOR2x1_ASAP7_75t_R _19000_ (.A(_02723_),
    .B(_03232_),
    .Y(_03259_));
 AO32x1_ASAP7_75t_R _19001_ (.A1(_03253_),
    .A2(_02722_),
    .A3(_03259_),
    .B1(_03252_),
    .B2(_04716_),
    .Y(_02200_));
 AND2x2_ASAP7_75t_R _19002_ (.A(_02807_),
    .B(_03240_),
    .Y(_03260_));
 AO22x1_ASAP7_75t_R _19003_ (.A1(_04608_),
    .A2(_03237_),
    .B1(_03260_),
    .B2(_02728_),
    .Y(_02201_));
 AND4x1_ASAP7_75t_R _19004_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_03246_),
    .Y(_03261_));
 INVx1_ASAP7_75t_R _19005_ (.A(_00143_),
    .Y(_03262_));
 AO32x1_ASAP7_75t_R _19006_ (.A1(_03253_),
    .A2(_02730_),
    .A3(_03261_),
    .B1(_03252_),
    .B2(_03262_),
    .Y(_02202_));
 AND3x1_ASAP7_75t_R _19007_ (.A(_02813_),
    .B(_02814_),
    .C(_03246_),
    .Y(_03263_));
 AO32x1_ASAP7_75t_R _19008_ (.A1(_03253_),
    .A2(_02733_),
    .A3(_03263_),
    .B1(_03252_),
    .B2(_04353_),
    .Y(_02203_));
 AO21x1_ASAP7_75t_R _19009_ (.A1(_09208_),
    .A2(_09529_),
    .B(_07082_),
    .Y(_03264_));
 OA21x2_ASAP7_75t_R _19010_ (.A1(_02816_),
    .A2(_03233_),
    .B(_03264_),
    .Y(_02204_));
 AND4x1_ASAP7_75t_R _19011_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_03246_),
    .Y(_03265_));
 AO32x1_ASAP7_75t_R _19012_ (.A1(_03253_),
    .A2(_02737_),
    .A3(_03265_),
    .B1(_03252_),
    .B2(_04203_),
    .Y(_02205_));
 AND3x1_ASAP7_75t_R _19013_ (.A(_02822_),
    .B(_02823_),
    .C(_03246_),
    .Y(_03266_));
 INVx1_ASAP7_75t_R _19014_ (.A(_00043_),
    .Y(_03267_));
 AO32x1_ASAP7_75t_R _19015_ (.A1(_03253_),
    .A2(_02740_),
    .A3(_03266_),
    .B1(_03232_),
    .B2(_03267_),
    .Y(_02206_));
 NAND2x1_ASAP7_75t_R _19016_ (.A(_00973_),
    .B(_03237_),
    .Y(_03268_));
 OA21x2_ASAP7_75t_R _19017_ (.A1(_02826_),
    .A2(_03233_),
    .B(_03268_),
    .Y(_02207_));
 NAND2x1_ASAP7_75t_R _19018_ (.A(_00940_),
    .B(_03237_),
    .Y(_03269_));
 OA21x2_ASAP7_75t_R _19019_ (.A1(_02828_),
    .A2(_03233_),
    .B(_03269_),
    .Y(_02208_));
 AND2x2_ASAP7_75t_R _19020_ (.A(_00906_),
    .B(_03232_),
    .Y(_03270_));
 AOI21x1_ASAP7_75t_R _19021_ (.A1(_02745_),
    .A2(_03240_),
    .B(_03270_),
    .Y(_02209_));
 AND2x2_ASAP7_75t_R _19022_ (.A(_06685_),
    .B(_03232_),
    .Y(_03271_));
 AO21x1_ASAP7_75t_R _19023_ (.A1(_02831_),
    .A2(_03240_),
    .B(_03271_),
    .Y(_02210_));
 AND2x2_ASAP7_75t_R _19024_ (.A(_06579_),
    .B(_03232_),
    .Y(_03272_));
 AO21x1_ASAP7_75t_R _19025_ (.A1(_02833_),
    .A2(_03240_),
    .B(_03272_),
    .Y(_02211_));
 AND2x2_ASAP7_75t_R _19026_ (.A(_06507_),
    .B(_03232_),
    .Y(_03273_));
 AO21x1_ASAP7_75t_R _19027_ (.A1(_02835_),
    .A2(_03240_),
    .B(_03273_),
    .Y(_02212_));
 AO21x1_ASAP7_75t_R _19028_ (.A1(_09208_),
    .A2(_09529_),
    .B(_06413_),
    .Y(_03274_));
 OA21x2_ASAP7_75t_R _19029_ (.A1(_02837_),
    .A2(_03237_),
    .B(_03274_),
    .Y(_02213_));
 NAND2x2_ASAP7_75t_R _19030_ (.A(_08607_),
    .B(_09590_),
    .Y(_03275_));
 BUFx6f_ASAP7_75t_R _19031_ (.A(_03275_),
    .Y(_03276_));
 AO21x1_ASAP7_75t_R _19032_ (.A1(_09208_),
    .A2(_09590_),
    .B(_03682_),
    .Y(_03277_));
 OA21x2_ASAP7_75t_R _19033_ (.A1(_08596_),
    .A2(_03276_),
    .B(_03277_),
    .Y(_02214_));
 BUFx16f_ASAP7_75t_R _19034_ (.A(_03275_),
    .Y(_03278_));
 NAND2x1_ASAP7_75t_R _19035_ (.A(_00741_),
    .B(_03278_),
    .Y(_03279_));
 OA21x2_ASAP7_75t_R _19036_ (.A1(_02755_),
    .A2(_03276_),
    .B(_03279_),
    .Y(_02215_));
 NAND2x1_ASAP7_75t_R _19037_ (.A(_00708_),
    .B(_03278_),
    .Y(_03280_));
 OA21x2_ASAP7_75t_R _19038_ (.A1(_02757_),
    .A2(_03276_),
    .B(_03280_),
    .Y(_02216_));
 NAND2x1_ASAP7_75t_R _19039_ (.A(_00675_),
    .B(_03278_),
    .Y(_03281_));
 OA21x2_ASAP7_75t_R _19040_ (.A1(_02759_),
    .A2(_03276_),
    .B(_03281_),
    .Y(_02217_));
 AND2x6_ASAP7_75t_R _19041_ (.A(_08606_),
    .B(_09590_),
    .Y(_03282_));
 BUFx10_ASAP7_75t_R _19042_ (.A(_03282_),
    .Y(_03283_));
 AND2x2_ASAP7_75t_R _19043_ (.A(_00642_),
    .B(_03275_),
    .Y(_03284_));
 AOI21x1_ASAP7_75t_R _19044_ (.A1(_08724_),
    .A2(_03283_),
    .B(_03284_),
    .Y(_02218_));
 NAND2x1_ASAP7_75t_R _19045_ (.A(_00609_),
    .B(_03278_),
    .Y(_03285_));
 OA21x2_ASAP7_75t_R _19046_ (.A1(_02765_),
    .A2(_03276_),
    .B(_03285_),
    .Y(_02219_));
 AO21x1_ASAP7_75t_R _19047_ (.A1(_09208_),
    .A2(_09597_),
    .B(_00575_),
    .Y(_03286_));
 OAI21x1_ASAP7_75t_R _19048_ (.A1(_09769_),
    .A2(_03276_),
    .B(_03286_),
    .Y(_02220_));
 AND3x1_ASAP7_75t_R _19049_ (.A(_02768_),
    .B(_02769_),
    .C(_03283_),
    .Y(_03287_));
 INVx1_ASAP7_75t_R _19050_ (.A(_00542_),
    .Y(_03288_));
 AO32x1_ASAP7_75t_R _19051_ (.A1(_08782_),
    .A2(_08798_),
    .A3(_03287_),
    .B1(_03278_),
    .B2(_03288_),
    .Y(_02221_));
 BUFx4f_ASAP7_75t_R _19052_ (.A(_09547_),
    .Y(_03289_));
 BUFx4f_ASAP7_75t_R _19053_ (.A(_03282_),
    .Y(_03290_));
 AND2x2_ASAP7_75t_R _19054_ (.A(_02773_),
    .B(_03290_),
    .Y(_03291_));
 INVx1_ASAP7_75t_R _19055_ (.A(_00509_),
    .Y(_03292_));
 AO32x1_ASAP7_75t_R _19056_ (.A1(_03289_),
    .A2(_08804_),
    .A3(_03291_),
    .B1(_03278_),
    .B2(_03292_),
    .Y(_02222_));
 AND3x1_ASAP7_75t_R _19057_ (.A(_02776_),
    .B(_02777_),
    .C(_03290_),
    .Y(_03293_));
 BUFx4f_ASAP7_75t_R _19058_ (.A(_03275_),
    .Y(_03294_));
 INVx1_ASAP7_75t_R _19059_ (.A(_00476_),
    .Y(_03295_));
 AO32x1_ASAP7_75t_R _19060_ (.A1(_03289_),
    .A2(_08829_),
    .A3(_03293_),
    .B1(_03294_),
    .B2(_03295_),
    .Y(_02223_));
 AND3x1_ASAP7_75t_R _19061_ (.A(_02780_),
    .B(_02781_),
    .C(_03290_),
    .Y(_03296_));
 INVx1_ASAP7_75t_R _19062_ (.A(_00443_),
    .Y(_03297_));
 AO32x1_ASAP7_75t_R _19063_ (.A1(_03289_),
    .A2(_08849_),
    .A3(_03296_),
    .B1(_03294_),
    .B2(_03297_),
    .Y(_02224_));
 INVx1_ASAP7_75t_R _19064_ (.A(_01040_),
    .Y(_03298_));
 AO21x1_ASAP7_75t_R _19065_ (.A1(_08607_),
    .A2(_09590_),
    .B(_03298_),
    .Y(_03299_));
 OA21x2_ASAP7_75t_R _19066_ (.A1(_02784_),
    .A2(_03276_),
    .B(_03299_),
    .Y(_02225_));
 AND2x2_ASAP7_75t_R _19067_ (.A(_02786_),
    .B(_03290_),
    .Y(_03300_));
 INVx1_ASAP7_75t_R _19068_ (.A(_00410_),
    .Y(_03301_));
 AO32x1_ASAP7_75t_R _19069_ (.A1(_03289_),
    .A2(_08878_),
    .A3(_03300_),
    .B1(_03294_),
    .B2(_03301_),
    .Y(_02226_));
 AND3x1_ASAP7_75t_R _19070_ (.A(_02789_),
    .B(_02790_),
    .C(_03290_),
    .Y(_03302_));
 INVx1_ASAP7_75t_R _19071_ (.A(_00377_),
    .Y(_03303_));
 AO32x1_ASAP7_75t_R _19072_ (.A1(_03289_),
    .A2(_08900_),
    .A3(_03302_),
    .B1(_03294_),
    .B2(_03303_),
    .Y(_02227_));
 AND2x2_ASAP7_75t_R _19073_ (.A(_02793_),
    .B(_03290_),
    .Y(_03304_));
 INVx1_ASAP7_75t_R _19074_ (.A(_00344_),
    .Y(_03305_));
 AO32x1_ASAP7_75t_R _19075_ (.A1(_03289_),
    .A2(_08917_),
    .A3(_03304_),
    .B1(_03294_),
    .B2(_03305_),
    .Y(_02228_));
 AND2x2_ASAP7_75t_R _19076_ (.A(_02796_),
    .B(_03290_),
    .Y(_03306_));
 INVx1_ASAP7_75t_R _19077_ (.A(_00310_),
    .Y(_03307_));
 AO32x1_ASAP7_75t_R _19078_ (.A1(_03289_),
    .A2(_08936_),
    .A3(_03306_),
    .B1(_03294_),
    .B2(_03307_),
    .Y(_02229_));
 AND2x2_ASAP7_75t_R _19079_ (.A(_02799_),
    .B(_03290_),
    .Y(_03308_));
 INVx1_ASAP7_75t_R _19080_ (.A(_00277_),
    .Y(_03309_));
 AO32x1_ASAP7_75t_R _19081_ (.A1(_03289_),
    .A2(_08950_),
    .A3(_03308_),
    .B1(_03294_),
    .B2(_03309_),
    .Y(_02230_));
 AND2x2_ASAP7_75t_R _19082_ (.A(_02802_),
    .B(_03282_),
    .Y(_03310_));
 INVx1_ASAP7_75t_R _19083_ (.A(_00244_),
    .Y(_03311_));
 AO32x1_ASAP7_75t_R _19084_ (.A1(_03289_),
    .A2(_08969_),
    .A3(_03310_),
    .B1(_03294_),
    .B2(_03311_),
    .Y(_02231_));
 NOR2x1_ASAP7_75t_R _19085_ (.A(_08996_),
    .B(_03275_),
    .Y(_03312_));
 INVx1_ASAP7_75t_R _19086_ (.A(_00211_),
    .Y(_03313_));
 AO32x1_ASAP7_75t_R _19087_ (.A1(_03289_),
    .A2(_08986_),
    .A3(_03312_),
    .B1(_03294_),
    .B2(_03313_),
    .Y(_02232_));
 INVx1_ASAP7_75t_R _19088_ (.A(_00177_),
    .Y(_03314_));
 AND2x2_ASAP7_75t_R _19089_ (.A(_02807_),
    .B(_03283_),
    .Y(_03315_));
 AO22x1_ASAP7_75t_R _19090_ (.A1(_03314_),
    .A2(_03278_),
    .B1(_03315_),
    .B2(_09005_),
    .Y(_02233_));
 AND4x1_ASAP7_75t_R _19091_ (.A(_02809_),
    .B(_02810_),
    .C(_02811_),
    .D(_03282_),
    .Y(_03316_));
 INVx1_ASAP7_75t_R _19092_ (.A(_00144_),
    .Y(_03317_));
 AO32x1_ASAP7_75t_R _19093_ (.A1(_08785_),
    .A2(_09024_),
    .A3(_03316_),
    .B1(_03294_),
    .B2(_03317_),
    .Y(_02234_));
 AND3x1_ASAP7_75t_R _19094_ (.A(_02813_),
    .B(_02814_),
    .C(_03290_),
    .Y(_03318_));
 INVx1_ASAP7_75t_R _19095_ (.A(_00110_),
    .Y(_03319_));
 AO32x1_ASAP7_75t_R _19096_ (.A1(_08785_),
    .A2(_09042_),
    .A3(_03318_),
    .B1(_03275_),
    .B2(_03319_),
    .Y(_02235_));
 AO21x1_ASAP7_75t_R _19097_ (.A1(_08607_),
    .A2(_09590_),
    .B(_07032_),
    .Y(_03320_));
 OA21x2_ASAP7_75t_R _19098_ (.A1(_02816_),
    .A2(_03276_),
    .B(_03320_),
    .Y(_02236_));
 AND4x1_ASAP7_75t_R _19099_ (.A(_02818_),
    .B(_02819_),
    .C(_02820_),
    .D(_03282_),
    .Y(_03321_));
 INVx1_ASAP7_75t_R _19100_ (.A(_00076_),
    .Y(_03322_));
 AO32x1_ASAP7_75t_R _19101_ (.A1(_08785_),
    .A2(_09069_),
    .A3(_03321_),
    .B1(_03275_),
    .B2(_03322_),
    .Y(_02237_));
 AND3x1_ASAP7_75t_R _19102_ (.A(_02822_),
    .B(_02823_),
    .C(_03290_),
    .Y(_03323_));
 INVx1_ASAP7_75t_R _19103_ (.A(_00044_),
    .Y(_03324_));
 AO32x1_ASAP7_75t_R _19104_ (.A1(_08785_),
    .A2(_09085_),
    .A3(_03323_),
    .B1(_03275_),
    .B2(_03324_),
    .Y(_02238_));
 NAND2x1_ASAP7_75t_R _19105_ (.A(_00974_),
    .B(_03278_),
    .Y(_03325_));
 OA21x2_ASAP7_75t_R _19106_ (.A1(_02826_),
    .A2(_03276_),
    .B(_03325_),
    .Y(_02239_));
 AO21x1_ASAP7_75t_R _19107_ (.A1(_08607_),
    .A2(_09590_),
    .B(_06854_),
    .Y(_03326_));
 OA21x2_ASAP7_75t_R _19108_ (.A1(_02828_),
    .A2(_03276_),
    .B(_03326_),
    .Y(_02240_));
 AND2x2_ASAP7_75t_R _19109_ (.A(_00907_),
    .B(_03275_),
    .Y(_03327_));
 AOI21x1_ASAP7_75t_R _19110_ (.A1(_09136_),
    .A2(_03283_),
    .B(_03327_),
    .Y(_02241_));
 NOR2x1_ASAP7_75t_R _19111_ (.A(_00874_),
    .B(_03283_),
    .Y(_03328_));
 AO21x1_ASAP7_75t_R _19112_ (.A1(_02831_),
    .A2(_03283_),
    .B(_03328_),
    .Y(_02242_));
 NOR2x1_ASAP7_75t_R _19113_ (.A(_00840_),
    .B(_03283_),
    .Y(_03329_));
 AO21x1_ASAP7_75t_R _19114_ (.A1(_02833_),
    .A2(_03283_),
    .B(_03329_),
    .Y(_02243_));
 NOR2x1_ASAP7_75t_R _19115_ (.A(_00807_),
    .B(_03283_),
    .Y(_03330_));
 AO21x1_ASAP7_75t_R _19116_ (.A1(_02835_),
    .A2(_03283_),
    .B(_03330_),
    .Y(_02244_));
 NAND2x1_ASAP7_75t_R _19117_ (.A(_00773_),
    .B(_03278_),
    .Y(_03331_));
 OA21x2_ASAP7_75t_R _19118_ (.A1(_02837_),
    .A2(_03278_),
    .B(_03331_),
    .Y(_02245_));
 AND2x2_ASAP7_75t_R _19119_ (.A(net64),
    .B(_05852_),
    .Y(_03332_));
 BUFx12f_ASAP7_75t_R _19120_ (.A(_03332_),
    .Y(_03333_));
 NAND2x2_ASAP7_75t_R _19121_ (.A(_05945_),
    .B(_03333_),
    .Y(_03334_));
 AND2x6_ASAP7_75t_R _19122_ (.A(_06284_),
    .B(_03334_),
    .Y(net100));
 AND2x6_ASAP7_75t_R _19123_ (.A(_06186_),
    .B(_03334_),
    .Y(net101));
 AND3x4_ASAP7_75t_R _19124_ (.A(net64),
    .B(_05852_),
    .C(_05945_),
    .Y(_03335_));
 NOR2x2_ASAP7_75t_R _19125_ (.A(_06081_),
    .B(_03335_),
    .Y(net102));
 AND2x6_ASAP7_75t_R _19126_ (.A(_08529_),
    .B(_03334_),
    .Y(net103));
 NOR2x2_ASAP7_75t_R _19127_ (.A(_05900_),
    .B(_03335_),
    .Y(net104));
 NOR2x2_ASAP7_75t_R _19128_ (.A(_05803_),
    .B(_03335_),
    .Y(net105));
 NOR2x2_ASAP7_75t_R _19129_ (.A(_05694_),
    .B(_03333_),
    .Y(net106));
 NAND2x2_ASAP7_75t_R _19130_ (.A(net64),
    .B(_05852_),
    .Y(_03336_));
 AND2x6_ASAP7_75t_R _19131_ (.A(_05596_),
    .B(_03336_),
    .Y(net107));
 AND2x6_ASAP7_75t_R _19132_ (.A(_05494_),
    .B(_03336_),
    .Y(net108));
 AND2x6_ASAP7_75t_R _19133_ (.A(_05396_),
    .B(_03336_),
    .Y(net109));
 AND2x6_ASAP7_75t_R _19134_ (.A(_05300_),
    .B(_03336_),
    .Y(net111));
 AND2x6_ASAP7_75t_R _19135_ (.A(_05209_),
    .B(_03336_),
    .Y(net112));
 NOR2x2_ASAP7_75t_R _19136_ (.A(_05104_),
    .B(_03333_),
    .Y(net113));
 NOR2x2_ASAP7_75t_R _19137_ (.A(_05014_),
    .B(_03333_),
    .Y(net114));
 NOR2x2_ASAP7_75t_R _19138_ (.A(_04895_),
    .B(_03333_),
    .Y(net115));
 NOR2x2_ASAP7_75t_R _19139_ (.A(_04784_),
    .B(_03333_),
    .Y(net116));
 AND2x6_ASAP7_75t_R _19140_ (.A(_04683_),
    .B(_03336_),
    .Y(net117));
 NOR2x2_ASAP7_75t_R _19141_ (.A(_04566_),
    .B(_03333_),
    .Y(net118));
 NOR2x2_ASAP7_75t_R _19142_ (.A(_04431_),
    .B(_03333_),
    .Y(net119));
 NOR2x2_ASAP7_75t_R _19143_ (.A(_04320_),
    .B(_03333_),
    .Y(net120));
 AND2x6_ASAP7_75t_R _19144_ (.A(_04161_),
    .B(_03336_),
    .Y(net122));
 AND2x6_ASAP7_75t_R _19145_ (.A(_04056_),
    .B(_03336_),
    .Y(net123));
 AND2x6_ASAP7_75t_R _19146_ (.A(_06472_),
    .B(_03334_),
    .Y(net129));
 AND2x6_ASAP7_75t_R _19147_ (.A(_06377_),
    .B(_03334_),
    .Y(net130));
 AND2x2_ASAP7_75t_R _19148_ (.A(net64),
    .B(\dmem.ce_mem[0] ),
    .Y(\dmem.we_mem[0] ));
 AND2x2_ASAP7_75t_R _19149_ (.A(net64),
    .B(\dmem.ce_mem[1] ),
    .Y(\dmem.we_mem[1] ));
 AND3x1_ASAP7_75t_R _19150_ (.A(net64),
    .B(net47),
    .C(_08658_),
    .Y(\dmem.we_mem[2] ));
 AND2x2_ASAP7_75t_R _19151_ (.A(net64),
    .B(\dmem.ce_mem[3] ),
    .Y(\dmem.we_mem[3] ));
 AND3x1_ASAP7_75t_R _19152_ (.A(_08550_),
    .B(_08571_),
    .C(_08652_),
    .Y(_03337_));
 AO21x1_ASAP7_75t_R _19153_ (.A1(_08572_),
    .A2(_08646_),
    .B(_03337_),
    .Y(\riscv.dp.ISRmux.d0[10] ));
 AO21x1_ASAP7_75t_R _19154_ (.A1(_08574_),
    .A2(_08575_),
    .B(_08673_),
    .Y(_03338_));
 OA21x2_ASAP7_75t_R _19155_ (.A1(_08573_),
    .A2(_08678_),
    .B(_03338_),
    .Y(\riscv.dp.ISRmux.d0[11] ));
 AND2x6_ASAP7_75t_R _19156_ (.A(_08550_),
    .B(_08571_),
    .Y(_03339_));
 BUFx4f_ASAP7_75t_R _19157_ (.A(_03339_),
    .Y(_03340_));
 NOR2x1_ASAP7_75t_R _19158_ (.A(_03339_),
    .B(_08691_),
    .Y(_03341_));
 AO21x1_ASAP7_75t_R _19159_ (.A1(_03340_),
    .A2(_08693_),
    .B(_03341_),
    .Y(\riscv.dp.ISRmux.d0[12] ));
 BUFx6f_ASAP7_75t_R _19160_ (.A(_08572_),
    .Y(_03342_));
 BUFx4f_ASAP7_75t_R _19161_ (.A(_08550_),
    .Y(_03343_));
 BUFx4f_ASAP7_75t_R _19162_ (.A(_08571_),
    .Y(_03344_));
 AND3x1_ASAP7_75t_R _19163_ (.A(_03343_),
    .B(_03344_),
    .C(_08717_),
    .Y(_03345_));
 AOI21x1_ASAP7_75t_R _19164_ (.A1(_03342_),
    .A2(_08721_),
    .B(_03345_),
    .Y(\riscv.dp.ISRmux.d0[13] ));
 NOR2x1_ASAP7_75t_R _19165_ (.A(_03339_),
    .B(_08740_),
    .Y(_03346_));
 AO21x1_ASAP7_75t_R _19166_ (.A1(_03340_),
    .A2(_08734_),
    .B(_03346_),
    .Y(\riscv.dp.ISRmux.d0[14] ));
 NAND2x1_ASAP7_75t_R _19167_ (.A(_03340_),
    .B(_08757_),
    .Y(_03347_));
 OA21x2_ASAP7_75t_R _19168_ (.A1(_03340_),
    .A2(_08762_),
    .B(_03347_),
    .Y(\riscv.dp.ISRmux.d0[15] ));
 AND3x1_ASAP7_75t_R _19169_ (.A(_03343_),
    .B(_03344_),
    .C(_08788_),
    .Y(_03348_));
 AOI21x1_ASAP7_75t_R _19170_ (.A1(_03342_),
    .A2(_08793_),
    .B(_03348_),
    .Y(\riscv.dp.ISRmux.d0[16] ));
 AO21x1_ASAP7_75t_R _19171_ (.A1(_08574_),
    .A2(_08575_),
    .B(_08818_),
    .Y(_03349_));
 OAI21x1_ASAP7_75t_R _19172_ (.A1(_03342_),
    .A2(_08811_),
    .B(_03349_),
    .Y(\riscv.dp.ISRmux.d0[17] ));
 AND3x1_ASAP7_75t_R _19173_ (.A(_03343_),
    .B(_03344_),
    .C(_08836_),
    .Y(_03350_));
 AOI21x1_ASAP7_75t_R _19174_ (.A1(_03342_),
    .A2(_08840_),
    .B(_03350_),
    .Y(\riscv.dp.ISRmux.d0[18] ));
 AND3x1_ASAP7_75t_R _19175_ (.A(_03343_),
    .B(_03344_),
    .C(_08854_),
    .Y(_03351_));
 AOI21x1_ASAP7_75t_R _19176_ (.A1(_03342_),
    .A2(_08859_),
    .B(_03351_),
    .Y(\riscv.dp.ISRmux.d0[19] ));
 AO21x1_ASAP7_75t_R _19177_ (.A1(_08574_),
    .A2(_08575_),
    .B(_08888_),
    .Y(_03352_));
 OA21x2_ASAP7_75t_R _19178_ (.A1(_08573_),
    .A2(_08890_),
    .B(_03352_),
    .Y(\riscv.dp.ISRmux.d0[20] ));
 AND3x1_ASAP7_75t_R _19179_ (.A(_03343_),
    .B(_03344_),
    .C(_08905_),
    .Y(_03353_));
 AOI21x1_ASAP7_75t_R _19180_ (.A1(_03342_),
    .A2(_08909_),
    .B(_03353_),
    .Y(\riscv.dp.ISRmux.d0[21] ));
 AO21x1_ASAP7_75t_R _19181_ (.A1(_08574_),
    .A2(_08575_),
    .B(_08924_),
    .Y(_03354_));
 OAI21x1_ASAP7_75t_R _19182_ (.A1(_03342_),
    .A2(_08927_),
    .B(_03354_),
    .Y(\riscv.dp.ISRmux.d0[22] ));
 OR2x2_ASAP7_75t_R _19183_ (.A(_08572_),
    .B(_08942_),
    .Y(_03355_));
 OA21x2_ASAP7_75t_R _19184_ (.A1(_03340_),
    .A2(_08940_),
    .B(_03355_),
    .Y(\riscv.dp.ISRmux.d0[23] ));
 AND3x1_ASAP7_75t_R _19185_ (.A(_03343_),
    .B(_03344_),
    .C(_08960_),
    .Y(_03356_));
 AOI21x1_ASAP7_75t_R _19186_ (.A1(_08573_),
    .A2(_08957_),
    .B(_03356_),
    .Y(\riscv.dp.ISRmux.d0[24] ));
 NOR2x1_ASAP7_75t_R _19187_ (.A(_03339_),
    .B(_08974_),
    .Y(_03357_));
 AO21x1_ASAP7_75t_R _19188_ (.A1(_03340_),
    .A2(_08976_),
    .B(_03357_),
    .Y(\riscv.dp.ISRmux.d0[25] ));
 AO21x1_ASAP7_75t_R _19189_ (.A1(_08574_),
    .A2(_08575_),
    .B(_08992_),
    .Y(_03358_));
 OAI21x1_ASAP7_75t_R _19190_ (.A1(_03342_),
    .A2(_08995_),
    .B(_03358_),
    .Y(\riscv.dp.ISRmux.d0[26] ));
 AND3x1_ASAP7_75t_R _19191_ (.A(_03343_),
    .B(_03344_),
    .C(_09009_),
    .Y(_03359_));
 AOI21x1_ASAP7_75t_R _19192_ (.A1(_08573_),
    .A2(_09015_),
    .B(_03359_),
    .Y(\riscv.dp.ISRmux.d0[27] ));
 NOR2x1_ASAP7_75t_R _19193_ (.A(_03339_),
    .B(_09029_),
    .Y(_03360_));
 AO21x1_ASAP7_75t_R _19194_ (.A1(_03340_),
    .A2(_09034_),
    .B(_03360_),
    .Y(\riscv.dp.ISRmux.d0[28] ));
 NOR2x1_ASAP7_75t_R _19195_ (.A(_03339_),
    .B(_09047_),
    .Y(_03361_));
 AO21x1_ASAP7_75t_R _19196_ (.A1(_03340_),
    .A2(_09050_),
    .B(_03361_),
    .Y(\riscv.dp.ISRmux.d0[29] ));
 AO21x1_ASAP7_75t_R _19197_ (.A1(_08574_),
    .A2(_08575_),
    .B(_09054_),
    .Y(_03362_));
 OA21x2_ASAP7_75t_R _19198_ (.A1(_10109_),
    .A2(_08572_),
    .B(_03362_),
    .Y(\riscv.dp.ISRmux.d0[2] ));
 NAND2x1_ASAP7_75t_R _19199_ (.A(_08572_),
    .B(_09073_),
    .Y(_03363_));
 OA21x2_ASAP7_75t_R _19200_ (.A1(_08573_),
    .A2(_09076_),
    .B(_03363_),
    .Y(\riscv.dp.ISRmux.d0[30] ));
 NAND2x1_ASAP7_75t_R _19201_ (.A(_03339_),
    .B(_09096_),
    .Y(_03364_));
 OA21x2_ASAP7_75t_R _19202_ (.A1(_03340_),
    .A2(_09093_),
    .B(_03364_),
    .Y(\riscv.dp.ISRmux.d0[31] ));
 AO21x1_ASAP7_75t_R _19203_ (.A1(_03343_),
    .A2(_03344_),
    .B(_09104_),
    .Y(_03365_));
 OA21x2_ASAP7_75t_R _19204_ (.A1(_09105_),
    .A2(_08572_),
    .B(_03365_),
    .Y(\riscv.dp.ISRmux.d0[3] ));
 AO21x1_ASAP7_75t_R _19205_ (.A1(_03343_),
    .A2(_03344_),
    .B(_09117_),
    .Y(_03366_));
 OA21x2_ASAP7_75t_R _19206_ (.A1(_08573_),
    .A2(_09118_),
    .B(_03366_),
    .Y(\riscv.dp.ISRmux.d0[4] ));
 NOR2x1_ASAP7_75t_R _19207_ (.A(_03339_),
    .B(_09126_),
    .Y(_03367_));
 AO21x1_ASAP7_75t_R _19208_ (.A1(_03340_),
    .A2(_09133_),
    .B(_03367_),
    .Y(\riscv.dp.ISRmux.d0[5] ));
 AO21x1_ASAP7_75t_R _19209_ (.A1(_08574_),
    .A2(_08575_),
    .B(_09145_),
    .Y(_03368_));
 OAI21x1_ASAP7_75t_R _19210_ (.A1(_03342_),
    .A2(_09146_),
    .B(_03368_),
    .Y(\riscv.dp.ISRmux.d0[6] ));
 AND3x1_ASAP7_75t_R _19211_ (.A(_08550_),
    .B(_08571_),
    .C(_09154_),
    .Y(_03369_));
 AOI21x1_ASAP7_75t_R _19212_ (.A1(_08573_),
    .A2(_09152_),
    .B(_03369_),
    .Y(\riscv.dp.ISRmux.d0[7] ));
 AO21x1_ASAP7_75t_R _19213_ (.A1(_03343_),
    .A2(_03344_),
    .B(_09169_),
    .Y(_03370_));
 OA21x2_ASAP7_75t_R _19214_ (.A1(_08573_),
    .A2(_09171_),
    .B(_03370_),
    .Y(\riscv.dp.ISRmux.d0[8] ));
 AO21x1_ASAP7_75t_R _19215_ (.A1(_08574_),
    .A2(_08575_),
    .B(_09179_),
    .Y(_03371_));
 OAI21x1_ASAP7_75t_R _19216_ (.A1(_03342_),
    .A2(_09176_),
    .B(_03371_),
    .Y(\riscv.dp.ISRmux.d0[9] ));
 AND4x2_ASAP7_75t_R _19217_ (.A(net89),
    .B(net27),
    .C(_03501_),
    .D(_08568_),
    .Y(net98));
 FAx1_ASAP7_75t_R _19218_ (.SN(_01066_),
    .A(_09940_),
    .B(_09941_),
    .CI(_09942_),
    .CON(_01064_));
 FAx1_ASAP7_75t_R _19219_ (.SN(_01072_),
    .A(_09943_),
    .B(_09944_),
    .CI(_09945_),
    .CON(_01160_));
 HAxp5_ASAP7_75t_R _19220_ (.A(_09947_),
    .B(_09948_),
    .CON(_01065_),
    .SN(_00034_));
 HAxp5_ASAP7_75t_R _19221_ (.A(_09949_),
    .B(_09950_),
    .CON(_01161_),
    .SN(_09951_));
 HAxp5_ASAP7_75t_R _19222_ (.A(_09952_),
    .B(_09953_),
    .CON(_01162_),
    .SN(_01163_));
 HAxp5_ASAP7_75t_R _19223_ (.A(_09954_),
    .B(_09955_),
    .CON(_01164_),
    .SN(_09956_));
 HAxp5_ASAP7_75t_R _19224_ (.A(_09957_),
    .B(_09958_),
    .CON(_01165_),
    .SN(_00100_));
 HAxp5_ASAP7_75t_R _19225_ (.A(_09959_),
    .B(_09960_),
    .CON(_00099_),
    .SN(_09961_));
 HAxp5_ASAP7_75t_R _19226_ (.A(_09962_),
    .B(_09963_),
    .CON(_01166_),
    .SN(_00134_));
 HAxp5_ASAP7_75t_R _19227_ (.A(_09964_),
    .B(_09965_),
    .CON(_00133_),
    .SN(_09966_));
 HAxp5_ASAP7_75t_R _19228_ (.A(_09967_),
    .B(_09968_),
    .CON(_01167_),
    .SN(_00167_));
 HAxp5_ASAP7_75t_R _19229_ (.A(_09969_),
    .B(_09970_),
    .CON(_01168_),
    .SN(_09971_));
 HAxp5_ASAP7_75t_R _19230_ (.A(_09972_),
    .B(_09973_),
    .CON(_01169_),
    .SN(_00201_));
 HAxp5_ASAP7_75t_R _19231_ (.A(_09974_),
    .B(_09975_),
    .CON(_00200_),
    .SN(_09976_));
 HAxp5_ASAP7_75t_R _19232_ (.A(_09977_),
    .B(_09978_),
    .CON(_01170_),
    .SN(_00234_));
 HAxp5_ASAP7_75t_R _19233_ (.A(_09979_),
    .B(_09980_),
    .CON(_01171_),
    .SN(_09981_));
 HAxp5_ASAP7_75t_R _19234_ (.A(_09982_),
    .B(_09983_),
    .CON(_01172_),
    .SN(_00267_));
 HAxp5_ASAP7_75t_R _19235_ (.A(_09984_),
    .B(_09985_),
    .CON(_01173_),
    .SN(_09986_));
 HAxp5_ASAP7_75t_R _19236_ (.A(_09987_),
    .B(_09988_),
    .CON(_01174_),
    .SN(_00300_));
 HAxp5_ASAP7_75t_R _19237_ (.A(_09989_),
    .B(_09990_),
    .CON(_01175_),
    .SN(_09991_));
 HAxp5_ASAP7_75t_R _19238_ (.A(_09992_),
    .B(_09993_),
    .CON(_00333_),
    .SN(_00334_));
 HAxp5_ASAP7_75t_R _19239_ (.A(_09994_),
    .B(_09995_),
    .CON(_01176_),
    .SN(_09996_));
 HAxp5_ASAP7_75t_R _19240_ (.A(_09997_),
    .B(_09998_),
    .CON(_01177_),
    .SN(_00367_));
 HAxp5_ASAP7_75t_R _19241_ (.A(_09999_),
    .B(_10000_),
    .CON(_01178_),
    .SN(_10001_));
 HAxp5_ASAP7_75t_R _19242_ (.A(_10002_),
    .B(_10003_),
    .CON(_01179_),
    .SN(_00400_));
 HAxp5_ASAP7_75t_R _19243_ (.A(_10004_),
    .B(_10005_),
    .CON(_01180_),
    .SN(_10006_));
 HAxp5_ASAP7_75t_R _19244_ (.A(_10007_),
    .B(_10008_),
    .CON(_01181_),
    .SN(_00433_));
 HAxp5_ASAP7_75t_R _19245_ (.A(_10009_),
    .B(_10010_),
    .CON(_01182_),
    .SN(_10011_));
 HAxp5_ASAP7_75t_R _19246_ (.A(_10012_),
    .B(_10013_),
    .CON(_01183_),
    .SN(_00466_));
 HAxp5_ASAP7_75t_R _19247_ (.A(_10014_),
    .B(_10015_),
    .CON(_01184_),
    .SN(_10016_));
 HAxp5_ASAP7_75t_R _19248_ (.A(_10017_),
    .B(_10018_),
    .CON(_01185_),
    .SN(_00499_));
 HAxp5_ASAP7_75t_R _19249_ (.A(_10019_),
    .B(_10020_),
    .CON(_01186_),
    .SN(_10021_));
 HAxp5_ASAP7_75t_R _19250_ (.A(_10022_),
    .B(_10023_),
    .CON(_01187_),
    .SN(_00532_));
 HAxp5_ASAP7_75t_R _19251_ (.A(_10024_),
    .B(_10025_),
    .CON(_01188_),
    .SN(_10026_));
 HAxp5_ASAP7_75t_R _19252_ (.A(_10027_),
    .B(_10028_),
    .CON(_01189_),
    .SN(_00565_));
 HAxp5_ASAP7_75t_R _19253_ (.A(_10029_),
    .B(_10030_),
    .CON(_01190_),
    .SN(_10031_));
 HAxp5_ASAP7_75t_R _19254_ (.A(_10032_),
    .B(_10033_),
    .CON(_00598_),
    .SN(_00599_));
 HAxp5_ASAP7_75t_R _19255_ (.A(_10034_),
    .B(_10035_),
    .CON(_01191_),
    .SN(_10036_));
 HAxp5_ASAP7_75t_R _19256_ (.A(_10037_),
    .B(_10038_),
    .CON(_01192_),
    .SN(_00632_));
 HAxp5_ASAP7_75t_R _19257_ (.A(_10039_),
    .B(_10040_),
    .CON(_01193_),
    .SN(_10041_));
 HAxp5_ASAP7_75t_R _19258_ (.A(_10042_),
    .B(_10043_),
    .CON(_01194_),
    .SN(_00665_));
 HAxp5_ASAP7_75t_R _19259_ (.A(_10044_),
    .B(_10045_),
    .CON(_01195_),
    .SN(_10046_));
 HAxp5_ASAP7_75t_R _19260_ (.A(_10047_),
    .B(_10048_),
    .CON(_01196_),
    .SN(_00698_));
 HAxp5_ASAP7_75t_R _19261_ (.A(_10049_),
    .B(_10050_),
    .CON(_01197_),
    .SN(_10051_));
 HAxp5_ASAP7_75t_R _19262_ (.A(_10052_),
    .B(_10053_),
    .CON(_01198_),
    .SN(_00731_));
 HAxp5_ASAP7_75t_R _19263_ (.A(_10054_),
    .B(_10055_),
    .CON(_01199_),
    .SN(_10056_));
 HAxp5_ASAP7_75t_R _19264_ (.A(_10057_),
    .B(_10058_),
    .CON(_00796_),
    .SN(_00797_));
 HAxp5_ASAP7_75t_R _19265_ (.A(_10059_),
    .B(_10060_),
    .CON(_01200_),
    .SN(_10061_));
 HAxp5_ASAP7_75t_R _19266_ (.A(_10062_),
    .B(_10063_),
    .CON(_01201_),
    .SN(_00830_));
 HAxp5_ASAP7_75t_R _19267_ (.A(_10064_),
    .B(_10065_),
    .CON(_01202_),
    .SN(_10066_));
 HAxp5_ASAP7_75t_R _19268_ (.A(_10067_),
    .B(_10068_),
    .CON(_00863_),
    .SN(_00864_));
 HAxp5_ASAP7_75t_R _19269_ (.A(_10069_),
    .B(_10070_),
    .CON(_01203_),
    .SN(_10071_));
 HAxp5_ASAP7_75t_R _19270_ (.A(_10072_),
    .B(_10073_),
    .CON(_01204_),
    .SN(_00897_));
 HAxp5_ASAP7_75t_R _19271_ (.A(_10074_),
    .B(_10075_),
    .CON(_01205_),
    .SN(_10076_));
 HAxp5_ASAP7_75t_R _19272_ (.A(_10077_),
    .B(_10078_),
    .CON(_00930_),
    .SN(_00931_));
 HAxp5_ASAP7_75t_R _19273_ (.A(_10079_),
    .B(_10080_),
    .CON(_01206_),
    .SN(_10081_));
 HAxp5_ASAP7_75t_R _19274_ (.A(_10082_),
    .B(_10083_),
    .CON(_01207_),
    .SN(_00964_));
 HAxp5_ASAP7_75t_R _19275_ (.A(_10084_),
    .B(_10085_),
    .CON(_01208_),
    .SN(_10086_));
 HAxp5_ASAP7_75t_R _19276_ (.A(_10087_),
    .B(_10088_),
    .CON(_01209_),
    .SN(_00997_));
 HAxp5_ASAP7_75t_R _19277_ (.A(_10089_),
    .B(_10090_),
    .CON(_01210_),
    .SN(_10091_));
 HAxp5_ASAP7_75t_R _19278_ (.A(_10092_),
    .B(_10093_),
    .CON(_01211_),
    .SN(_01030_));
 HAxp5_ASAP7_75t_R _19279_ (.A(_10094_),
    .B(_10095_),
    .CON(_01212_),
    .SN(_10096_));
 HAxp5_ASAP7_75t_R _19280_ (.A(_09941_),
    .B(_09942_),
    .CON(_01213_),
    .SN(_01063_));
 HAxp5_ASAP7_75t_R _19281_ (.A(_10097_),
    .B(_10098_),
    .CON(_01214_),
    .SN(_10099_));
 HAxp5_ASAP7_75t_R _19282_ (.A(_10100_),
    .B(_10101_),
    .CON(_01215_),
    .SN(_01067_));
 HAxp5_ASAP7_75t_R _19283_ (.A(_10102_),
    .B(_10103_),
    .CON(_01216_),
    .SN(_10104_));
 HAxp5_ASAP7_75t_R _19284_ (.A(_10105_),
    .B(_10106_),
    .CON(_09946_),
    .SN(_01069_));
 HAxp5_ASAP7_75t_R _19285_ (.A(_09944_),
    .B(_09945_),
    .CON(_01074_),
    .SN(_01071_));
 HAxp5_ASAP7_75t_R _19286_ (.A(_10107_),
    .B(_10108_),
    .CON(_01076_),
    .SN(_01073_));
 HAxp5_ASAP7_75t_R _19287_ (.A(_10109_),
    .B(_10110_),
    .CON(_00032_),
    .SN(_01217_));
 HAxp5_ASAP7_75t_R _19288_ (.A(net87),
    .B(_10110_),
    .CON(_00033_),
    .SN(_10111_));
 HAxp5_ASAP7_75t_R _19289_ (.A(net87),
    .B(net90),
    .CON(_01218_),
    .SN(_10112_));
 HAxp5_ASAP7_75t_R _19290_ (.A(_10113_),
    .B(_10114_),
    .CON(_01079_),
    .SN(_01075_));
 HAxp5_ASAP7_75t_R _19291_ (.A(_10115_),
    .B(_10116_),
    .CON(_01082_),
    .SN(_01078_));
 HAxp5_ASAP7_75t_R _19292_ (.A(_10117_),
    .B(_10118_),
    .CON(_01085_),
    .SN(_01081_));
 HAxp5_ASAP7_75t_R _19293_ (.A(_10119_),
    .B(_10120_),
    .CON(_01088_),
    .SN(_01084_));
 HAxp5_ASAP7_75t_R _19294_ (.A(_10121_),
    .B(_10122_),
    .CON(_01091_),
    .SN(_01087_));
 HAxp5_ASAP7_75t_R _19295_ (.A(_10123_),
    .B(_10124_),
    .CON(_01094_),
    .SN(_01090_));
 HAxp5_ASAP7_75t_R _19296_ (.A(_10125_),
    .B(_10126_),
    .CON(_01097_),
    .SN(_01093_));
 HAxp5_ASAP7_75t_R _19297_ (.A(_10127_),
    .B(_10128_),
    .CON(_01100_),
    .SN(_01096_));
 HAxp5_ASAP7_75t_R _19298_ (.A(_10129_),
    .B(_10130_),
    .CON(_01103_),
    .SN(_01099_));
 HAxp5_ASAP7_75t_R _19299_ (.A(_10131_),
    .B(_10132_),
    .CON(_01106_),
    .SN(_01102_));
 HAxp5_ASAP7_75t_R _19300_ (.A(_10133_),
    .B(_10134_),
    .CON(_01109_),
    .SN(_01105_));
 HAxp5_ASAP7_75t_R _19301_ (.A(_10135_),
    .B(_10136_),
    .CON(_01112_),
    .SN(_01108_));
 HAxp5_ASAP7_75t_R _19302_ (.A(_10137_),
    .B(_10138_),
    .CON(_01115_),
    .SN(_01111_));
 HAxp5_ASAP7_75t_R _19303_ (.A(_10139_),
    .B(_10140_),
    .CON(_01118_),
    .SN(_01114_));
 HAxp5_ASAP7_75t_R _19304_ (.A(_10141_),
    .B(_10142_),
    .CON(_01121_),
    .SN(_01117_));
 HAxp5_ASAP7_75t_R _19305_ (.A(_10143_),
    .B(_10144_),
    .CON(_01124_),
    .SN(_01120_));
 HAxp5_ASAP7_75t_R _19306_ (.A(_10145_),
    .B(_10146_),
    .CON(_01127_),
    .SN(_01123_));
 HAxp5_ASAP7_75t_R _19307_ (.A(_10147_),
    .B(_10148_),
    .CON(_01130_),
    .SN(_01126_));
 HAxp5_ASAP7_75t_R _19308_ (.A(_10149_),
    .B(_10150_),
    .CON(_01133_),
    .SN(_01129_));
 HAxp5_ASAP7_75t_R _19309_ (.A(_10151_),
    .B(_10152_),
    .CON(_01136_),
    .SN(_01132_));
 HAxp5_ASAP7_75t_R _19310_ (.A(_10153_),
    .B(_10154_),
    .CON(_01139_),
    .SN(_01135_));
 HAxp5_ASAP7_75t_R _19311_ (.A(_10155_),
    .B(_10156_),
    .CON(_01142_),
    .SN(_01138_));
 HAxp5_ASAP7_75t_R _19312_ (.A(_10157_),
    .B(_10158_),
    .CON(_01145_),
    .SN(_01141_));
 HAxp5_ASAP7_75t_R _19313_ (.A(_10159_),
    .B(_10160_),
    .CON(_01148_),
    .SN(_01144_));
 HAxp5_ASAP7_75t_R _19314_ (.A(_10161_),
    .B(_10162_),
    .CON(_01151_),
    .SN(_01147_));
 HAxp5_ASAP7_75t_R _19315_ (.A(_10163_),
    .B(_10164_),
    .CON(_01154_),
    .SN(_01150_));
 HAxp5_ASAP7_75t_R _19316_ (.A(_10165_),
    .B(_10166_),
    .CON(_01157_),
    .SN(_01153_));
 HAxp5_ASAP7_75t_R _19317_ (.A(_10167_),
    .B(_10168_),
    .CON(_01158_),
    .SN(_01156_));
 BUFx16f_ASAP7_75t_R clkbuf_regs_0_clk (.A(clk),
    .Y(clk_regs));
 BUFx3_ASAP7_75t_R _19319_ (.A(\dmem.ce_mem[3] ),
    .Y(net56));
 BUFx2_ASAP7_75t_R _19320_ (.A(valid),
    .Y(net97));
 fakeram7_256x32 \dmem.dmem0  (.ce_in(\dmem.ce_mem[0] ),
    .clk(clknet_1_1__leaf_clk),
    .we_in(\dmem.we_mem[0] ),
    .addr_in({net61,
    net60,
    net59,
    net58,
    net57,
    net54,
    net43,
    net32}),
    .rd_out({\dmem.inter_dmem0[31] ,
    \dmem.inter_dmem0[30] ,
    \dmem.inter_dmem0[29] ,
    \dmem.inter_dmem0[28] ,
    \dmem.inter_dmem0[27] ,
    \dmem.inter_dmem0[26] ,
    \dmem.inter_dmem0[25] ,
    \dmem.inter_dmem0[24] ,
    \dmem.inter_dmem0[23] ,
    \dmem.inter_dmem0[22] ,
    \dmem.inter_dmem0[21] ,
    \dmem.inter_dmem0[20] ,
    \dmem.inter_dmem0[19] ,
    \dmem.inter_dmem0[18] ,
    \dmem.inter_dmem0[17] ,
    \dmem.inter_dmem0[16] ,
    \dmem.inter_dmem0[15] ,
    \dmem.inter_dmem0[14] ,
    \dmem.inter_dmem0[13] ,
    \dmem.inter_dmem0[12] ,
    \dmem.inter_dmem0[11] ,
    \dmem.inter_dmem0[10] ,
    \dmem.inter_dmem0[9] ,
    \dmem.inter_dmem0[8] ,
    \dmem.inter_dmem0[7] ,
    \dmem.inter_dmem0[6] ,
    \dmem.inter_dmem0[5] ,
    \dmem.inter_dmem0[4] ,
    \dmem.inter_dmem0[3] ,
    \dmem.inter_dmem0[2] ,
    \dmem.inter_dmem0[1] ,
    \dmem.inter_dmem0[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net126,
    net125,
    net124,
    net121,
    net110,
    net99}));
 fakeram7_256x32 \dmem.dmem1  (.ce_in(\dmem.ce_mem[1] ),
    .clk(clknet_1_0__leaf_clk),
    .we_in(\dmem.we_mem[1] ),
    .addr_in({net38,
    net37,
    net36,
    net35,
    net34,
    net33,
    net63,
    net62}),
    .rd_out({\dmem.inter_dmem1[31] ,
    \dmem.inter_dmem1[30] ,
    \dmem.inter_dmem1[29] ,
    \dmem.inter_dmem1[28] ,
    \dmem.inter_dmem1[27] ,
    \dmem.inter_dmem1[26] ,
    \dmem.inter_dmem1[25] ,
    \dmem.inter_dmem1[24] ,
    \dmem.inter_dmem1[23] ,
    \dmem.inter_dmem1[22] ,
    \dmem.inter_dmem1[21] ,
    \dmem.inter_dmem1[20] ,
    \dmem.inter_dmem1[19] ,
    \dmem.inter_dmem1[18] ,
    \dmem.inter_dmem1[17] ,
    \dmem.inter_dmem1[16] ,
    \dmem.inter_dmem1[15] ,
    \dmem.inter_dmem1[14] ,
    \dmem.inter_dmem1[13] ,
    \dmem.inter_dmem1[12] ,
    \dmem.inter_dmem1[11] ,
    \dmem.inter_dmem1[10] ,
    \dmem.inter_dmem1[9] ,
    \dmem.inter_dmem1[8] ,
    \dmem.inter_dmem1[7] ,
    \dmem.inter_dmem1[6] ,
    \dmem.inter_dmem1[5] ,
    \dmem.inter_dmem1[4] ,
    \dmem.inter_dmem1[3] ,
    \dmem.inter_dmem1[2] ,
    \dmem.inter_dmem1[1] ,
    \dmem.inter_dmem1[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net126,
    net125,
    net124,
    net121,
    net110,
    net99}));
 fakeram7_256x32 \dmem.dmem2  (.ce_in(\dmem.ce_mem[2] ),
    .clk(clknet_1_0__leaf_clk),
    .we_in(\dmem.we_mem[2] ),
    .addr_in({net47,
    net46,
    net45,
    net44,
    net42,
    net41,
    net40,
    net39}),
    .rd_out({\dmem.inter_dmem2[31] ,
    \dmem.inter_dmem2[30] ,
    \dmem.inter_dmem2[29] ,
    \dmem.inter_dmem2[28] ,
    \dmem.inter_dmem2[27] ,
    \dmem.inter_dmem2[26] ,
    \dmem.inter_dmem2[25] ,
    \dmem.inter_dmem2[24] ,
    \dmem.inter_dmem2[23] ,
    \dmem.inter_dmem2[22] ,
    \dmem.inter_dmem2[21] ,
    \dmem.inter_dmem2[20] ,
    \dmem.inter_dmem2[19] ,
    \dmem.inter_dmem2[18] ,
    \dmem.inter_dmem2[17] ,
    \dmem.inter_dmem2[16] ,
    \dmem.inter_dmem2[15] ,
    \dmem.inter_dmem2[14] ,
    \dmem.inter_dmem2[13] ,
    \dmem.inter_dmem2[12] ,
    \dmem.inter_dmem2[11] ,
    \dmem.inter_dmem2[10] ,
    \dmem.inter_dmem2[9] ,
    \dmem.inter_dmem2[8] ,
    \dmem.inter_dmem2[7] ,
    \dmem.inter_dmem2[6] ,
    \dmem.inter_dmem2[5] ,
    \dmem.inter_dmem2[4] ,
    \dmem.inter_dmem2[3] ,
    \dmem.inter_dmem2[2] ,
    \dmem.inter_dmem2[1] ,
    \dmem.inter_dmem2[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net126,
    net125,
    net124,
    net121,
    net110,
    net99}));
 fakeram7_256x32 \dmem.dmem3  (.ce_in(\dmem.ce_mem[3] ),
    .clk(clknet_1_1__leaf_clk),
    .we_in(\dmem.we_mem[3] ),
    .addr_in({\dmem.ce_mem[3] ,
    net55,
    net53,
    net52,
    net51,
    net50,
    net49,
    net48}),
    .rd_out({\dmem.inter_dmem3[31] ,
    \dmem.inter_dmem3[30] ,
    \dmem.inter_dmem3[29] ,
    \dmem.inter_dmem3[28] ,
    \dmem.inter_dmem3[27] ,
    \dmem.inter_dmem3[26] ,
    \dmem.inter_dmem3[25] ,
    \dmem.inter_dmem3[24] ,
    \dmem.inter_dmem3[23] ,
    \dmem.inter_dmem3[22] ,
    \dmem.inter_dmem3[21] ,
    \dmem.inter_dmem3[20] ,
    \dmem.inter_dmem3[19] ,
    \dmem.inter_dmem3[18] ,
    \dmem.inter_dmem3[17] ,
    \dmem.inter_dmem3[16] ,
    \dmem.inter_dmem3[15] ,
    \dmem.inter_dmem3[14] ,
    \dmem.inter_dmem3[13] ,
    \dmem.inter_dmem3[12] ,
    \dmem.inter_dmem3[11] ,
    \dmem.inter_dmem3[10] ,
    \dmem.inter_dmem3[9] ,
    \dmem.inter_dmem3[8] ,
    \dmem.inter_dmem3[7] ,
    \dmem.inter_dmem3[6] ,
    \dmem.inter_dmem3[5] ,
    \dmem.inter_dmem3[4] ,
    \dmem.inter_dmem3[3] ,
    \dmem.inter_dmem3[2] ,
    \dmem.inter_dmem3[1] ,
    \dmem.inter_dmem3[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net126,
    net125,
    net124,
    net121,
    net110,
    net99}));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk_regs),
    .D(_01220_),
    .QN(_01068_),
    .RESETN(net131),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[10]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[10] ),
    .QN(_01095_),
    .RESETN(net132),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[11]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[11] ),
    .QN(_01098_),
    .RESETN(net133),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[12]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[12] ),
    .QN(_01101_),
    .RESETN(net134),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[13]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[13] ),
    .QN(_01104_),
    .RESETN(net135),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[14]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[14] ),
    .QN(_01107_),
    .RESETN(net136),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[15]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[15] ),
    .QN(_01110_),
    .RESETN(net137),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[16]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[16] ),
    .QN(_01113_),
    .RESETN(net138),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[17]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[17] ),
    .QN(_01116_),
    .RESETN(net139),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[18]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[18] ),
    .QN(_01119_),
    .RESETN(net140),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[19]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[19] ),
    .QN(_01122_),
    .RESETN(net141),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_2_clk_regs),
    .D(_01221_),
    .QN(_01070_),
    .RESETN(net142),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[20]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[20] ),
    .QN(_01125_),
    .RESETN(net143),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[21]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[21] ),
    .QN(_01128_),
    .RESETN(net144),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[22]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[22] ),
    .QN(_01131_),
    .RESETN(net145),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[23]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[23] ),
    .QN(_01134_),
    .RESETN(net146),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[24]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[24] ),
    .QN(_01137_),
    .RESETN(net147),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[25]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[25] ),
    .QN(_01140_),
    .RESETN(net148),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[26]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[26] ),
    .QN(_01143_),
    .RESETN(net149),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[27]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[27] ),
    .QN(_01146_),
    .RESETN(net150),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[28]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[28] ),
    .QN(_01149_),
    .RESETN(net151),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[29]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[29] ),
    .QN(_01152_),
    .RESETN(net152),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[2]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[2] ),
    .QN(_10109_),
    .RESETN(net153),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[30]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[30] ),
    .QN(_01155_),
    .RESETN(net154),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[31]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[31] ),
    .QN(_01159_),
    .RESETN(net155),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[3]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[3] ),
    .QN(_10110_),
    .RESETN(net156),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[4]$_DFF_PP0_  (.CLK(clknet_leaf_2_clk_regs),
    .D(\riscv.dp.ISRmux.d0[4] ),
    .QN(_01077_),
    .RESETN(net157),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[5]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[5] ),
    .QN(_01080_),
    .RESETN(net158),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[6]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[6] ),
    .QN(_01083_),
    .RESETN(net159),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[7]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[7] ),
    .QN(_01086_),
    .RESETN(net160),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[8]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[8] ),
    .QN(_01089_),
    .RESETN(net161),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[9]$_DFF_PP0_  (.CLK(clknet_leaf_3_clk_regs),
    .D(\riscv.dp.ISRmux.d0[9] ),
    .QN(_01092_),
    .RESETN(net162),
    .SETN(_01219_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01222_),
    .QN(_00000_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01223_),
    .QN(_00732_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01224_),
    .QN(_00699_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01225_),
    .QN(_00666_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01226_),
    .QN(_00633_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01227_),
    .QN(_00600_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01228_),
    .QN(_00566_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01229_),
    .QN(_00533_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01230_),
    .QN(_00500_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_01231_),
    .QN(_00467_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_01232_),
    .QN(_00434_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_01233_),
    .QN(_01031_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_01234_),
    .QN(_00401_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_01235_),
    .QN(_00368_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01236_),
    .QN(_00335_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01237_),
    .QN(_00301_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01238_),
    .QN(_00268_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01239_),
    .QN(_00235_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_01240_),
    .QN(_00202_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01241_),
    .QN(_00168_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01242_),
    .QN(_00135_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_01243_),
    .QN(_00101_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01244_),
    .QN(_00998_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_01245_),
    .QN(_00067_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01246_),
    .QN(_00035_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01247_),
    .QN(_00965_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01248_),
    .QN(_00932_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01249_),
    .QN(_00898_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01250_),
    .QN(_00865_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_01251_),
    .QN(_00831_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01252_),
    .QN(_00798_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01253_),
    .QN(_00764_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01254_),
    .QN(_00010_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01255_),
    .QN(_00742_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01256_),
    .QN(_00709_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01257_),
    .QN(_00676_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01258_),
    .QN(_00643_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01259_),
    .QN(_00610_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][15]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01260_),
    .QN(_00576_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][16]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01261_),
    .QN(_00543_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][17]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01262_),
    .QN(_00510_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][18]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01263_),
    .QN(_00477_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][19]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01264_),
    .QN(_00444_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01265_),
    .QN(_01041_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][20]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01266_),
    .QN(_00411_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01267_),
    .QN(_00378_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][22]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01268_),
    .QN(_00345_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][23]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01269_),
    .QN(_00311_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][24]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01270_),
    .QN(_00278_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][25]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01271_),
    .QN(_00245_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][26]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01272_),
    .QN(_00212_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][27]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01273_),
    .QN(_00178_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][28]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01274_),
    .QN(_00145_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01275_),
    .QN(_00111_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01276_),
    .QN(_01008_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][30]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01277_),
    .QN(_00077_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][31]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01278_),
    .QN(_00045_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01279_),
    .QN(_00975_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01280_),
    .QN(_00942_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01281_),
    .QN(_00908_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01282_),
    .QN(_00875_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01283_),
    .QN(_00841_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01284_),
    .QN(_00808_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01285_),
    .QN(_00774_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01286_),
    .QN(_00011_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01287_),
    .QN(_00743_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01288_),
    .QN(_00710_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01289_),
    .QN(_00677_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01290_),
    .QN(_00644_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01291_),
    .QN(_00611_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][15]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01292_),
    .QN(_00577_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01293_),
    .QN(_00544_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01294_),
    .QN(_00511_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][18]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01295_),
    .QN(_00478_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][19]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01296_),
    .QN(_00445_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01297_),
    .QN(_01042_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][20]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01298_),
    .QN(_00412_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01299_),
    .QN(_00379_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][22]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01300_),
    .QN(_00346_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][23]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01301_),
    .QN(_00312_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][24]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01302_),
    .QN(_00279_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][25]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01303_),
    .QN(_00246_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][26]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01304_),
    .QN(_00213_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01305_),
    .QN(_00179_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][28]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01306_),
    .QN(_00146_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01307_),
    .QN(_00112_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01308_),
    .QN(_01009_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][30]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01309_),
    .QN(_00078_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][31]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01310_),
    .QN(_00046_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01311_),
    .QN(_00976_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01312_),
    .QN(_00943_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01313_),
    .QN(_00909_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01314_),
    .QN(_00876_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01315_),
    .QN(_00842_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01316_),
    .QN(_00809_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01317_),
    .QN(_00775_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01318_),
    .QN(_00012_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01319_),
    .QN(_00744_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01320_),
    .QN(_00711_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01321_),
    .QN(_00678_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01322_),
    .QN(_00645_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][14]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01323_),
    .QN(_00612_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][15]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01324_),
    .QN(_00578_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][16]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01325_),
    .QN(_00545_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][17]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01326_),
    .QN(_00512_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][18]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01327_),
    .QN(_00479_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][19]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01328_),
    .QN(_00446_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01329_),
    .QN(_01043_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][20]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01330_),
    .QN(_00413_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01331_),
    .QN(_00380_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][22]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01332_),
    .QN(_00347_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][23]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01333_),
    .QN(_00313_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][24]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01334_),
    .QN(_00280_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][25]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01335_),
    .QN(_00247_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][26]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01336_),
    .QN(_00214_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][27]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01337_),
    .QN(_00180_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][28]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01338_),
    .QN(_00147_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01339_),
    .QN(_00113_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01340_),
    .QN(_01010_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][30]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01341_),
    .QN(_00079_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][31]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01342_),
    .QN(_00047_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01343_),
    .QN(_00977_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01344_),
    .QN(_00944_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01345_),
    .QN(_00910_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01346_),
    .QN(_00877_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01347_),
    .QN(_00843_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01348_),
    .QN(_00810_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01349_),
    .QN(_00776_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01350_),
    .QN(_00013_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01351_),
    .QN(_00745_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01352_),
    .QN(_00712_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01353_),
    .QN(_00679_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01354_),
    .QN(_00646_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01355_),
    .QN(_00613_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][15]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01356_),
    .QN(_00579_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][16]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01357_),
    .QN(_00546_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01358_),
    .QN(_00513_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][18]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01359_),
    .QN(_00480_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][19]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01360_),
    .QN(_00447_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01361_),
    .QN(_01044_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][20]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01362_),
    .QN(_00414_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01363_),
    .QN(_00381_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][22]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01364_),
    .QN(_00348_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][23]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01365_),
    .QN(_00314_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][24]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01366_),
    .QN(_00281_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][25]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01367_),
    .QN(_00248_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][26]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01368_),
    .QN(_00215_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01369_),
    .QN(_00181_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][28]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01370_),
    .QN(_00148_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01371_),
    .QN(_00114_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01372_),
    .QN(_01011_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][30]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01373_),
    .QN(_00080_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][31]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01374_),
    .QN(_00048_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01375_),
    .QN(_00978_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01376_),
    .QN(_00945_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01377_),
    .QN(_00911_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01378_),
    .QN(_00878_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01379_),
    .QN(_00844_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01380_),
    .QN(_00811_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01381_),
    .QN(_00777_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01382_),
    .QN(_00014_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01383_),
    .QN(_00746_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01384_),
    .QN(_00713_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01385_),
    .QN(_00680_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01386_),
    .QN(_00647_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][14]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01387_),
    .QN(_00614_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][15]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01388_),
    .QN(_00580_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][16]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01389_),
    .QN(_00547_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01390_),
    .QN(_00514_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][18]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01391_),
    .QN(_00481_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][19]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01392_),
    .QN(_00448_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01393_),
    .QN(_01045_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][20]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01394_),
    .QN(_00415_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01395_),
    .QN(_00382_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][22]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01396_),
    .QN(_00349_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][23]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01397_),
    .QN(_00315_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][24]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01398_),
    .QN(_00282_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][25]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01399_),
    .QN(_00249_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][26]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01400_),
    .QN(_00216_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][27]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01401_),
    .QN(_00182_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][28]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01402_),
    .QN(_00149_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][29]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01403_),
    .QN(_00115_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01404_),
    .QN(_01012_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][30]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01405_),
    .QN(_00081_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][31]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01406_),
    .QN(_00049_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01407_),
    .QN(_00979_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01408_),
    .QN(_00946_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01409_),
    .QN(_00912_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01410_),
    .QN(_00879_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01411_),
    .QN(_00845_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01412_),
    .QN(_00812_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01413_),
    .QN(_00778_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01414_),
    .QN(_00015_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01415_),
    .QN(_00747_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01416_),
    .QN(_00714_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01417_),
    .QN(_00681_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01418_),
    .QN(_00648_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01419_),
    .QN(_00615_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][15]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01420_),
    .QN(_00581_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][16]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01421_),
    .QN(_00548_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][17]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01422_),
    .QN(_00515_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][18]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01423_),
    .QN(_00482_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][19]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01424_),
    .QN(_00449_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01425_),
    .QN(_01046_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][20]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01426_),
    .QN(_00416_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][21]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01427_),
    .QN(_00383_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][22]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01428_),
    .QN(_00350_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][23]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01429_),
    .QN(_00316_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][24]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01430_),
    .QN(_00283_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][25]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01431_),
    .QN(_00250_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][26]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01432_),
    .QN(_00217_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][27]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01433_),
    .QN(_00183_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][28]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01434_),
    .QN(_00150_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk_regs),
    .D(_01435_),
    .QN(_00116_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01436_),
    .QN(_01013_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][30]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk_regs),
    .D(_01437_),
    .QN(_00082_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][31]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01438_),
    .QN(_00050_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01439_),
    .QN(_00980_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01440_),
    .QN(_00947_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01441_),
    .QN(_00913_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01442_),
    .QN(_00880_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01443_),
    .QN(_00846_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01444_),
    .QN(_00813_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01445_),
    .QN(_00779_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01446_),
    .QN(_00016_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01447_),
    .QN(_00748_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01448_),
    .QN(_00715_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01449_),
    .QN(_00682_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01450_),
    .QN(_00649_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01451_),
    .QN(_00616_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][15]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01452_),
    .QN(_00582_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01453_),
    .QN(_00549_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][17]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01454_),
    .QN(_00516_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][18]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01455_),
    .QN(_00483_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][19]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01456_),
    .QN(_00450_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01457_),
    .QN(_01047_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][20]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01458_),
    .QN(_00417_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01459_),
    .QN(_00384_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01460_),
    .QN(_00351_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][23]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01461_),
    .QN(_00317_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][24]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01462_),
    .QN(_00284_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01463_),
    .QN(_00251_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][26]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01464_),
    .QN(_00218_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01465_),
    .QN(_00184_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][28]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01466_),
    .QN(_00151_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][29]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01467_),
    .QN(_00117_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01468_),
    .QN(_01014_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][30]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01469_),
    .QN(_00083_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][31]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01470_),
    .QN(_00051_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01471_),
    .QN(_00981_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01472_),
    .QN(_00948_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01473_),
    .QN(_00914_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01474_),
    .QN(_00881_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01475_),
    .QN(_00847_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01476_),
    .QN(_00814_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01477_),
    .QN(_00780_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01478_),
    .QN(_00017_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01479_),
    .QN(_00749_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01480_),
    .QN(_00716_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][12]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01481_),
    .QN(_00683_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01482_),
    .QN(_00650_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01483_),
    .QN(_00617_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][15]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01484_),
    .QN(_00583_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01485_),
    .QN(_00550_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][17]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01486_),
    .QN(_00517_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][18]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01487_),
    .QN(_00484_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][19]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01488_),
    .QN(_00451_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01489_),
    .QN(_01048_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][20]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01490_),
    .QN(_00418_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][21]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01491_),
    .QN(_00385_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01492_),
    .QN(_00352_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][23]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01493_),
    .QN(_00318_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][24]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01494_),
    .QN(_00285_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01495_),
    .QN(_00252_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][26]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01496_),
    .QN(_00219_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01497_),
    .QN(_00185_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][28]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01498_),
    .QN(_00152_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][29]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01499_),
    .QN(_00118_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01500_),
    .QN(_01015_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][30]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01501_),
    .QN(_00084_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01502_),
    .QN(_00052_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01503_),
    .QN(_00982_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01504_),
    .QN(_00949_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01505_),
    .QN(_00915_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01506_),
    .QN(_00882_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01507_),
    .QN(_00848_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01508_),
    .QN(_00815_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01509_),
    .QN(_00781_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01510_),
    .QN(_00018_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01511_),
    .QN(_00750_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01512_),
    .QN(_00717_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01513_),
    .QN(_00684_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01514_),
    .QN(_00651_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01515_),
    .QN(_00618_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][15]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01516_),
    .QN(_00584_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01517_),
    .QN(_00551_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][17]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01518_),
    .QN(_00518_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][18]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01519_),
    .QN(_00485_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][19]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01520_),
    .QN(_00452_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01521_),
    .QN(_01049_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][20]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01522_),
    .QN(_00419_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][21]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01523_),
    .QN(_00386_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01524_),
    .QN(_00353_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][23]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01525_),
    .QN(_00319_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][24]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01526_),
    .QN(_00286_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01527_),
    .QN(_00253_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][26]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01528_),
    .QN(_00220_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01529_),
    .QN(_00186_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][28]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01530_),
    .QN(_00153_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][29]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01531_),
    .QN(_00119_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01532_),
    .QN(_01016_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][30]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01533_),
    .QN(_00085_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][31]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01534_),
    .QN(_00053_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01535_),
    .QN(_00983_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01536_),
    .QN(_00950_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01537_),
    .QN(_00916_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01538_),
    .QN(_00883_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01539_),
    .QN(_00849_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01540_),
    .QN(_00816_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01541_),
    .QN(_00782_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01542_),
    .QN(_00019_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01543_),
    .QN(_00751_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01544_),
    .QN(_00718_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01545_),
    .QN(_00685_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01546_),
    .QN(_00652_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01547_),
    .QN(_00619_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][15]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01548_),
    .QN(_00585_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01549_),
    .QN(_00552_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][17]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01550_),
    .QN(_00519_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][18]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01551_),
    .QN(_00486_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][19]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01552_),
    .QN(_00453_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01553_),
    .QN(_01050_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][20]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01554_),
    .QN(_00420_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][21]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01555_),
    .QN(_00387_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][22]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01556_),
    .QN(_00354_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][23]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01557_),
    .QN(_00320_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][24]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01558_),
    .QN(_00287_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01559_),
    .QN(_00254_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][26]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01560_),
    .QN(_00221_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01561_),
    .QN(_00187_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][28]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01562_),
    .QN(_00154_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][29]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01563_),
    .QN(_00120_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01564_),
    .QN(_01017_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][30]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01565_),
    .QN(_00086_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk_regs),
    .D(_01566_),
    .QN(_00054_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01567_),
    .QN(_00984_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01568_),
    .QN(_00951_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01569_),
    .QN(_00917_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01570_),
    .QN(_00884_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01571_),
    .QN(_00850_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01572_),
    .QN(_00817_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01573_),
    .QN(_00783_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01574_),
    .QN(_00001_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01575_),
    .QN(_00733_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01576_),
    .QN(_00700_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_01577_),
    .QN(_00667_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01578_),
    .QN(_00634_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01579_),
    .QN(_00601_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01580_),
    .QN(_00567_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01581_),
    .QN(_00534_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01582_),
    .QN(_00501_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01583_),
    .QN(_00468_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01584_),
    .QN(_00435_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01585_),
    .QN(_01032_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk_regs),
    .D(_01586_),
    .QN(_00402_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01587_),
    .QN(_00369_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01588_),
    .QN(_00336_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01589_),
    .QN(_00302_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk_regs),
    .D(_01590_),
    .QN(_00269_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01591_),
    .QN(_00236_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01592_),
    .QN(_00203_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01593_),
    .QN(_00169_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01594_),
    .QN(_00136_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01595_),
    .QN(_00102_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01596_),
    .QN(_00999_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01597_),
    .QN(_00068_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01598_),
    .QN(_00036_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01599_),
    .QN(_00966_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01600_),
    .QN(_00933_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01601_),
    .QN(_00899_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01602_),
    .QN(_00866_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01603_),
    .QN(_00832_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01604_),
    .QN(_00799_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_01605_),
    .QN(_00765_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01606_),
    .QN(_00020_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01607_),
    .QN(_00752_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01608_),
    .QN(_00719_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][12]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01609_),
    .QN(_00686_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01610_),
    .QN(_00653_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][14]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01611_),
    .QN(_00620_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][15]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01612_),
    .QN(_00586_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01613_),
    .QN(_00553_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][17]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01614_),
    .QN(_00520_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][18]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01615_),
    .QN(_00487_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][19]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01616_),
    .QN(_00454_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01617_),
    .QN(_01051_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][20]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01618_),
    .QN(_00421_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][21]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01619_),
    .QN(_00388_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][22]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01620_),
    .QN(_00355_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][23]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01621_),
    .QN(_00321_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][24]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01622_),
    .QN(_00288_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][25]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01623_),
    .QN(_00255_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01624_),
    .QN(_00222_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01625_),
    .QN(_00188_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01626_),
    .QN(_00155_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][29]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01627_),
    .QN(_00121_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01628_),
    .QN(_01018_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01629_),
    .QN(_00087_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][31]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01630_),
    .QN(_00055_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01631_),
    .QN(_00985_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01632_),
    .QN(_00952_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01633_),
    .QN(_00918_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01634_),
    .QN(_00885_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01635_),
    .QN(_00851_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01636_),
    .QN(_00818_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01637_),
    .QN(_00784_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01638_),
    .QN(_00021_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01639_),
    .QN(_00753_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01640_),
    .QN(_00720_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01641_),
    .QN(_00687_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01642_),
    .QN(_00654_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01643_),
    .QN(_00621_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][15]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01644_),
    .QN(_00587_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01645_),
    .QN(_00554_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][17]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01646_),
    .QN(_00521_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][18]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01647_),
    .QN(_00488_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][19]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01648_),
    .QN(_00455_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01649_),
    .QN(_01052_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][20]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01650_),
    .QN(_00422_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01651_),
    .QN(_00389_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][22]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01652_),
    .QN(_00356_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][23]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01653_),
    .QN(_00322_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][24]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01654_),
    .QN(_00289_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][25]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01655_),
    .QN(_00256_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01656_),
    .QN(_00223_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01657_),
    .QN(_00189_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][28]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01658_),
    .QN(_00156_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][29]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01659_),
    .QN(_00122_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01660_),
    .QN(_01019_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01661_),
    .QN(_00088_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01662_),
    .QN(_00056_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01663_),
    .QN(_00986_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01664_),
    .QN(_00953_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01665_),
    .QN(_00919_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01666_),
    .QN(_00886_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01667_),
    .QN(_00852_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01668_),
    .QN(_00819_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01669_),
    .QN(_00785_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01670_),
    .QN(_00022_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01671_),
    .QN(_00754_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01672_),
    .QN(_00721_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01673_),
    .QN(_00688_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][13]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01674_),
    .QN(_00655_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][14]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01675_),
    .QN(_00622_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][15]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01676_),
    .QN(_00588_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01677_),
    .QN(_00555_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][17]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01678_),
    .QN(_00522_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][18]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01679_),
    .QN(_00489_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][19]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01680_),
    .QN(_00456_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01681_),
    .QN(_01053_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][20]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01682_),
    .QN(_00423_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk_regs),
    .D(_01683_),
    .QN(_00390_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][22]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01684_),
    .QN(_00357_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01685_),
    .QN(_00323_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][24]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01686_),
    .QN(_00290_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][25]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01687_),
    .QN(_00257_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][26]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01688_),
    .QN(_00224_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01689_),
    .QN(_00190_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01690_),
    .QN(_00157_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][29]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01691_),
    .QN(_00123_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01692_),
    .QN(_01020_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01693_),
    .QN(_00089_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01694_),
    .QN(_00057_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01695_),
    .QN(_00987_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01696_),
    .QN(_00954_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01697_),
    .QN(_00920_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01698_),
    .QN(_00887_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01699_),
    .QN(_00853_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01700_),
    .QN(_00820_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01701_),
    .QN(_00786_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01702_),
    .QN(_00023_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01703_),
    .QN(_00755_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01704_),
    .QN(_00722_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01705_),
    .QN(_00689_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01706_),
    .QN(_00656_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][14]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01707_),
    .QN(_00623_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][15]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01708_),
    .QN(_00589_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01709_),
    .QN(_00556_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][17]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01710_),
    .QN(_00523_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][18]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01711_),
    .QN(_00490_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][19]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01712_),
    .QN(_00457_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01713_),
    .QN(_01054_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][20]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01714_),
    .QN(_00424_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01715_),
    .QN(_00391_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01716_),
    .QN(_00358_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][23]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01717_),
    .QN(_00324_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][24]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01718_),
    .QN(_00291_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][25]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01719_),
    .QN(_00258_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01720_),
    .QN(_00225_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01721_),
    .QN(_00191_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01722_),
    .QN(_00158_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][29]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01723_),
    .QN(_00124_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01724_),
    .QN(_01021_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01725_),
    .QN(_00090_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][31]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01726_),
    .QN(_00058_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01727_),
    .QN(_00988_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01728_),
    .QN(_00955_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01729_),
    .QN(_00921_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01730_),
    .QN(_00888_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01731_),
    .QN(_00854_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01732_),
    .QN(_00821_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01733_),
    .QN(_00787_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01734_),
    .QN(_00024_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01735_),
    .QN(_00756_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01736_),
    .QN(_00723_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01737_),
    .QN(_00690_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][13]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01738_),
    .QN(_00657_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01739_),
    .QN(_00624_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][15]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01740_),
    .QN(_00590_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01741_),
    .QN(_00557_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][17]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01742_),
    .QN(_00524_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][18]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01743_),
    .QN(_00491_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][19]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01744_),
    .QN(_00458_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01745_),
    .QN(_01055_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][20]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01746_),
    .QN(_00425_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01747_),
    .QN(_00392_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][22]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01748_),
    .QN(_00359_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][23]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01749_),
    .QN(_00325_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][24]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01750_),
    .QN(_00292_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][25]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01751_),
    .QN(_00259_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01752_),
    .QN(_00226_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01753_),
    .QN(_00192_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][28]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01754_),
    .QN(_00159_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][29]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01755_),
    .QN(_00125_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01756_),
    .QN(_01022_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01757_),
    .QN(_00091_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][31]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01758_),
    .QN(_00059_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01759_),
    .QN(_00989_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01760_),
    .QN(_00956_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01761_),
    .QN(_00922_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01762_),
    .QN(_00889_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01763_),
    .QN(_00855_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01764_),
    .QN(_00822_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01765_),
    .QN(_00788_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01766_),
    .QN(_00025_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01767_),
    .QN(_00757_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01768_),
    .QN(_00724_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01769_),
    .QN(_00691_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01770_),
    .QN(_00658_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01771_),
    .QN(_00625_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][15]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01772_),
    .QN(_00591_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][16]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01773_),
    .QN(_00558_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][17]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01774_),
    .QN(_00525_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][18]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01775_),
    .QN(_00492_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][19]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01776_),
    .QN(_00459_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01777_),
    .QN(_01056_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][20]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01778_),
    .QN(_00426_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01779_),
    .QN(_00393_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][22]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01780_),
    .QN(_00360_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][23]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01781_),
    .QN(_00326_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][24]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01782_),
    .QN(_00293_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][25]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01783_),
    .QN(_00260_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][26]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01784_),
    .QN(_00227_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01785_),
    .QN(_00193_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01786_),
    .QN(_00160_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][29]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01787_),
    .QN(_00126_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01788_),
    .QN(_01023_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01789_),
    .QN(_00092_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01790_),
    .QN(_00060_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01791_),
    .QN(_00990_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01792_),
    .QN(_00957_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01793_),
    .QN(_00923_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01794_),
    .QN(_00890_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01795_),
    .QN(_00856_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01796_),
    .QN(_00823_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01797_),
    .QN(_00789_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01798_),
    .QN(_00026_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01799_),
    .QN(_00758_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01800_),
    .QN(_00725_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][12]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01801_),
    .QN(_00692_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01802_),
    .QN(_00659_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01803_),
    .QN(_00626_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][15]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01804_),
    .QN(_00592_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01805_),
    .QN(_00559_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][17]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01806_),
    .QN(_00526_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][18]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01807_),
    .QN(_00493_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][19]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01808_),
    .QN(_00460_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01809_),
    .QN(_01057_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][20]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01810_),
    .QN(_00427_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][21]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01811_),
    .QN(_00394_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][22]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01812_),
    .QN(_00361_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][23]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk_regs),
    .D(_01813_),
    .QN(_00327_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][24]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01814_),
    .QN(_00294_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][25]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01815_),
    .QN(_00261_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01816_),
    .QN(_00228_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01817_),
    .QN(_00194_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][28]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01818_),
    .QN(_00161_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][29]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01819_),
    .QN(_00127_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01820_),
    .QN(_01024_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01821_),
    .QN(_00093_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][31]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01822_),
    .QN(_00061_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01823_),
    .QN(_00991_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01824_),
    .QN(_00958_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01825_),
    .QN(_00924_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01826_),
    .QN(_00891_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01827_),
    .QN(_00857_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01828_),
    .QN(_00824_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01829_),
    .QN(_00790_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01830_),
    .QN(_00027_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01831_),
    .QN(_00759_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01832_),
    .QN(_00726_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01833_),
    .QN(_00693_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01834_),
    .QN(_00660_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][14]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01835_),
    .QN(_00627_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][15]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01836_),
    .QN(_00593_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01837_),
    .QN(_00560_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][17]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01838_),
    .QN(_00527_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][18]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01839_),
    .QN(_00494_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][19]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01840_),
    .QN(_00461_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01841_),
    .QN(_01058_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][20]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01842_),
    .QN(_00428_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][21]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01843_),
    .QN(_00395_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][22]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01844_),
    .QN(_00362_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][23]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01845_),
    .QN(_00328_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][24]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01846_),
    .QN(_00295_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][25]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01847_),
    .QN(_00262_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01848_),
    .QN(_00229_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01849_),
    .QN(_00195_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01850_),
    .QN(_00162_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][29]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01851_),
    .QN(_00128_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01852_),
    .QN(_01025_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][30]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk_regs),
    .D(_01853_),
    .QN(_00094_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][31]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01854_),
    .QN(_00062_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01855_),
    .QN(_00992_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01856_),
    .QN(_00959_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01857_),
    .QN(_00925_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01858_),
    .QN(_00892_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01859_),
    .QN(_00858_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01860_),
    .QN(_00825_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01861_),
    .QN(_00791_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01862_),
    .QN(_00028_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01863_),
    .QN(_00760_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01864_),
    .QN(_00727_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][12]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_01865_),
    .QN(_00694_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01866_),
    .QN(_00661_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01867_),
    .QN(_00628_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][15]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01868_),
    .QN(_00594_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk_regs),
    .D(_01869_),
    .QN(_00561_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][17]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01870_),
    .QN(_00528_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][18]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01871_),
    .QN(_00495_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][19]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01872_),
    .QN(_00462_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01873_),
    .QN(_01059_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][20]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk_regs),
    .D(_01874_),
    .QN(_00429_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][21]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01875_),
    .QN(_00396_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][22]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01876_),
    .QN(_00363_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01877_),
    .QN(_00329_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][24]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk_regs),
    .D(_01878_),
    .QN(_00296_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][25]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01879_),
    .QN(_00263_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][26]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01880_),
    .QN(_00230_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01881_),
    .QN(_00196_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][28]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01882_),
    .QN(_00163_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][29]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01883_),
    .QN(_00129_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01884_),
    .QN(_01026_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][30]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01885_),
    .QN(_00095_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk_regs),
    .D(_01886_),
    .QN(_00063_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01887_),
    .QN(_00993_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01888_),
    .QN(_00960_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk_regs),
    .D(_01889_),
    .QN(_00926_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01890_),
    .QN(_00893_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01891_),
    .QN(_00859_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01892_),
    .QN(_00826_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk_regs),
    .D(_01893_),
    .QN(_00792_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01894_),
    .QN(_00029_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01895_),
    .QN(_00761_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01896_),
    .QN(_00728_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_01897_),
    .QN(_00695_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][13]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01898_),
    .QN(_00662_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk_regs),
    .D(_01899_),
    .QN(_00629_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][15]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_01900_),
    .QN(_00595_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][16]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01901_),
    .QN(_00562_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][17]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01902_),
    .QN(_00529_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][18]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01903_),
    .QN(_00496_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][19]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01904_),
    .QN(_00463_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01905_),
    .QN(_01060_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][20]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01906_),
    .QN(_00430_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][21]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk_regs),
    .D(_01907_),
    .QN(_00397_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][22]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01908_),
    .QN(_00364_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][23]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01909_),
    .QN(_00330_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][24]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01910_),
    .QN(_00297_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][25]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01911_),
    .QN(_00264_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][26]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01912_),
    .QN(_00231_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_01913_),
    .QN(_00197_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][28]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01914_),
    .QN(_00164_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][29]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01915_),
    .QN(_00130_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01916_),
    .QN(_01027_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][30]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_01917_),
    .QN(_00096_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01918_),
    .QN(_00064_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_01919_),
    .QN(_00994_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk_regs),
    .D(_01920_),
    .QN(_00961_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01921_),
    .QN(_00927_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01922_),
    .QN(_00894_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_01923_),
    .QN(_00860_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk_regs),
    .D(_01924_),
    .QN(_00827_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_01925_),
    .QN(_00793_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01926_),
    .QN(_00002_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01927_),
    .QN(_00734_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01928_),
    .QN(_00701_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01929_),
    .QN(_00668_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_01930_),
    .QN(_00635_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01931_),
    .QN(_00602_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_01932_),
    .QN(_00568_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_01933_),
    .QN(_00535_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_01934_),
    .QN(_00502_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_01935_),
    .QN(_00469_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_01936_),
    .QN(_00436_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01937_),
    .QN(_01033_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_01938_),
    .QN(_00403_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_01939_),
    .QN(_00370_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_01940_),
    .QN(_00337_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_01941_),
    .QN(_00303_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_01942_),
    .QN(_00270_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_01943_),
    .QN(_00237_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_01944_),
    .QN(_00204_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01945_),
    .QN(_00170_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_01946_),
    .QN(_00137_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_01947_),
    .QN(_00103_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_01948_),
    .QN(_01000_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_01949_),
    .QN(_00069_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_01950_),
    .QN(_00037_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_01951_),
    .QN(_00967_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_01952_),
    .QN(_00934_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_01953_),
    .QN(_00900_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_01954_),
    .QN(_00867_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_01955_),
    .QN(_00833_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_01956_),
    .QN(_00800_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_01957_),
    .QN(_00766_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01958_),
    .QN(_00030_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01959_),
    .QN(_00762_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01960_),
    .QN(_00729_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01961_),
    .QN(_00696_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][13]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01962_),
    .QN(_00663_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01963_),
    .QN(_00630_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][15]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01964_),
    .QN(_00596_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][16]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_01965_),
    .QN(_00563_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01966_),
    .QN(_00530_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][18]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_01967_),
    .QN(_00497_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][19]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_01968_),
    .QN(_00464_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01969_),
    .QN(_01061_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][20]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_01970_),
    .QN(_00431_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][21]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_01971_),
    .QN(_00398_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][22]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_01972_),
    .QN(_00365_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][23]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_01973_),
    .QN(_00331_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][24]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_01974_),
    .QN(_00298_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][25]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_01975_),
    .QN(_00265_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][26]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_01976_),
    .QN(_00232_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][27]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01977_),
    .QN(_00198_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][28]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_01978_),
    .QN(_00165_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][29]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_01979_),
    .QN(_00131_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01980_),
    .QN(_01028_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][30]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_01981_),
    .QN(_00097_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01982_),
    .QN(_00065_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01983_),
    .QN(_00995_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01984_),
    .QN(_00962_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_01985_),
    .QN(_00928_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_01986_),
    .QN(_00895_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_01987_),
    .QN(_00861_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_01988_),
    .QN(_00828_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_01989_),
    .QN(_00794_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01990_),
    .QN(_00031_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01991_),
    .QN(_00763_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01992_),
    .QN(_00730_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_01993_),
    .QN(_00697_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][13]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_01994_),
    .QN(_00664_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01995_),
    .QN(_00631_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][15]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_01996_),
    .QN(_00597_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][16]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_01997_),
    .QN(_00564_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01998_),
    .QN(_00531_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][18]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_01999_),
    .QN(_00498_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][19]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02000_),
    .QN(_00465_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_02001_),
    .QN(_01062_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][20]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02002_),
    .QN(_00432_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02003_),
    .QN(_00399_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][22]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02004_),
    .QN(_00366_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][23]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02005_),
    .QN(_00332_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][24]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02006_),
    .QN(_00299_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][25]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_02007_),
    .QN(_00266_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][26]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_02008_),
    .QN(_00233_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][27]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_02009_),
    .QN(_00199_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][28]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_02010_),
    .QN(_00166_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][29]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_02011_),
    .QN(_00132_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_02012_),
    .QN(_01029_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][30]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk_regs),
    .D(_02013_),
    .QN(_00098_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk_regs),
    .D(_02014_),
    .QN(_00066_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_02015_),
    .QN(_00996_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_02016_),
    .QN(_00963_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_02017_),
    .QN(_00929_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_02018_),
    .QN(_00896_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk_regs),
    .D(_02019_),
    .QN(_00862_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk_regs),
    .D(_02020_),
    .QN(_00829_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_02021_),
    .QN(_00795_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02022_),
    .QN(_00003_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02023_),
    .QN(_00735_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02024_),
    .QN(_00702_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02025_),
    .QN(_00669_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02026_),
    .QN(_00636_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02027_),
    .QN(_00603_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02028_),
    .QN(_00569_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02029_),
    .QN(_00536_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02030_),
    .QN(_00503_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02031_),
    .QN(_00470_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02032_),
    .QN(_00437_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02033_),
    .QN(_01034_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02034_),
    .QN(_00404_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02035_),
    .QN(_00371_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02036_),
    .QN(_00338_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02037_),
    .QN(_00304_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02038_),
    .QN(_00271_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02039_),
    .QN(_00238_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02040_),
    .QN(_00205_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02041_),
    .QN(_00171_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02042_),
    .QN(_00138_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02043_),
    .QN(_00104_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02044_),
    .QN(_01001_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02045_),
    .QN(_00070_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02046_),
    .QN(_00038_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02047_),
    .QN(_00968_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk_regs),
    .D(_02048_),
    .QN(_00935_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02049_),
    .QN(_00901_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02050_),
    .QN(_00868_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02051_),
    .QN(_00834_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk_regs),
    .D(_02052_),
    .QN(_00801_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02053_),
    .QN(_00767_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02054_),
    .QN(_00004_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02055_),
    .QN(_00736_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02056_),
    .QN(_00703_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02057_),
    .QN(_00670_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02058_),
    .QN(_00637_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02059_),
    .QN(_00604_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02060_),
    .QN(_00570_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02061_),
    .QN(_00537_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02062_),
    .QN(_00504_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02063_),
    .QN(_00471_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02064_),
    .QN(_00438_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02065_),
    .QN(_01035_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02066_),
    .QN(_00405_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02067_),
    .QN(_00372_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02068_),
    .QN(_00339_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02069_),
    .QN(_00305_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_02070_),
    .QN(_00272_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02071_),
    .QN(_00239_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_02072_),
    .QN(_00206_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02073_),
    .QN(_00172_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02074_),
    .QN(_00139_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_02075_),
    .QN(_00105_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02076_),
    .QN(_01002_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02077_),
    .QN(_00071_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02078_),
    .QN(_00039_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02079_),
    .QN(_00969_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02080_),
    .QN(_00936_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02081_),
    .QN(_00902_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02082_),
    .QN(_00869_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02083_),
    .QN(_00835_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02084_),
    .QN(_00802_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02085_),
    .QN(_00768_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02086_),
    .QN(_00005_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02087_),
    .QN(_00737_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02088_),
    .QN(_00704_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02089_),
    .QN(_00671_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02090_),
    .QN(_00638_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02091_),
    .QN(_00605_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02092_),
    .QN(_00571_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02093_),
    .QN(_00538_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02094_),
    .QN(_00505_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02095_),
    .QN(_00472_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02096_),
    .QN(_00439_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02097_),
    .QN(_01036_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02098_),
    .QN(_00406_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02099_),
    .QN(_00373_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02100_),
    .QN(_00340_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02101_),
    .QN(_00306_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02102_),
    .QN(_00273_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02103_),
    .QN(_00240_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02104_),
    .QN(_00207_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02105_),
    .QN(_00173_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02106_),
    .QN(_00140_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02107_),
    .QN(_00106_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02108_),
    .QN(_01003_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02109_),
    .QN(_00072_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02110_),
    .QN(_00040_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02111_),
    .QN(_00970_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02112_),
    .QN(_00937_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02113_),
    .QN(_00903_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02114_),
    .QN(_00870_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02115_),
    .QN(_00836_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk_regs),
    .D(_02116_),
    .QN(_00803_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02117_),
    .QN(_00769_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02118_),
    .QN(_00006_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02119_),
    .QN(_00738_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02120_),
    .QN(_00705_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02121_),
    .QN(_00672_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02122_),
    .QN(_00639_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02123_),
    .QN(_00606_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02124_),
    .QN(_00572_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02125_),
    .QN(_00539_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02126_),
    .QN(_00506_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02127_),
    .QN(_00473_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02128_),
    .QN(_00440_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02129_),
    .QN(_01037_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02130_),
    .QN(_00407_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02131_),
    .QN(_00374_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02132_),
    .QN(_00341_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02133_),
    .QN(_00307_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02134_),
    .QN(_00274_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02135_),
    .QN(_00241_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_02136_),
    .QN(_00208_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02137_),
    .QN(_00174_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02138_),
    .QN(_00141_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02139_),
    .QN(_00107_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02140_),
    .QN(_01004_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02141_),
    .QN(_00073_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02142_),
    .QN(_00041_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02143_),
    .QN(_00971_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02144_),
    .QN(_00938_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02145_),
    .QN(_00904_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02146_),
    .QN(_00871_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02147_),
    .QN(_00837_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02148_),
    .QN(_00804_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02149_),
    .QN(_00770_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02150_),
    .QN(_00007_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk_regs),
    .D(_02151_),
    .QN(_00739_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02152_),
    .QN(_00706_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02153_),
    .QN(_00673_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02154_),
    .QN(_00640_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02155_),
    .QN(_00607_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02156_),
    .QN(_00573_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02157_),
    .QN(_00540_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02158_),
    .QN(_00507_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02159_),
    .QN(_00474_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02160_),
    .QN(_00441_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02161_),
    .QN(_01038_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02162_),
    .QN(_00408_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02163_),
    .QN(_00375_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02164_),
    .QN(_00342_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02165_),
    .QN(_00308_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02166_),
    .QN(_00275_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02167_),
    .QN(_00242_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_02168_),
    .QN(_00209_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02169_),
    .QN(_00175_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02170_),
    .QN(_00142_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02171_),
    .QN(_00108_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02172_),
    .QN(_01005_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02173_),
    .QN(_00074_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02174_),
    .QN(_00042_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02175_),
    .QN(_00972_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk_regs),
    .D(_02176_),
    .QN(_00939_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02177_),
    .QN(_00905_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02178_),
    .QN(_00872_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02179_),
    .QN(_00838_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk_regs),
    .D(_02180_),
    .QN(_00805_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk_regs),
    .D(_02181_),
    .QN(_00771_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_02182_),
    .QN(_00008_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_02183_),
    .QN(_00740_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_02184_),
    .QN(_00707_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][12]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk_regs),
    .D(_02185_),
    .QN(_00674_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][13]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_02186_),
    .QN(_00641_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][14]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_02187_),
    .QN(_00608_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][15]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_02188_),
    .QN(_00574_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][16]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02189_),
    .QN(_00541_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02190_),
    .QN(_00508_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][18]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02191_),
    .QN(_00475_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][19]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02192_),
    .QN(_00442_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_02193_),
    .QN(_01039_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][20]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02194_),
    .QN(_00409_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][21]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02195_),
    .QN(_00376_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][22]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02196_),
    .QN(_00343_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][23]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02197_),
    .QN(_00309_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][24]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02198_),
    .QN(_00276_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][25]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02199_),
    .QN(_00243_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][26]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02200_),
    .QN(_00210_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][27]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_02201_),
    .QN(_00176_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][28]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk_regs),
    .D(_02202_),
    .QN(_00143_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][29]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02203_),
    .QN(_00109_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_02204_),
    .QN(_01006_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][30]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk_regs),
    .D(_02205_),
    .QN(_00075_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02206_),
    .QN(_00043_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk_regs),
    .D(_02207_),
    .QN(_00973_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_02208_),
    .QN(_00940_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_02209_),
    .QN(_00906_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_02210_),
    .QN(_00873_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_02211_),
    .QN(_00839_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk_regs),
    .D(_02212_),
    .QN(_00806_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_02213_),
    .QN(_00772_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk_regs),
    .D(_02214_),
    .QN(_00009_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_02215_),
    .QN(_00741_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_02216_),
    .QN(_00708_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][12]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_02217_),
    .QN(_00675_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][13]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk_regs),
    .D(_02218_),
    .QN(_00642_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][14]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_02219_),
    .QN(_00609_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][15]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk_regs),
    .D(_02220_),
    .QN(_00575_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][16]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk_regs),
    .D(_02221_),
    .QN(_00542_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][17]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02222_),
    .QN(_00509_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][18]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02223_),
    .QN(_00476_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][19]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02224_),
    .QN(_00443_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_02225_),
    .QN(_01040_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][20]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02226_),
    .QN(_00410_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][21]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02227_),
    .QN(_00377_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][22]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02228_),
    .QN(_00344_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][23]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02229_),
    .QN(_00310_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][24]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02230_),
    .QN(_00277_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][25]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk_regs),
    .D(_02231_),
    .QN(_00244_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][26]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02232_),
    .QN(_00211_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk_regs),
    .D(_02233_),
    .QN(_00177_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][28]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk_regs),
    .D(_02234_),
    .QN(_00144_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][29]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk_regs),
    .D(_02235_),
    .QN(_00110_));
 DFFHQNx3_ASAP7_75t_R \riscv.dp.rf.rf[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk_regs),
    .D(_02236_),
    .QN(_01007_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][30]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk_regs),
    .D(_02237_),
    .QN(_00076_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][31]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk_regs),
    .D(_02238_),
    .QN(_00044_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk_regs),
    .D(_02239_),
    .QN(_00974_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk_regs),
    .D(_02240_),
    .QN(_00941_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk_regs),
    .D(_02241_),
    .QN(_00907_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_02242_),
    .QN(_00874_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk_regs),
    .D(_02243_),
    .QN(_00840_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk_regs),
    .D(_02244_),
    .QN(_00807_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk_regs),
    .D(_02245_),
    .QN(_00773_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Left_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Left_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Left_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Left_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Left_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Left_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Left_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Left_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Left_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Left_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Left_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Left_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Left_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Left_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Left_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Left_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Left_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Left_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Left_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Left_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Left_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Left_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Left_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Left_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Left_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Left_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Left_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Left_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Left_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Left_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Left_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Left_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Left_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Left_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Left_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Left_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Left_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Left_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Left_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Left_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Left_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Left_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Left_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Left_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Left_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Left_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Left_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Left_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Left_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Left_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Left_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Left_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Left_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Left_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_4_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_4_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_4_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_4_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_4_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_4_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_4_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_4_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_4_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_4_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_4_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_4_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_4_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_4_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_4_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_4_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_4_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_4_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_4_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_4_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_4_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_4_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_4_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_4_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_4_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_4_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_4_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_4_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_4_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_4_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_4_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_4_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_4_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_4_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_4_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_4_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_4_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_4_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_4_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_4_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_4_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_4_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_4_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_4_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_4_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_4_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_4_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_4_Left_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_4_Left_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_4_Left_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_4_Left_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_4_Left_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_4_Left_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_4_Left_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_4_Left_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_4_Left_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_4_Left_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_4_Left_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_4_Left_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_4_Left_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_4_Left_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_4_Left_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_4_Left_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_4_Left_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_4_Left_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_4_Left_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_4_Left_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_4_Left_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_4_Left_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_4_Left_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_4_Left_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_4_Left_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_4_Left_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_4_Left_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_4_Left_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_4_Left_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_4_Left_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_4_Left_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_4_Left_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_4_Left_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_4_Left_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_4_Left_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_4_Left_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_4_Left_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_4_Left_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_4_Left_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_4_Left_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_4_Left_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_4_Left_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_4_Left_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_4_Left_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_4_Left_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_4_Left_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_4_Left_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_4_Left_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_4_Left_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_4_Left_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_4_Left_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_4_Left_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_4_Left_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_4_Left_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_4_Left_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_4_Left_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_4_Left_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_4_Left_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_4_Left_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_4_Left_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_4_Left_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_4_Left_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_4_Left_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_4_Left_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_4_Left_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_4_Left_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_4_Left_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_4_Left_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_4_Left_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_4_Left_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_4_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_4_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_4_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_4_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_4_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_4_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_4_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_4_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_4_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_4_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_4_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_4_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_4_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_4_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_4_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_4_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_4_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_4_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_4_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_4_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_4_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_4_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_4_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_4_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_4_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_4_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_4_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_4_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_4_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_4_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_4_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_4_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_4_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_4_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_4_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_4_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_4_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_4_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_4_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_4_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_4_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_4_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_4_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_4_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_4_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_4_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_4_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_4_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_4_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_4_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_4_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_4_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_4_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_4_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_4_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_4_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_4_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_4_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_4_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_4_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_4_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_4_Right_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_4_Right_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_4_Right_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_4_Right_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_4_Right_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_4_Right_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_4_Right_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_4_Right_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_4_Right_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_4_Right_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_4_Right_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_4_Right_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_4_Right_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_4_Right_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_4_Right_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_4_Right_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_4_Right_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_4_Right_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_4_Right_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_4_Right_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_4_Right_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_4_Right_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_4_Right_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_4_Right_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_4_Right_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_4_Right_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_4_Right_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_4_Right_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_4_Right_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_4_Right_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_4_Right_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_4_Right_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_4_Right_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_4_Right_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_4_Right_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_4_Right_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_4_Right_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_4_Right_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_4_Right_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_4_Right_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_4_Right_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_4_Right_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_4_Right_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_4_Right_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_4_Right_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_4_Right_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_4_Right_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_4_Right_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_4_Right_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_4_Right_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_4_Right_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_4_Right_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_4_Right_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_4_Right_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_4_Right_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_2_Right_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Right_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Right_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Right_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Right_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Right_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Right_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Right_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Right_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Right_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Right_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Right_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Right_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Right_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Right_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Right_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Right_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Right_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Right_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Right_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Right_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Right_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Right_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Right_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Right_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Right_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Right_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Right_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Right_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Right_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Right_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Right_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Right_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Right_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Right_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Right_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_Right_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_Right_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_Right_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_Right_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_Right_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_Right_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_Right_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_Right_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_Right_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_Right_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Right_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Right_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Right_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Right_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Right_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Right_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Right_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Right_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Right_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Right_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Right_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Right_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_Right_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_Right_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_Right_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_Right_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Right_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_2_Right_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_2_Right_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_2_Right_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_2_Right_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_2_Right_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_2_Right_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_2_Right_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_2_Right_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_2_Right_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_2_Right_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_2_Right_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_2_Right_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_2_Right_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_2_Right_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_2_Right_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_2_Right_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_2_Right_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_2_Right_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_2_Right_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_2_Right_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_2_Right_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_2_Right_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_2_Right_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_2_Right_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_2_Right_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_2_Right_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_2_Right_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_2_Right_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_2_Right_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_2_Right_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_2_Right_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_2_Right_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_2_Right_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_2_Right_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_2_Right_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_2_Right_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_2_Right_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_2_Right_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_2_Right_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_2_Right_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_2_Right_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_2_Right_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_2_Right_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_2_Right_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_2_Right_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_2_Right_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_2_Right_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_2_Right_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_2_Right_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_2_Right_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_2_Right_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_2_Right_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_2_Right_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_2_Right_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_2_Right_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_2_Right_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_2_Right_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_2_Right_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_2_Right_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_2_Right_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_2_Right_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_2_Right_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_2_Right_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_2_Right_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_2_Right_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_2_Right_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_2_Right_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_2_Right_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_2_Right_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_2_Right_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_2_Right_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_2_Right_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_2_Right_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_2_Right_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_2_Right_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_2_Right_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_2_Right_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_2_Right_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_2_Right_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_2_Right_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_2_Right_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_2_Right_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_2_Right_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_2_Right_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_2_Right_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_2_Right_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_2_Right_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_2_Right_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_2_Right_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_2_Right_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_2_Right_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_2_Right_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_2_Right_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_2_Right_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_2_Right_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_2_Right_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_2_Right_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_2_Right_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_2_Right_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_2_Right_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_2_Right_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_2_Right_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_2_Right_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_2_Right_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_2_Right_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_2_Right_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_2_Right_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_2_Right_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_2_Right_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_2_Right_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_2_Right_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_2_Right_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_2_Right_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_2_Right_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_2_Right_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_4_Right_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_2_Left_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_2_Left_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_2_Left_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_2_Left_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_2_Left_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_2_Left_479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_2_Left_480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_2_Left_481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_2_Left_482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_2_Left_483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_2_Left_484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_2_Left_485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_2_Left_486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_2_Left_487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_2_Left_488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_2_Left_489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_2_Left_490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_2_Left_491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_2_Left_492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_2_Left_493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_2_Left_494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_2_Left_495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_2_Left_496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_2_Left_497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_2_Left_498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_2_Left_499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_2_Left_500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_2_Left_501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_2_Left_502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_2_Left_503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_2_Left_504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_2_Left_505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_2_Left_506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_2_Left_507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_2_Left_508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_2_Left_509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_2_Left_510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_2_Left_511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_2_Left_512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_2_Left_513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_2_Left_514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_2_Left_515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_2_Left_516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_2_Left_517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_2_Left_518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_2_Left_519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_2_Left_520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_2_Left_521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_2_Left_522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_2_Left_523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_2_Left_524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_2_Left_525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_2_Left_526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_2_Left_527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_2_Left_528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_2_Left_529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_2_Left_530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_2_Left_531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_2_Left_532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_2_Left_533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_2_Left_534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_2_Left_535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_2_Left_536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_2_Left_537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_2_Left_538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_2_Left_539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_2_Left_540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_2_Left_541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_2_Left_542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_2_Left_543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_2_Left_544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_2_Left_545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_2_Left_546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_2_Left_547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_2_Left_548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_2_Left_549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_2_Left_550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_2_Left_551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_2_Left_552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_2_Left_553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_2_Left_554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_2_Left_555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_2_Left_556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_2_Left_557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_2_Left_558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_2_Left_559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_2_Left_560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_2_Left_561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_2_Left_562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_2_Left_563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_2_Left_564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_2_Left_565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_2_Left_566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_2_Left_567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_2_Left_568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_2_Left_569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_2_Left_570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_2_Left_571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_2_Left_572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_2_Left_573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_2_Left_574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_2_Left_575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_2_Left_576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_2_Left_577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_2_Left_578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_2_Left_579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_2_Left_580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_2_Left_581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_2_Left_582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_2_Left_583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_2_Left_584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_2_Left_585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_2_Left_586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_2_Left_587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_2_Left_588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_2_Left_589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_4_590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_4_591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_4_592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_4_593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_4_594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_4_595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_4_596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_4_597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_4_598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_4_599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_4_600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_4_601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_4_602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_4_603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_4_604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_4_605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_4_606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_4_607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_4_608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_4_609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_4_610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_4_611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_4_612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_4_613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_4_614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_4_615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_4_616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_4_617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_4_618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_4_619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_4_620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_4_621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_4_622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_4_623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_4_624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_4_625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_4_626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_4_627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_4_628 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_4_629 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_4_630 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_4_631 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_4_632 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_4_633 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_4_634 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_4_635 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_4_636 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_4_637 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_4_638 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_4_639 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_4_640 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_4_641 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_4_642 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_4_643 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_4_644 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_4_645 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_4_646 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_4_647 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_2_648 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_117_649 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_117_650 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_651 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_119_652 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_653 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_121_654 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_655 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_123_656 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_657 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_125_658 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_659 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_127_660 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_661 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_129_662 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_663 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_131_664 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_665 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_133_666 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_667 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_135_668 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_669 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_137_670 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_671 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_139_672 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_673 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_141_674 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_675 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_143_676 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_677 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_145_678 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_679 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_147_680 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_681 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_149_682 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_683 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_151_684 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_152_685 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_153_686 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_154_687 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_155_688 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_156_689 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_157_690 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_158_691 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_159_692 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_160_693 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_161_694 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_695 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_163_696 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_697 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_165_698 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_699 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_167_700 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_701 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_169_702 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_703 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_171_704 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_705 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_706 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_174_707 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_175_708 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_176_709 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_177_710 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_711 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_712 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_2_713 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_2_714 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_2_715 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_2_716 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_2_717 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_2_718 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_2_719 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_2_720 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_2_721 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_2_722 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_190_2_723 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_191_2_724 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_192_2_725 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_193_2_726 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_194_2_727 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_195_2_728 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_196_2_729 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_197_2_730 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_198_2_731 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_199_2_732 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_200_2_733 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_201_2_734 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_202_2_735 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_203_2_736 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_204_2_737 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_205_2_738 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_206_2_739 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_207_2_740 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_208_2_741 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_209_2_742 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_210_2_743 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_211_2_744 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_212_2_745 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_213_2_746 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_214_2_747 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_215_2_748 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_216_2_749 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_217_2_750 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_218_2_751 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_219_2_752 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_220_2_753 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_221_2_754 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_222_2_755 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_223_2_756 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_224_2_757 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_225_2_758 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_226_2_759 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_227_2_760 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_228_2_761 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_229_2_762 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_230_2_763 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_231_2_764 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_232_2_765 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_233_2_766 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_234_2_767 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_235_2_768 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_236_2_769 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_237_2_770 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_238_2_771 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_239_2_772 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_240_2_773 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_241_2_774 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_2_775 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_243_2_776 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_244_2_777 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_245_2_778 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_246_2_779 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_247_2_780 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_248_2_781 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_249_2_782 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_250_2_783 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_251_2_784 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_252_2_785 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_253_2_786 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_254_2_787 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_255_2_788 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_256_2_789 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_257_2_790 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_258_2_791 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_259_2_792 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_260_2_793 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_261_2_794 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_262_2_795 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_263_2_796 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_264_2_797 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_265_2_798 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_266_2_799 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_267_2_800 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_268_2_801 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_269_2_802 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_270_2_803 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_271_2_804 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_272_2_805 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_273_2_806 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_274_2_807 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_275_2_808 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_276_2_809 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_277_2_810 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_278_2_811 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_279_2_812 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_280_2_813 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_281_2_814 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_282_2_815 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_283_2_816 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_284_2_817 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_285_2_818 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_286_2_819 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_287_2_820 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_288_2_821 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_289_2_822 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_290_2_823 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_291_2_824 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_292_2_825 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_293_2_826 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_294_2_827 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_294_2_828 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_4_829 ();
 BUFx4f_ASAP7_75t_R input1 (.A(instr[0]),
    .Y(net1));
 BUFx4f_ASAP7_75t_R input2 (.A(instr[10]),
    .Y(net2));
 BUFx3_ASAP7_75t_R input3 (.A(instr[11]),
    .Y(net3));
 BUFx4f_ASAP7_75t_R input4 (.A(instr[12]),
    .Y(net4));
 BUFx3_ASAP7_75t_R input5 (.A(instr[13]),
    .Y(net5));
 BUFx4f_ASAP7_75t_R input6 (.A(instr[14]),
    .Y(net6));
 BUFx6f_ASAP7_75t_R input7 (.A(instr[15]),
    .Y(net7));
 BUFx4f_ASAP7_75t_R input8 (.A(instr[17]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input9 (.A(instr[18]),
    .Y(net9));
 BUFx4f_ASAP7_75t_R input10 (.A(instr[19]),
    .Y(net10));
 BUFx3_ASAP7_75t_R input11 (.A(instr[1]),
    .Y(net11));
 BUFx3_ASAP7_75t_R input12 (.A(instr[20]),
    .Y(net12));
 BUFx4f_ASAP7_75t_R input13 (.A(instr[21]),
    .Y(net13));
 BUFx4f_ASAP7_75t_R input14 (.A(instr[23]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input15 (.A(instr[24]),
    .Y(net15));
 BUFx3_ASAP7_75t_R input16 (.A(instr[25]),
    .Y(net16));
 BUFx3_ASAP7_75t_R input17 (.A(instr[26]),
    .Y(net17));
 BUFx3_ASAP7_75t_R input18 (.A(instr[27]),
    .Y(net18));
 BUFx3_ASAP7_75t_R input19 (.A(instr[28]),
    .Y(net19));
 BUFx3_ASAP7_75t_R input20 (.A(instr[29]),
    .Y(net20));
 BUFx4f_ASAP7_75t_R input21 (.A(instr[2]),
    .Y(net21));
 BUFx6f_ASAP7_75t_R input22 (.A(instr[30]),
    .Y(net22));
 BUFx3_ASAP7_75t_R input23 (.A(instr[31]),
    .Y(net23));
 BUFx4f_ASAP7_75t_R input24 (.A(instr[3]),
    .Y(net24));
 BUFx4f_ASAP7_75t_R input25 (.A(instr[4]),
    .Y(net25));
 BUFx3_ASAP7_75t_R input26 (.A(instr[5]),
    .Y(net26));
 BUFx4f_ASAP7_75t_R input27 (.A(instr[6]),
    .Y(net27));
 BUFx4f_ASAP7_75t_R input28 (.A(instr[7]),
    .Y(net28));
 BUFx3_ASAP7_75t_R input29 (.A(instr[8]),
    .Y(net29));
 BUFx3_ASAP7_75t_R input30 (.A(instr[9]),
    .Y(net30));
 BUFx12f_ASAP7_75t_R input31 (.A(reset),
    .Y(net31));
 BUFx2_ASAP7_75t_R output32 (.A(net32),
    .Y(dataadr[0]));
 BUFx2_ASAP7_75t_R output33 (.A(net33),
    .Y(dataadr[10]));
 BUFx2_ASAP7_75t_R output34 (.A(net34),
    .Y(dataadr[11]));
 BUFx2_ASAP7_75t_R output35 (.A(net35),
    .Y(dataadr[12]));
 BUFx2_ASAP7_75t_R output36 (.A(net36),
    .Y(dataadr[13]));
 BUFx2_ASAP7_75t_R output37 (.A(net37),
    .Y(dataadr[14]));
 BUFx2_ASAP7_75t_R output38 (.A(net38),
    .Y(dataadr[15]));
 BUFx2_ASAP7_75t_R output39 (.A(net39),
    .Y(dataadr[16]));
 BUFx2_ASAP7_75t_R output40 (.A(net40),
    .Y(dataadr[17]));
 BUFx2_ASAP7_75t_R output41 (.A(net41),
    .Y(dataadr[18]));
 BUFx2_ASAP7_75t_R output42 (.A(net42),
    .Y(dataadr[19]));
 BUFx2_ASAP7_75t_R output43 (.A(net43),
    .Y(dataadr[1]));
 BUFx2_ASAP7_75t_R output44 (.A(net44),
    .Y(dataadr[20]));
 BUFx2_ASAP7_75t_R output45 (.A(net45),
    .Y(dataadr[21]));
 BUFx2_ASAP7_75t_R output46 (.A(net46),
    .Y(dataadr[22]));
 BUFx2_ASAP7_75t_R output47 (.A(net47),
    .Y(dataadr[23]));
 BUFx2_ASAP7_75t_R output48 (.A(net48),
    .Y(dataadr[24]));
 BUFx2_ASAP7_75t_R output49 (.A(net49),
    .Y(dataadr[25]));
 BUFx2_ASAP7_75t_R output50 (.A(net50),
    .Y(dataadr[26]));
 BUFx2_ASAP7_75t_R output51 (.A(net51),
    .Y(dataadr[27]));
 BUFx2_ASAP7_75t_R output52 (.A(net52),
    .Y(dataadr[28]));
 BUFx2_ASAP7_75t_R output53 (.A(net53),
    .Y(dataadr[29]));
 BUFx2_ASAP7_75t_R output54 (.A(net54),
    .Y(dataadr[2]));
 BUFx2_ASAP7_75t_R output55 (.A(net55),
    .Y(dataadr[30]));
 BUFx2_ASAP7_75t_R output56 (.A(net56),
    .Y(dataadr[31]));
 BUFx2_ASAP7_75t_R output57 (.A(net57),
    .Y(dataadr[3]));
 BUFx2_ASAP7_75t_R output58 (.A(net58),
    .Y(dataadr[4]));
 BUFx2_ASAP7_75t_R output59 (.A(net59),
    .Y(dataadr[5]));
 BUFx2_ASAP7_75t_R output60 (.A(net60),
    .Y(dataadr[6]));
 BUFx2_ASAP7_75t_R output61 (.A(net61),
    .Y(dataadr[7]));
 BUFx2_ASAP7_75t_R output62 (.A(net62),
    .Y(dataadr[8]));
 BUFx2_ASAP7_75t_R output63 (.A(net63),
    .Y(dataadr[9]));
 BUFx2_ASAP7_75t_R output64 (.A(net64),
    .Y(memwrite));
 BUFx2_ASAP7_75t_R output65 (.A(net65),
    .Y(pc[0]));
 BUFx2_ASAP7_75t_R output66 (.A(net66),
    .Y(pc[10]));
 BUFx2_ASAP7_75t_R output67 (.A(net67),
    .Y(pc[11]));
 BUFx2_ASAP7_75t_R output68 (.A(net68),
    .Y(pc[12]));
 BUFx2_ASAP7_75t_R output69 (.A(net69),
    .Y(pc[13]));
 BUFx2_ASAP7_75t_R output70 (.A(net70),
    .Y(pc[14]));
 BUFx2_ASAP7_75t_R output71 (.A(net71),
    .Y(pc[15]));
 BUFx2_ASAP7_75t_R output72 (.A(net72),
    .Y(pc[16]));
 BUFx2_ASAP7_75t_R output73 (.A(net73),
    .Y(pc[17]));
 BUFx2_ASAP7_75t_R output74 (.A(net74),
    .Y(pc[18]));
 BUFx2_ASAP7_75t_R output75 (.A(net75),
    .Y(pc[19]));
 BUFx2_ASAP7_75t_R output76 (.A(net76),
    .Y(pc[1]));
 BUFx2_ASAP7_75t_R output77 (.A(net77),
    .Y(pc[20]));
 BUFx2_ASAP7_75t_R output78 (.A(net78),
    .Y(pc[21]));
 BUFx2_ASAP7_75t_R output79 (.A(net79),
    .Y(pc[22]));
 BUFx2_ASAP7_75t_R output80 (.A(net80),
    .Y(pc[23]));
 BUFx2_ASAP7_75t_R output81 (.A(net81),
    .Y(pc[24]));
 BUFx2_ASAP7_75t_R output82 (.A(net82),
    .Y(pc[25]));
 BUFx2_ASAP7_75t_R output83 (.A(net83),
    .Y(pc[26]));
 BUFx2_ASAP7_75t_R output84 (.A(net84),
    .Y(pc[27]));
 BUFx2_ASAP7_75t_R output85 (.A(net85),
    .Y(pc[28]));
 BUFx2_ASAP7_75t_R output86 (.A(net86),
    .Y(pc[29]));
 BUFx2_ASAP7_75t_R output87 (.A(net87),
    .Y(pc[2]));
 BUFx2_ASAP7_75t_R output88 (.A(net88),
    .Y(pc[30]));
 BUFx2_ASAP7_75t_R output89 (.A(net89),
    .Y(pc[31]));
 BUFx2_ASAP7_75t_R output90 (.A(net90),
    .Y(pc[3]));
 BUFx2_ASAP7_75t_R output91 (.A(net91),
    .Y(pc[4]));
 BUFx2_ASAP7_75t_R output92 (.A(net92),
    .Y(pc[5]));
 BUFx2_ASAP7_75t_R output93 (.A(net93),
    .Y(pc[6]));
 BUFx2_ASAP7_75t_R output94 (.A(net94),
    .Y(pc[7]));
 BUFx2_ASAP7_75t_R output95 (.A(net95),
    .Y(pc[8]));
 BUFx2_ASAP7_75t_R output96 (.A(net96),
    .Y(pc[9]));
 BUFx2_ASAP7_75t_R output97 (.A(net97),
    .Y(ready));
 BUFx2_ASAP7_75t_R output98 (.A(net98),
    .Y(suspend));
 BUFx2_ASAP7_75t_R output99 (.A(net99),
    .Y(writedata[0]));
 BUFx2_ASAP7_75t_R output100 (.A(net100),
    .Y(writedata[10]));
 BUFx2_ASAP7_75t_R output101 (.A(net101),
    .Y(writedata[11]));
 BUFx2_ASAP7_75t_R output102 (.A(net102),
    .Y(writedata[12]));
 BUFx2_ASAP7_75t_R output103 (.A(net103),
    .Y(writedata[13]));
 BUFx2_ASAP7_75t_R output104 (.A(net104),
    .Y(writedata[14]));
 BUFx2_ASAP7_75t_R output105 (.A(net105),
    .Y(writedata[15]));
 BUFx2_ASAP7_75t_R output106 (.A(net106),
    .Y(writedata[16]));
 BUFx2_ASAP7_75t_R output107 (.A(net107),
    .Y(writedata[17]));
 BUFx2_ASAP7_75t_R output108 (.A(net108),
    .Y(writedata[18]));
 BUFx2_ASAP7_75t_R output109 (.A(net109),
    .Y(writedata[19]));
 BUFx2_ASAP7_75t_R output110 (.A(net110),
    .Y(writedata[1]));
 BUFx2_ASAP7_75t_R output111 (.A(net111),
    .Y(writedata[20]));
 BUFx2_ASAP7_75t_R output112 (.A(net112),
    .Y(writedata[21]));
 BUFx2_ASAP7_75t_R output113 (.A(net113),
    .Y(writedata[22]));
 BUFx2_ASAP7_75t_R output114 (.A(net114),
    .Y(writedata[23]));
 BUFx2_ASAP7_75t_R output115 (.A(net115),
    .Y(writedata[24]));
 BUFx2_ASAP7_75t_R output116 (.A(net116),
    .Y(writedata[25]));
 BUFx2_ASAP7_75t_R output117 (.A(net117),
    .Y(writedata[26]));
 BUFx2_ASAP7_75t_R output118 (.A(net118),
    .Y(writedata[27]));
 BUFx2_ASAP7_75t_R output119 (.A(net119),
    .Y(writedata[28]));
 BUFx2_ASAP7_75t_R output120 (.A(net120),
    .Y(writedata[29]));
 BUFx2_ASAP7_75t_R output121 (.A(net121),
    .Y(writedata[2]));
 BUFx2_ASAP7_75t_R output122 (.A(net122),
    .Y(writedata[30]));
 BUFx2_ASAP7_75t_R output123 (.A(net123),
    .Y(writedata[31]));
 BUFx2_ASAP7_75t_R output124 (.A(net124),
    .Y(writedata[3]));
 BUFx2_ASAP7_75t_R output125 (.A(net125),
    .Y(writedata[4]));
 BUFx2_ASAP7_75t_R output126 (.A(net126),
    .Y(writedata[5]));
 BUFx2_ASAP7_75t_R output127 (.A(net127),
    .Y(writedata[6]));
 BUFx2_ASAP7_75t_R output128 (.A(net128),
    .Y(writedata[7]));
 BUFx2_ASAP7_75t_R output129 (.A(net129),
    .Y(writedata[8]));
 BUFx2_ASAP7_75t_R output130 (.A(net130),
    .Y(writedata[9]));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[0]$_DFFE_PP0P__131  (.H(net131));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[10]$_DFF_PP0__132  (.H(net132));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[11]$_DFF_PP0__133  (.H(net133));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[12]$_DFF_PP0__134  (.H(net134));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[13]$_DFF_PP0__135  (.H(net135));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[14]$_DFF_PP0__136  (.H(net136));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[15]$_DFF_PP0__137  (.H(net137));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[16]$_DFF_PP0__138  (.H(net138));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[17]$_DFF_PP0__139  (.H(net139));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[18]$_DFF_PP0__140  (.H(net140));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[19]$_DFF_PP0__141  (.H(net141));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[1]$_DFFE_PP0P__142  (.H(net142));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[20]$_DFF_PP0__143  (.H(net143));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[21]$_DFF_PP0__144  (.H(net144));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[22]$_DFF_PP0__145  (.H(net145));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[23]$_DFF_PP0__146  (.H(net146));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[24]$_DFF_PP0__147  (.H(net147));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[25]$_DFF_PP0__148  (.H(net148));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[26]$_DFF_PP0__149  (.H(net149));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[27]$_DFF_PP0__150  (.H(net150));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[28]$_DFF_PP0__151  (.H(net151));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[29]$_DFF_PP0__152  (.H(net152));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[2]$_DFF_PP0__153  (.H(net153));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[30]$_DFF_PP0__154  (.H(net154));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[31]$_DFF_PP0__155  (.H(net155));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[3]$_DFF_PP0__156  (.H(net156));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[4]$_DFF_PP0__157  (.H(net157));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[5]$_DFF_PP0__158  (.H(net158));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[6]$_DFF_PP0__159  (.H(net159));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[7]$_DFF_PP0__160  (.H(net160));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[8]$_DFF_PP0__161  (.H(net161));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[9]$_DFF_PP0__162  (.H(net162));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx16f_ASAP7_75t_R clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_0__leaf_clk));
 BUFx16f_ASAP7_75t_R clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_1__leaf_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_0_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_1_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_2_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_3_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_4_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_5_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_6_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_7_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_8_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk_regs (.A(clknet_2_2_0_clk_regs),
    .Y(clknet_leaf_9_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_10_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_11_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_12_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_13_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_14_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_15_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_16_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_17_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_18_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_19_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_20_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_21_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_22_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_23_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_24_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk_regs (.A(clknet_2_3_0_clk_regs),
    .Y(clknet_leaf_25_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_26_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_27_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_28_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_28_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_29_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_29_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_30_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_30_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_31_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_31_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_32_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_32_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_33_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_33_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_34_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_34_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_35_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_35_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_36_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_36_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_37_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_37_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_38_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_38_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_39_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_39_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_40_clk_regs (.A(clknet_2_1_0_clk_regs),
    .Y(clknet_leaf_40_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_41_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_41_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_42_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_42_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_43_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_43_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_44_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_44_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_45_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_45_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_46_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_46_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_47_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_47_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_48_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_48_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_49_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_49_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_50_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_50_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_51_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_51_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_leaf_52_clk_regs (.A(clknet_2_0_0_clk_regs),
    .Y(clknet_leaf_52_clk_regs));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk_regs (.A(clk_regs),
    .Y(clknet_0_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_2_0_0_clk_regs (.A(clknet_0_clk_regs),
    .Y(clknet_2_0_0_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_2_1_0_clk_regs (.A(clknet_0_clk_regs),
    .Y(clknet_2_1_0_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_2_2_0_clk_regs (.A(clknet_0_clk_regs),
    .Y(clknet_2_2_0_clk_regs));
 BUFx24_ASAP7_75t_R clkbuf_2_3_0_clk_regs (.A(clknet_0_clk_regs),
    .Y(clknet_2_3_0_clk_regs));
 CKINVDCx16_ASAP7_75t_R clkload0 (.A(clknet_2_0_0_clk_regs));
 CKINVDCx20_ASAP7_75t_R clkload1 (.A(clknet_2_2_0_clk_regs));
 BUFx24_ASAP7_75t_R clkload2 (.A(clknet_2_3_0_clk_regs));
 BUFx4f_ASAP7_75t_R clkload3 (.A(clknet_leaf_42_clk_regs));
 INVxp33_ASAP7_75t_R clkload4 (.A(clknet_leaf_43_clk_regs));
 INVx6_ASAP7_75t_R clkload5 (.A(clknet_leaf_44_clk_regs));
 INVx8_ASAP7_75t_R clkload6 (.A(clknet_leaf_45_clk_regs));
 CKINVDCx5p33_ASAP7_75t_R clkload7 (.A(clknet_leaf_46_clk_regs));
 INVx5_ASAP7_75t_R clkload8 (.A(clknet_leaf_47_clk_regs));
 INVxp67_ASAP7_75t_R clkload9 (.A(clknet_leaf_48_clk_regs));
 INVx3_ASAP7_75t_R clkload10 (.A(clknet_leaf_49_clk_regs));
 INVx5_ASAP7_75t_R clkload11 (.A(clknet_leaf_50_clk_regs));
 CKINVDCx8_ASAP7_75t_R clkload12 (.A(clknet_leaf_51_clk_regs));
 BUFx12_ASAP7_75t_R clkload13 (.A(clknet_leaf_52_clk_regs));
 CKINVDCx8_ASAP7_75t_R clkload14 (.A(clknet_leaf_26_clk_regs));
 INVx8_ASAP7_75t_R clkload15 (.A(clknet_leaf_27_clk_regs));
 INVx3_ASAP7_75t_R clkload16 (.A(clknet_leaf_28_clk_regs));
 BUFx4f_ASAP7_75t_R clkload17 (.A(clknet_leaf_29_clk_regs));
 BUFx12_ASAP7_75t_R clkload18 (.A(clknet_leaf_30_clk_regs));
 BUFx4f_ASAP7_75t_R clkload19 (.A(clknet_leaf_31_clk_regs));
 INVx8_ASAP7_75t_R clkload20 (.A(clknet_leaf_32_clk_regs));
 INVx3_ASAP7_75t_R clkload21 (.A(clknet_leaf_33_clk_regs));
 BUFx4f_ASAP7_75t_R clkload22 (.A(clknet_leaf_34_clk_regs));
 INVxp67_ASAP7_75t_R clkload23 (.A(clknet_leaf_35_clk_regs));
 BUFx12_ASAP7_75t_R clkload24 (.A(clknet_leaf_36_clk_regs));
 INVx3_ASAP7_75t_R clkload25 (.A(clknet_leaf_37_clk_regs));
 CKINVDCx6p67_ASAP7_75t_R clkload26 (.A(clknet_leaf_38_clk_regs));
 INVx5_ASAP7_75t_R clkload27 (.A(clknet_leaf_39_clk_regs));
 INVxp67_ASAP7_75t_R clkload28 (.A(clknet_leaf_0_clk_regs));
 BUFx24_ASAP7_75t_R clkload29 (.A(clknet_leaf_1_clk_regs));
 INVx5_ASAP7_75t_R clkload30 (.A(clknet_leaf_2_clk_regs));
 CKINVDCx8_ASAP7_75t_R clkload31 (.A(clknet_leaf_3_clk_regs));
 BUFx24_ASAP7_75t_R clkload32 (.A(clknet_leaf_5_clk_regs));
 BUFx24_ASAP7_75t_R clkload33 (.A(clknet_leaf_6_clk_regs));
 BUFx4f_ASAP7_75t_R clkload34 (.A(clknet_leaf_7_clk_regs));
 BUFx24_ASAP7_75t_R clkload35 (.A(clknet_leaf_8_clk_regs));
 CKINVDCx10_ASAP7_75t_R clkload36 (.A(clknet_leaf_9_clk_regs));
 CKINVDCx8_ASAP7_75t_R clkload37 (.A(clknet_leaf_10_clk_regs));
 BUFx4f_ASAP7_75t_R clkload38 (.A(clknet_leaf_11_clk_regs));
 INVx3_ASAP7_75t_R clkload39 (.A(clknet_leaf_12_clk_regs));
 INVx3_ASAP7_75t_R clkload40 (.A(clknet_leaf_14_clk_regs));
 INVxp67_ASAP7_75t_R clkload41 (.A(clknet_leaf_15_clk_regs));
 BUFx12_ASAP7_75t_R clkload42 (.A(clknet_leaf_16_clk_regs));
 BUFx24_ASAP7_75t_R clkload43 (.A(clknet_leaf_17_clk_regs));
 BUFx4f_ASAP7_75t_R clkload44 (.A(clknet_leaf_18_clk_regs));
 CKINVDCx11_ASAP7_75t_R clkload45 (.A(clknet_leaf_19_clk_regs));
 BUFx4f_ASAP7_75t_R clkload46 (.A(clknet_leaf_20_clk_regs));
 CKINVDCx6p67_ASAP7_75t_R clkload47 (.A(clknet_leaf_21_clk_regs));
 INVx3_ASAP7_75t_R clkload48 (.A(clknet_leaf_22_clk_regs));
 INVx6_ASAP7_75t_R clkload49 (.A(clknet_leaf_23_clk_regs));
 CKINVDCx11_ASAP7_75t_R clkload50 (.A(clknet_leaf_25_clk_regs));
 DECAPx10_ASAP7_75t_R FILLER_0_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_675 ();
 DECAPx6_ASAP7_75t_R FILLER_0_697 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711 ();
 DECAPx1_ASAP7_75t_R FILLER_0_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_745 ();
 DECAPx1_ASAP7_75t_R FILLER_0_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_764 ();
 FILLER_ASAP7_75t_R FILLER_0_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_775 ();
 DECAPx4_ASAP7_75t_R FILLER_0_799 ();
 FILLER_ASAP7_75t_R FILLER_0_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_847 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851 ();
 DECAPx10_ASAP7_75t_R FILLER_0_873 ();
 DECAPx10_ASAP7_75t_R FILLER_0_895 ();
 DECAPx10_ASAP7_75t_R FILLER_0_917 ();
 DECAPx1_ASAP7_75t_R FILLER_0_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_943 ();
 DECAPx10_ASAP7_75t_R FILLER_0_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_971 ();
 DECAPx10_ASAP7_75t_R FILLER_0_974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_546 ();
 DECAPx2_ASAP7_75t_R FILLER_1_586 ();
 FILLER_ASAP7_75t_R FILLER_1_613 ();
 DECAPx1_ASAP7_75t_R FILLER_1_636 ();
 DECAPx1_ASAP7_75t_R FILLER_1_646 ();
 DECAPx2_ASAP7_75t_R FILLER_1_678 ();
 FILLER_ASAP7_75t_R FILLER_1_684 ();
 DECAPx10_ASAP7_75t_R FILLER_1_707 ();
 FILLER_ASAP7_75t_R FILLER_1_729 ();
 FILLER_ASAP7_75t_R FILLER_1_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_740 ();
 FILLER_ASAP7_75t_R FILLER_1_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_764 ();
 FILLER_ASAP7_75t_R FILLER_1_793 ();
 FILLER_ASAP7_75t_R FILLER_1_837 ();
 DECAPx2_ASAP7_75t_R FILLER_1_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_866 ();
 DECAPx6_ASAP7_75t_R FILLER_1_874 ();
 FILLER_ASAP7_75t_R FILLER_1_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_890 ();
 DECAPx2_ASAP7_75t_R FILLER_1_898 ();
 FILLER_ASAP7_75t_R FILLER_1_904 ();
 DECAPx4_ASAP7_75t_R FILLER_1_934 ();
 FILLER_ASAP7_75t_R FILLER_1_944 ();
 DECAPx4_ASAP7_75t_R FILLER_1_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_977 ();
 DECAPx10_ASAP7_75t_R FILLER_1_984 ();
 DECAPx4_ASAP7_75t_R FILLER_1_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_1_1038 ();
 FILLER_ASAP7_75t_R FILLER_1_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1058 ();
 FILLER_ASAP7_75t_R FILLER_1_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1066 ();
 FILLER_ASAP7_75t_R FILLER_1_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1229 ();
 DECAPx4_ASAP7_75t_R FILLER_1_1251 ();
 FILLER_ASAP7_75t_R FILLER_1_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1269 ();
 FILLER_ASAP7_75t_R FILLER_1_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_537 ();
 DECAPx2_ASAP7_75t_R FILLER_2_586 ();
 FILLER_ASAP7_75t_R FILLER_2_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_601 ();
 DECAPx2_ASAP7_75t_R FILLER_2_608 ();
 DECAPx2_ASAP7_75t_R FILLER_2_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_633 ();
 DECAPx6_ASAP7_75t_R FILLER_2_641 ();
 FILLER_ASAP7_75t_R FILLER_2_655 ();
 DECAPx2_ASAP7_75t_R FILLER_2_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_666 ();
 DECAPx6_ASAP7_75t_R FILLER_2_701 ();
 DECAPx2_ASAP7_75t_R FILLER_2_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_742 ();
 DECAPx4_ASAP7_75t_R FILLER_2_756 ();
 FILLER_ASAP7_75t_R FILLER_2_766 ();
 FILLER_ASAP7_75t_R FILLER_2_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_783 ();
 FILLER_ASAP7_75t_R FILLER_2_805 ();
 DECAPx4_ASAP7_75t_R FILLER_2_814 ();
 FILLER_ASAP7_75t_R FILLER_2_824 ();
 DECAPx6_ASAP7_75t_R FILLER_2_833 ();
 DECAPx2_ASAP7_75t_R FILLER_2_854 ();
 FILLER_ASAP7_75t_R FILLER_2_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_862 ();
 DECAPx2_ASAP7_75t_R FILLER_2_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_952 ();
 DECAPx2_ASAP7_75t_R FILLER_2_959 ();
 DECAPx1_ASAP7_75t_R FILLER_2_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_978 ();
 FILLER_ASAP7_75t_R FILLER_2_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_2_1074 ();
 FILLER_ASAP7_75t_R FILLER_2_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_2_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1287 ();
 DECAPx1_ASAP7_75t_R FILLER_3_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_569 ();
 DECAPx10_ASAP7_75t_R FILLER_3_585 ();
 DECAPx10_ASAP7_75t_R FILLER_3_607 ();
 DECAPx6_ASAP7_75t_R FILLER_3_657 ();
 DECAPx2_ASAP7_75t_R FILLER_3_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_677 ();
 DECAPx10_ASAP7_75t_R FILLER_3_684 ();
 DECAPx10_ASAP7_75t_R FILLER_3_706 ();
 DECAPx1_ASAP7_75t_R FILLER_3_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_732 ();
 DECAPx6_ASAP7_75t_R FILLER_3_739 ();
 FILLER_ASAP7_75t_R FILLER_3_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_755 ();
 DECAPx10_ASAP7_75t_R FILLER_3_763 ();
 DECAPx2_ASAP7_75t_R FILLER_3_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_791 ();
 DECAPx4_ASAP7_75t_R FILLER_3_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_808 ();
 DECAPx6_ASAP7_75t_R FILLER_3_815 ();
 FILLER_ASAP7_75t_R FILLER_3_829 ();
 DECAPx2_ASAP7_75t_R FILLER_3_837 ();
 FILLER_ASAP7_75t_R FILLER_3_843 ();
 DECAPx2_ASAP7_75t_R FILLER_3_866 ();
 DECAPx6_ASAP7_75t_R FILLER_3_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_892 ();
 DECAPx1_ASAP7_75t_R FILLER_3_899 ();
 DECAPx1_ASAP7_75t_R FILLER_3_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_913 ();
 FILLER_ASAP7_75t_R FILLER_3_921 ();
 DECAPx6_ASAP7_75t_R FILLER_3_950 ();
 FILLER_ASAP7_75t_R FILLER_3_985 ();
 DECAPx4_ASAP7_75t_R FILLER_3_993 ();
 FILLER_ASAP7_75t_R FILLER_3_1003 ();
 FILLER_ASAP7_75t_R FILLER_3_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_4_580 ();
 DECAPx10_ASAP7_75t_R FILLER_4_620 ();
 DECAPx2_ASAP7_75t_R FILLER_4_642 ();
 FILLER_ASAP7_75t_R FILLER_4_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_671 ();
 DECAPx10_ASAP7_75t_R FILLER_4_679 ();
 DECAPx10_ASAP7_75t_R FILLER_4_701 ();
 DECAPx10_ASAP7_75t_R FILLER_4_723 ();
 DECAPx2_ASAP7_75t_R FILLER_4_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_751 ();
 DECAPx4_ASAP7_75t_R FILLER_4_773 ();
 FILLER_ASAP7_75t_R FILLER_4_783 ();
 DECAPx10_ASAP7_75t_R FILLER_4_788 ();
 DECAPx4_ASAP7_75t_R FILLER_4_810 ();
 FILLER_ASAP7_75t_R FILLER_4_820 ();
 DECAPx6_ASAP7_75t_R FILLER_4_832 ();
 DECAPx2_ASAP7_75t_R FILLER_4_846 ();
 DECAPx10_ASAP7_75t_R FILLER_4_858 ();
 DECAPx10_ASAP7_75t_R FILLER_4_880 ();
 DECAPx10_ASAP7_75t_R FILLER_4_902 ();
 DECAPx10_ASAP7_75t_R FILLER_4_924 ();
 DECAPx10_ASAP7_75t_R FILLER_4_946 ();
 DECAPx1_ASAP7_75t_R FILLER_4_968 ();
 DECAPx10_ASAP7_75t_R FILLER_4_974 ();
 DECAPx6_ASAP7_75t_R FILLER_4_996 ();
 FILLER_ASAP7_75t_R FILLER_4_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_4_1281 ();
 FILLER_ASAP7_75t_R FILLER_4_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_5_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_587 ();
 DECAPx6_ASAP7_75t_R FILLER_5_637 ();
 DECAPx1_ASAP7_75t_R FILLER_5_651 ();
 DECAPx2_ASAP7_75t_R FILLER_5_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_667 ();
 DECAPx2_ASAP7_75t_R FILLER_5_731 ();
 FILLER_ASAP7_75t_R FILLER_5_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_739 ();
 FILLER_ASAP7_75t_R FILLER_5_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_769 ();
 DECAPx10_ASAP7_75t_R FILLER_5_783 ();
 DECAPx2_ASAP7_75t_R FILLER_5_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_811 ();
 DECAPx10_ASAP7_75t_R FILLER_5_839 ();
 DECAPx4_ASAP7_75t_R FILLER_5_861 ();
 FILLER_ASAP7_75t_R FILLER_5_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_873 ();
 DECAPx6_ASAP7_75t_R FILLER_5_895 ();
 DECAPx2_ASAP7_75t_R FILLER_5_909 ();
 DECAPx6_ASAP7_75t_R FILLER_5_922 ();
 DECAPx1_ASAP7_75t_R FILLER_5_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_940 ();
 DECAPx6_ASAP7_75t_R FILLER_5_948 ();
 DECAPx10_ASAP7_75t_R FILLER_5_983 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_5_1281 ();
 FILLER_ASAP7_75t_R FILLER_5_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_6_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_566 ();
 DECAPx6_ASAP7_75t_R FILLER_6_572 ();
 FILLER_ASAP7_75t_R FILLER_6_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_588 ();
 DECAPx6_ASAP7_75t_R FILLER_6_596 ();
 FILLER_ASAP7_75t_R FILLER_6_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_634 ();
 DECAPx6_ASAP7_75t_R FILLER_6_656 ();
 DECAPx1_ASAP7_75t_R FILLER_6_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_674 ();
 DECAPx2_ASAP7_75t_R FILLER_6_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_687 ();
 DECAPx6_ASAP7_75t_R FILLER_6_701 ();
 FILLER_ASAP7_75t_R FILLER_6_715 ();
 DECAPx4_ASAP7_75t_R FILLER_6_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_740 ();
 FILLER_ASAP7_75t_R FILLER_6_756 ();
 FILLER_ASAP7_75t_R FILLER_6_765 ();
 DECAPx4_ASAP7_75t_R FILLER_6_794 ();
 FILLER_ASAP7_75t_R FILLER_6_804 ();
 DECAPx10_ASAP7_75t_R FILLER_6_827 ();
 FILLER_ASAP7_75t_R FILLER_6_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_851 ();
 DECAPx1_ASAP7_75t_R FILLER_6_886 ();
 DECAPx1_ASAP7_75t_R FILLER_6_911 ();
 DECAPx6_ASAP7_75t_R FILLER_6_948 ();
 FILLER_ASAP7_75t_R FILLER_6_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_980 ();
 DECAPx1_ASAP7_75t_R FILLER_6_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_998 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1055 ();
 FILLER_ASAP7_75t_R FILLER_6_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_7_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_546 ();
 DECAPx2_ASAP7_75t_R FILLER_7_562 ();
 FILLER_ASAP7_75t_R FILLER_7_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_570 ();
 DECAPx2_ASAP7_75t_R FILLER_7_578 ();
 FILLER_ASAP7_75t_R FILLER_7_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_586 ();
 DECAPx6_ASAP7_75t_R FILLER_7_608 ();
 DECAPx2_ASAP7_75t_R FILLER_7_622 ();
 DECAPx10_ASAP7_75t_R FILLER_7_658 ();
 DECAPx10_ASAP7_75t_R FILLER_7_680 ();
 DECAPx6_ASAP7_75t_R FILLER_7_702 ();
 DECAPx1_ASAP7_75t_R FILLER_7_716 ();
 DECAPx10_ASAP7_75t_R FILLER_7_771 ();
 DECAPx10_ASAP7_75t_R FILLER_7_793 ();
 DECAPx6_ASAP7_75t_R FILLER_7_815 ();
 FILLER_ASAP7_75t_R FILLER_7_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_831 ();
 DECAPx6_ASAP7_75t_R FILLER_7_839 ();
 FILLER_ASAP7_75t_R FILLER_7_853 ();
 DECAPx2_ASAP7_75t_R FILLER_7_868 ();
 FILLER_ASAP7_75t_R FILLER_7_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_876 ();
 DECAPx6_ASAP7_75t_R FILLER_7_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_904 ();
 FILLER_ASAP7_75t_R FILLER_7_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_920 ();
 DECAPx2_ASAP7_75t_R FILLER_7_927 ();
 FILLER_ASAP7_75t_R FILLER_7_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_942 ();
 DECAPx6_ASAP7_75t_R FILLER_7_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_978 ();
 DECAPx1_ASAP7_75t_R FILLER_7_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_7_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_7_1042 ();
 FILLER_ASAP7_75t_R FILLER_7_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1058 ();
 FILLER_ASAP7_75t_R FILLER_7_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1077 ();
 FILLER_ASAP7_75t_R FILLER_7_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_7_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_8_552 ();
 FILLER_ASAP7_75t_R FILLER_8_566 ();
 DECAPx1_ASAP7_75t_R FILLER_8_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_599 ();
 DECAPx2_ASAP7_75t_R FILLER_8_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_612 ();
 FILLER_ASAP7_75t_R FILLER_8_626 ();
 DECAPx2_ASAP7_75t_R FILLER_8_635 ();
 FILLER_ASAP7_75t_R FILLER_8_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_643 ();
 DECAPx10_ASAP7_75t_R FILLER_8_650 ();
 DECAPx1_ASAP7_75t_R FILLER_8_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_676 ();
 DECAPx10_ASAP7_75t_R FILLER_8_683 ();
 DECAPx2_ASAP7_75t_R FILLER_8_705 ();
 FILLER_ASAP7_75t_R FILLER_8_711 ();
 DECAPx4_ASAP7_75t_R FILLER_8_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_747 ();
 FILLER_ASAP7_75t_R FILLER_8_769 ();
 DECAPx2_ASAP7_75t_R FILLER_8_778 ();
 FILLER_ASAP7_75t_R FILLER_8_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_820 ();
 FILLER_ASAP7_75t_R FILLER_8_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_851 ();
 DECAPx6_ASAP7_75t_R FILLER_8_859 ();
 DECAPx1_ASAP7_75t_R FILLER_8_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_877 ();
 DECAPx10_ASAP7_75t_R FILLER_8_899 ();
 DECAPx4_ASAP7_75t_R FILLER_8_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_931 ();
 DECAPx6_ASAP7_75t_R FILLER_8_953 ();
 DECAPx1_ASAP7_75t_R FILLER_8_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_971 ();
 FILLER_ASAP7_75t_R FILLER_8_974 ();
 DECAPx6_ASAP7_75t_R FILLER_8_997 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1029 ();
 FILLER_ASAP7_75t_R FILLER_8_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_9_537 ();
 DECAPx10_ASAP7_75t_R FILLER_9_559 ();
 DECAPx10_ASAP7_75t_R FILLER_9_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_603 ();
 DECAPx10_ASAP7_75t_R FILLER_9_611 ();
 DECAPx10_ASAP7_75t_R FILLER_9_633 ();
 DECAPx1_ASAP7_75t_R FILLER_9_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_708 ();
 FILLER_ASAP7_75t_R FILLER_9_715 ();
 DECAPx1_ASAP7_75t_R FILLER_9_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_728 ();
 DECAPx10_ASAP7_75t_R FILLER_9_735 ();
 DECAPx1_ASAP7_75t_R FILLER_9_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_768 ();
 DECAPx10_ASAP7_75t_R FILLER_9_803 ();
 DECAPx2_ASAP7_75t_R FILLER_9_825 ();
 FILLER_ASAP7_75t_R FILLER_9_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_833 ();
 DECAPx4_ASAP7_75t_R FILLER_9_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_850 ();
 DECAPx10_ASAP7_75t_R FILLER_9_881 ();
 DECAPx1_ASAP7_75t_R FILLER_9_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_907 ();
 DECAPx10_ASAP7_75t_R FILLER_9_915 ();
 DECAPx10_ASAP7_75t_R FILLER_9_937 ();
 DECAPx1_ASAP7_75t_R FILLER_9_959 ();
 FILLER_ASAP7_75t_R FILLER_9_973 ();
 DECAPx2_ASAP7_75t_R FILLER_9_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_994 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_9_1024 ();
 FILLER_ASAP7_75t_R FILLER_9_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_9_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_10_532 ();
 DECAPx1_ASAP7_75t_R FILLER_10_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_558 ();
 DECAPx10_ASAP7_75t_R FILLER_10_569 ();
 DECAPx4_ASAP7_75t_R FILLER_10_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_601 ();
 DECAPx4_ASAP7_75t_R FILLER_10_629 ();
 DECAPx4_ASAP7_75t_R FILLER_10_686 ();
 FILLER_ASAP7_75t_R FILLER_10_696 ();
 DECAPx10_ASAP7_75t_R FILLER_10_705 ();
 DECAPx2_ASAP7_75t_R FILLER_10_727 ();
 FILLER_ASAP7_75t_R FILLER_10_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_735 ();
 DECAPx10_ASAP7_75t_R FILLER_10_764 ();
 DECAPx10_ASAP7_75t_R FILLER_10_786 ();
 DECAPx4_ASAP7_75t_R FILLER_10_836 ();
 FILLER_ASAP7_75t_R FILLER_10_846 ();
 DECAPx10_ASAP7_75t_R FILLER_10_869 ();
 DECAPx4_ASAP7_75t_R FILLER_10_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_901 ();
 DECAPx6_ASAP7_75t_R FILLER_10_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_937 ();
 DECAPx2_ASAP7_75t_R FILLER_10_966 ();
 DECAPx6_ASAP7_75t_R FILLER_10_974 ();
 DECAPx2_ASAP7_75t_R FILLER_10_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1022 ();
 FILLER_ASAP7_75t_R FILLER_10_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_10_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_11_527 ();
 DECAPx10_ASAP7_75t_R FILLER_11_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_571 ();
 DECAPx10_ASAP7_75t_R FILLER_11_582 ();
 DECAPx4_ASAP7_75t_R FILLER_11_604 ();
 FILLER_ASAP7_75t_R FILLER_11_614 ();
 FILLER_ASAP7_75t_R FILLER_11_624 ();
 DECAPx1_ASAP7_75t_R FILLER_11_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_637 ();
 DECAPx6_ASAP7_75t_R FILLER_11_659 ();
 FILLER_ASAP7_75t_R FILLER_11_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_675 ();
 FILLER_ASAP7_75t_R FILLER_11_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_686 ();
 DECAPx10_ASAP7_75t_R FILLER_11_694 ();
 DECAPx10_ASAP7_75t_R FILLER_11_716 ();
 DECAPx1_ASAP7_75t_R FILLER_11_738 ();
 DECAPx6_ASAP7_75t_R FILLER_11_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_762 ();
 DECAPx6_ASAP7_75t_R FILLER_11_771 ();
 DECAPx6_ASAP7_75t_R FILLER_11_792 ();
 DECAPx1_ASAP7_75t_R FILLER_11_806 ();
 DECAPx1_ASAP7_75t_R FILLER_11_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_820 ();
 DECAPx10_ASAP7_75t_R FILLER_11_828 ();
 DECAPx4_ASAP7_75t_R FILLER_11_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_867 ();
 DECAPx10_ASAP7_75t_R FILLER_11_875 ();
 DECAPx6_ASAP7_75t_R FILLER_11_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_911 ();
 DECAPx10_ASAP7_75t_R FILLER_11_952 ();
 DECAPx10_ASAP7_75t_R FILLER_11_974 ();
 DECAPx4_ASAP7_75t_R FILLER_11_1002 ();
 FILLER_ASAP7_75t_R FILLER_11_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_11_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_11_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_11_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1285 ();
 FILLER_ASAP7_75t_R FILLER_11_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_12_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_519 ();
 DECAPx10_ASAP7_75t_R FILLER_12_523 ();
 DECAPx2_ASAP7_75t_R FILLER_12_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_551 ();
 DECAPx4_ASAP7_75t_R FILLER_12_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_593 ();
 DECAPx6_ASAP7_75t_R FILLER_12_604 ();
 FILLER_ASAP7_75t_R FILLER_12_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_620 ();
 DECAPx10_ASAP7_75t_R FILLER_12_648 ();
 DECAPx2_ASAP7_75t_R FILLER_12_670 ();
 DECAPx6_ASAP7_75t_R FILLER_12_703 ();
 FILLER_ASAP7_75t_R FILLER_12_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_719 ();
 DECAPx4_ASAP7_75t_R FILLER_12_730 ();
 DECAPx6_ASAP7_75t_R FILLER_12_803 ();
 FILLER_ASAP7_75t_R FILLER_12_817 ();
 DECAPx10_ASAP7_75t_R FILLER_12_840 ();
 DECAPx2_ASAP7_75t_R FILLER_12_862 ();
 FILLER_ASAP7_75t_R FILLER_12_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_870 ();
 DECAPx4_ASAP7_75t_R FILLER_12_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_887 ();
 DECAPx2_ASAP7_75t_R FILLER_12_901 ();
 FILLER_ASAP7_75t_R FILLER_12_907 ();
 DECAPx10_ASAP7_75t_R FILLER_12_936 ();
 DECAPx2_ASAP7_75t_R FILLER_12_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_964 ();
 DECAPx10_ASAP7_75t_R FILLER_12_980 ();
 DECAPx4_ASAP7_75t_R FILLER_12_1002 ();
 FILLER_ASAP7_75t_R FILLER_12_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_12_1050 ();
 FILLER_ASAP7_75t_R FILLER_12_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_12_1073 ();
 FILLER_ASAP7_75t_R FILLER_12_1087 ();
 FILLER_ASAP7_75t_R FILLER_12_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_12_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_13_518 ();
 DECAPx4_ASAP7_75t_R FILLER_13_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_550 ();
 FILLER_ASAP7_75t_R FILLER_13_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_574 ();
 DECAPx6_ASAP7_75t_R FILLER_13_582 ();
 DECAPx2_ASAP7_75t_R FILLER_13_596 ();
 DECAPx10_ASAP7_75t_R FILLER_13_612 ();
 DECAPx4_ASAP7_75t_R FILLER_13_634 ();
 DECAPx6_ASAP7_75t_R FILLER_13_668 ();
 FILLER_ASAP7_75t_R FILLER_13_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_684 ();
 DECAPx10_ASAP7_75t_R FILLER_13_693 ();
 DECAPx10_ASAP7_75t_R FILLER_13_715 ();
 DECAPx2_ASAP7_75t_R FILLER_13_737 ();
 DECAPx2_ASAP7_75t_R FILLER_13_750 ();
 DECAPx6_ASAP7_75t_R FILLER_13_759 ();
 FILLER_ASAP7_75t_R FILLER_13_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_775 ();
 DECAPx2_ASAP7_75t_R FILLER_13_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_789 ();
 DECAPx2_ASAP7_75t_R FILLER_13_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_802 ();
 DECAPx4_ASAP7_75t_R FILLER_13_831 ();
 FILLER_ASAP7_75t_R FILLER_13_841 ();
 DECAPx6_ASAP7_75t_R FILLER_13_916 ();
 DECAPx2_ASAP7_75t_R FILLER_13_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_936 ();
 FILLER_ASAP7_75t_R FILLER_13_944 ();
 DECAPx2_ASAP7_75t_R FILLER_13_997 ();
 FILLER_ASAP7_75t_R FILLER_13_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_13_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_13_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_14_512 ();
 DECAPx1_ASAP7_75t_R FILLER_14_534 ();
 DECAPx4_ASAP7_75t_R FILLER_14_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_556 ();
 DECAPx1_ASAP7_75t_R FILLER_14_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_574 ();
 DECAPx4_ASAP7_75t_R FILLER_14_581 ();
 DECAPx4_ASAP7_75t_R FILLER_14_600 ();
 FILLER_ASAP7_75t_R FILLER_14_610 ();
 FILLER_ASAP7_75t_R FILLER_14_619 ();
 DECAPx10_ASAP7_75t_R FILLER_14_627 ();
 DECAPx10_ASAP7_75t_R FILLER_14_649 ();
 DECAPx10_ASAP7_75t_R FILLER_14_671 ();
 DECAPx2_ASAP7_75t_R FILLER_14_693 ();
 FILLER_ASAP7_75t_R FILLER_14_699 ();
 DECAPx10_ASAP7_75t_R FILLER_14_726 ();
 DECAPx2_ASAP7_75t_R FILLER_14_748 ();
 DECAPx6_ASAP7_75t_R FILLER_14_760 ();
 DECAPx6_ASAP7_75t_R FILLER_14_780 ();
 DECAPx2_ASAP7_75t_R FILLER_14_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_800 ();
 DECAPx2_ASAP7_75t_R FILLER_14_814 ();
 FILLER_ASAP7_75t_R FILLER_14_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_822 ();
 DECAPx10_ASAP7_75t_R FILLER_14_826 ();
 DECAPx10_ASAP7_75t_R FILLER_14_848 ();
 DECAPx10_ASAP7_75t_R FILLER_14_870 ();
 DECAPx10_ASAP7_75t_R FILLER_14_892 ();
 DECAPx10_ASAP7_75t_R FILLER_14_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_936 ();
 DECAPx6_ASAP7_75t_R FILLER_14_958 ();
 DECAPx1_ASAP7_75t_R FILLER_14_974 ();
 DECAPx2_ASAP7_75t_R FILLER_14_985 ();
 FILLER_ASAP7_75t_R FILLER_14_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1040 ();
 FILLER_ASAP7_75t_R FILLER_14_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_14_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1281 ();
 FILLER_ASAP7_75t_R FILLER_14_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_15_512 ();
 DECAPx1_ASAP7_75t_R FILLER_15_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_530 ();
 DECAPx4_ASAP7_75t_R FILLER_15_541 ();
 DECAPx10_ASAP7_75t_R FILLER_15_564 ();
 DECAPx1_ASAP7_75t_R FILLER_15_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_593 ();
 DECAPx10_ASAP7_75t_R FILLER_15_636 ();
 DECAPx10_ASAP7_75t_R FILLER_15_658 ();
 DECAPx6_ASAP7_75t_R FILLER_15_680 ();
 FILLER_ASAP7_75t_R FILLER_15_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_696 ();
 DECAPx10_ASAP7_75t_R FILLER_15_723 ();
 DECAPx2_ASAP7_75t_R FILLER_15_755 ();
 FILLER_ASAP7_75t_R FILLER_15_761 ();
 DECAPx1_ASAP7_75t_R FILLER_15_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_774 ();
 DECAPx10_ASAP7_75t_R FILLER_15_778 ();
 DECAPx10_ASAP7_75t_R FILLER_15_800 ();
 DECAPx2_ASAP7_75t_R FILLER_15_822 ();
 FILLER_ASAP7_75t_R FILLER_15_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_830 ();
 DECAPx6_ASAP7_75t_R FILLER_15_837 ();
 FILLER_ASAP7_75t_R FILLER_15_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_853 ();
 DECAPx10_ASAP7_75t_R FILLER_15_876 ();
 FILLER_ASAP7_75t_R FILLER_15_898 ();
 DECAPx4_ASAP7_75t_R FILLER_15_907 ();
 FILLER_ASAP7_75t_R FILLER_15_917 ();
 DECAPx10_ASAP7_75t_R FILLER_15_948 ();
 FILLER_ASAP7_75t_R FILLER_15_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_972 ();
 DECAPx6_ASAP7_75t_R FILLER_15_994 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_15_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1086 ();
 FILLER_ASAP7_75t_R FILLER_15_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1098 ();
 DECAPx4_ASAP7_75t_R FILLER_15_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_15_1281 ();
 FILLER_ASAP7_75t_R FILLER_15_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_16_512 ();
 DECAPx2_ASAP7_75t_R FILLER_16_534 ();
 DECAPx4_ASAP7_75t_R FILLER_16_561 ();
 DECAPx10_ASAP7_75t_R FILLER_16_584 ();
 DECAPx10_ASAP7_75t_R FILLER_16_606 ();
 DECAPx10_ASAP7_75t_R FILLER_16_628 ();
 DECAPx6_ASAP7_75t_R FILLER_16_656 ();
 FILLER_ASAP7_75t_R FILLER_16_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_709 ();
 DECAPx4_ASAP7_75t_R FILLER_16_736 ();
 FILLER_ASAP7_75t_R FILLER_16_746 ();
 DECAPx6_ASAP7_75t_R FILLER_16_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_789 ();
 DECAPx4_ASAP7_75t_R FILLER_16_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_814 ();
 FILLER_ASAP7_75t_R FILLER_16_830 ();
 DECAPx2_ASAP7_75t_R FILLER_16_840 ();
 FILLER_ASAP7_75t_R FILLER_16_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_848 ();
 FILLER_ASAP7_75t_R FILLER_16_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_873 ();
 DECAPx1_ASAP7_75t_R FILLER_16_880 ();
 FILLER_ASAP7_75t_R FILLER_16_896 ();
 DECAPx4_ASAP7_75t_R FILLER_16_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_945 ();
 DECAPx6_ASAP7_75t_R FILLER_16_953 ();
 DECAPx1_ASAP7_75t_R FILLER_16_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_971 ();
 DECAPx10_ASAP7_75t_R FILLER_16_974 ();
 DECAPx2_ASAP7_75t_R FILLER_16_996 ();
 FILLER_ASAP7_75t_R FILLER_16_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1110 ();
 DECAPx4_ASAP7_75t_R FILLER_16_1132 ();
 FILLER_ASAP7_75t_R FILLER_16_1142 ();
 FILLER_ASAP7_75t_R FILLER_16_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_16_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_17_518 ();
 DECAPx10_ASAP7_75t_R FILLER_17_540 ();
 DECAPx2_ASAP7_75t_R FILLER_17_562 ();
 FILLER_ASAP7_75t_R FILLER_17_568 ();
 DECAPx10_ASAP7_75t_R FILLER_17_597 ();
 DECAPx6_ASAP7_75t_R FILLER_17_619 ();
 FILLER_ASAP7_75t_R FILLER_17_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_635 ();
 DECAPx1_ASAP7_75t_R FILLER_17_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_654 ();
 DECAPx1_ASAP7_75t_R FILLER_17_682 ();
 DECAPx1_ASAP7_75t_R FILLER_17_704 ();
 DECAPx10_ASAP7_75t_R FILLER_17_714 ();
 DECAPx1_ASAP7_75t_R FILLER_17_736 ();
 DECAPx4_ASAP7_75t_R FILLER_17_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_773 ();
 FILLER_ASAP7_75t_R FILLER_17_780 ();
 DECAPx1_ASAP7_75t_R FILLER_17_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_798 ();
 DECAPx4_ASAP7_75t_R FILLER_17_813 ();
 DECAPx10_ASAP7_75t_R FILLER_17_830 ();
 DECAPx4_ASAP7_75t_R FILLER_17_852 ();
 FILLER_ASAP7_75t_R FILLER_17_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_864 ();
 DECAPx1_ASAP7_75t_R FILLER_17_873 ();
 FILLER_ASAP7_75t_R FILLER_17_887 ();
 DECAPx2_ASAP7_75t_R FILLER_17_895 ();
 FILLER_ASAP7_75t_R FILLER_17_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_903 ();
 DECAPx10_ASAP7_75t_R FILLER_17_910 ();
 DECAPx2_ASAP7_75t_R FILLER_17_932 ();
 FILLER_ASAP7_75t_R FILLER_17_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_940 ();
 DECAPx10_ASAP7_75t_R FILLER_17_983 ();
 FILLER_ASAP7_75t_R FILLER_17_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1059 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_17_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1105 ();
 FILLER_ASAP7_75t_R FILLER_17_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_17_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_18_518 ();
 DECAPx10_ASAP7_75t_R FILLER_18_540 ();
 DECAPx1_ASAP7_75t_R FILLER_18_562 ();
 DECAPx2_ASAP7_75t_R FILLER_18_574 ();
 DECAPx10_ASAP7_75t_R FILLER_18_590 ();
 DECAPx4_ASAP7_75t_R FILLER_18_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_622 ();
 DECAPx4_ASAP7_75t_R FILLER_18_648 ();
 FILLER_ASAP7_75t_R FILLER_18_658 ();
 DECAPx2_ASAP7_75t_R FILLER_18_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_674 ();
 DECAPx10_ASAP7_75t_R FILLER_18_681 ();
 DECAPx2_ASAP7_75t_R FILLER_18_703 ();
 FILLER_ASAP7_75t_R FILLER_18_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_711 ();
 DECAPx6_ASAP7_75t_R FILLER_18_724 ();
 DECAPx1_ASAP7_75t_R FILLER_18_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_742 ();
 DECAPx6_ASAP7_75t_R FILLER_18_751 ();
 DECAPx1_ASAP7_75t_R FILLER_18_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_783 ();
 DECAPx6_ASAP7_75t_R FILLER_18_792 ();
 DECAPx2_ASAP7_75t_R FILLER_18_812 ();
 FILLER_ASAP7_75t_R FILLER_18_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_834 ();
 FILLER_ASAP7_75t_R FILLER_18_838 ();
 DECAPx2_ASAP7_75t_R FILLER_18_848 ();
 FILLER_ASAP7_75t_R FILLER_18_854 ();
 DECAPx10_ASAP7_75t_R FILLER_18_864 ();
 DECAPx10_ASAP7_75t_R FILLER_18_886 ();
 DECAPx10_ASAP7_75t_R FILLER_18_908 ();
 DECAPx6_ASAP7_75t_R FILLER_18_930 ();
 DECAPx2_ASAP7_75t_R FILLER_18_944 ();
 DECAPx2_ASAP7_75t_R FILLER_18_956 ();
 FILLER_ASAP7_75t_R FILLER_18_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_971 ();
 DECAPx6_ASAP7_75t_R FILLER_18_974 ();
 FILLER_ASAP7_75t_R FILLER_18_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_990 ();
 DECAPx4_ASAP7_75t_R FILLER_18_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_18_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1137 ();
 FILLER_ASAP7_75t_R FILLER_18_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_19_512 ();
 FILLER_ASAP7_75t_R FILLER_19_522 ();
 DECAPx6_ASAP7_75t_R FILLER_19_540 ();
 DECAPx2_ASAP7_75t_R FILLER_19_582 ();
 DECAPx10_ASAP7_75t_R FILLER_19_603 ();
 DECAPx1_ASAP7_75t_R FILLER_19_625 ();
 DECAPx6_ASAP7_75t_R FILLER_19_647 ();
 DECAPx6_ASAP7_75t_R FILLER_19_681 ();
 FILLER_ASAP7_75t_R FILLER_19_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_708 ();
 DECAPx10_ASAP7_75t_R FILLER_19_721 ();
 DECAPx6_ASAP7_75t_R FILLER_19_743 ();
 DECAPx1_ASAP7_75t_R FILLER_19_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_761 ();
 DECAPx10_ASAP7_75t_R FILLER_19_768 ();
 DECAPx4_ASAP7_75t_R FILLER_19_790 ();
 DECAPx1_ASAP7_75t_R FILLER_19_808 ();
 DECAPx10_ASAP7_75t_R FILLER_19_838 ();
 DECAPx2_ASAP7_75t_R FILLER_19_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_872 ();
 DECAPx6_ASAP7_75t_R FILLER_19_895 ();
 DECAPx2_ASAP7_75t_R FILLER_19_930 ();
 DECAPx2_ASAP7_75t_R FILLER_19_942 ();
 FILLER_ASAP7_75t_R FILLER_19_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_950 ();
 DECAPx2_ASAP7_75t_R FILLER_19_954 ();
 FILLER_ASAP7_75t_R FILLER_19_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_962 ();
 FILLER_ASAP7_75t_R FILLER_19_969 ();
 DECAPx10_ASAP7_75t_R FILLER_19_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1031 ();
 FILLER_ASAP7_75t_R FILLER_19_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1096 ();
 FILLER_ASAP7_75t_R FILLER_19_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_19_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_19_1171 ();
 FILLER_ASAP7_75t_R FILLER_19_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1183 ();
 FILLER_ASAP7_75t_R FILLER_19_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_20_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_547 ();
 DECAPx6_ASAP7_75t_R FILLER_20_576 ();
 FILLER_ASAP7_75t_R FILLER_20_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_592 ();
 DECAPx10_ASAP7_75t_R FILLER_20_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_639 ();
 DECAPx1_ASAP7_75t_R FILLER_20_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_662 ();
 DECAPx2_ASAP7_75t_R FILLER_20_669 ();
 FILLER_ASAP7_75t_R FILLER_20_675 ();
 DECAPx6_ASAP7_75t_R FILLER_20_693 ();
 DECAPx2_ASAP7_75t_R FILLER_20_707 ();
 DECAPx4_ASAP7_75t_R FILLER_20_722 ();
 FILLER_ASAP7_75t_R FILLER_20_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_734 ();
 DECAPx2_ASAP7_75t_R FILLER_20_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_763 ();
 DECAPx10_ASAP7_75t_R FILLER_20_770 ();
 DECAPx10_ASAP7_75t_R FILLER_20_792 ();
 DECAPx10_ASAP7_75t_R FILLER_20_814 ();
 DECAPx6_ASAP7_75t_R FILLER_20_836 ();
 DECAPx2_ASAP7_75t_R FILLER_20_850 ();
 DECAPx6_ASAP7_75t_R FILLER_20_871 ();
 FILLER_ASAP7_75t_R FILLER_20_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_887 ();
 DECAPx6_ASAP7_75t_R FILLER_20_898 ();
 FILLER_ASAP7_75t_R FILLER_20_949 ();
 DECAPx10_ASAP7_75t_R FILLER_20_974 ();
 DECAPx6_ASAP7_75t_R FILLER_20_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1010 ();
 FILLER_ASAP7_75t_R FILLER_20_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_20_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_20_1066 ();
 FILLER_ASAP7_75t_R FILLER_20_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1129 ();
 FILLER_ASAP7_75t_R FILLER_20_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_20_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_20_1277 ();
 FILLER_ASAP7_75t_R FILLER_20_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_21_512 ();
 DECAPx1_ASAP7_75t_R FILLER_21_534 ();
 FILLER_ASAP7_75t_R FILLER_21_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_553 ();
 DECAPx10_ASAP7_75t_R FILLER_21_605 ();
 DECAPx10_ASAP7_75t_R FILLER_21_627 ();
 DECAPx10_ASAP7_75t_R FILLER_21_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_671 ();
 DECAPx4_ASAP7_75t_R FILLER_21_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_700 ();
 DECAPx2_ASAP7_75t_R FILLER_21_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_727 ();
 DECAPx4_ASAP7_75t_R FILLER_21_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_764 ();
 DECAPx2_ASAP7_75t_R FILLER_21_774 ();
 FILLER_ASAP7_75t_R FILLER_21_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_782 ();
 FILLER_ASAP7_75t_R FILLER_21_795 ();
 DECAPx6_ASAP7_75t_R FILLER_21_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_825 ();
 DECAPx6_ASAP7_75t_R FILLER_21_834 ();
 DECAPx2_ASAP7_75t_R FILLER_21_848 ();
 DECAPx2_ASAP7_75t_R FILLER_21_864 ();
 FILLER_ASAP7_75t_R FILLER_21_876 ();
 DECAPx1_ASAP7_75t_R FILLER_21_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_890 ();
 DECAPx1_ASAP7_75t_R FILLER_21_905 ();
 DECAPx6_ASAP7_75t_R FILLER_21_923 ();
 FILLER_ASAP7_75t_R FILLER_21_937 ();
 FILLER_ASAP7_75t_R FILLER_21_946 ();
 DECAPx10_ASAP7_75t_R FILLER_21_961 ();
 DECAPx6_ASAP7_75t_R FILLER_21_983 ();
 DECAPx4_ASAP7_75t_R FILLER_21_1003 ();
 FILLER_ASAP7_75t_R FILLER_21_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_21_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_21_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_21_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_21_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_22_512 ();
 DECAPx4_ASAP7_75t_R FILLER_22_534 ();
 FILLER_ASAP7_75t_R FILLER_22_544 ();
 DECAPx1_ASAP7_75t_R FILLER_22_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_578 ();
 DECAPx2_ASAP7_75t_R FILLER_22_586 ();
 DECAPx4_ASAP7_75t_R FILLER_22_598 ();
 DECAPx6_ASAP7_75t_R FILLER_22_629 ();
 DECAPx1_ASAP7_75t_R FILLER_22_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_647 ();
 FILLER_ASAP7_75t_R FILLER_22_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_672 ();
 DECAPx10_ASAP7_75t_R FILLER_22_679 ();
 FILLER_ASAP7_75t_R FILLER_22_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_729 ();
 FILLER_ASAP7_75t_R FILLER_22_739 ();
 FILLER_ASAP7_75t_R FILLER_22_755 ();
 FILLER_ASAP7_75t_R FILLER_22_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_799 ();
 DECAPx2_ASAP7_75t_R FILLER_22_834 ();
 DECAPx4_ASAP7_75t_R FILLER_22_849 ();
 DECAPx2_ASAP7_75t_R FILLER_22_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_895 ();
 FILLER_ASAP7_75t_R FILLER_22_904 ();
 DECAPx10_ASAP7_75t_R FILLER_22_912 ();
 DECAPx4_ASAP7_75t_R FILLER_22_934 ();
 FILLER_ASAP7_75t_R FILLER_22_944 ();
 DECAPx1_ASAP7_75t_R FILLER_22_968 ();
 DECAPx6_ASAP7_75t_R FILLER_22_974 ();
 DECAPx1_ASAP7_75t_R FILLER_22_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_992 ();
 DECAPx6_ASAP7_75t_R FILLER_22_1005 ();
 FILLER_ASAP7_75t_R FILLER_22_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1021 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1040 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1084 ();
 FILLER_ASAP7_75t_R FILLER_22_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_22_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1161 ();
 FILLER_ASAP7_75t_R FILLER_22_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1280 ();
 FILLER_ASAP7_75t_R FILLER_22_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_23_512 ();
 DECAPx6_ASAP7_75t_R FILLER_23_534 ();
 DECAPx1_ASAP7_75t_R FILLER_23_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_552 ();
 FILLER_ASAP7_75t_R FILLER_23_560 ();
 DECAPx1_ASAP7_75t_R FILLER_23_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_593 ();
 DECAPx1_ASAP7_75t_R FILLER_23_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_618 ();
 DECAPx10_ASAP7_75t_R FILLER_23_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_665 ();
 DECAPx6_ASAP7_75t_R FILLER_23_682 ();
 DECAPx4_ASAP7_75t_R FILLER_23_714 ();
 DECAPx10_ASAP7_75t_R FILLER_23_740 ();
 DECAPx10_ASAP7_75t_R FILLER_23_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_798 ();
 DECAPx4_ASAP7_75t_R FILLER_23_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_823 ();
 DECAPx4_ASAP7_75t_R FILLER_23_830 ();
 DECAPx1_ASAP7_75t_R FILLER_23_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_881 ();
 DECAPx2_ASAP7_75t_R FILLER_23_888 ();
 FILLER_ASAP7_75t_R FILLER_23_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_896 ();
 DECAPx1_ASAP7_75t_R FILLER_23_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_907 ();
 DECAPx6_ASAP7_75t_R FILLER_23_916 ();
 FILLER_ASAP7_75t_R FILLER_23_944 ();
 DECAPx10_ASAP7_75t_R FILLER_23_961 ();
 DECAPx4_ASAP7_75t_R FILLER_23_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_993 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1004 ();
 FILLER_ASAP7_75t_R FILLER_23_1026 ();
 FILLER_ASAP7_75t_R FILLER_23_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_23_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1149 ();
 FILLER_ASAP7_75t_R FILLER_23_1159 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_23_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_23_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_24_512 ();
 FILLER_ASAP7_75t_R FILLER_24_518 ();
 DECAPx6_ASAP7_75t_R FILLER_24_557 ();
 DECAPx4_ASAP7_75t_R FILLER_24_577 ();
 FILLER_ASAP7_75t_R FILLER_24_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_611 ();
 DECAPx6_ASAP7_75t_R FILLER_24_640 ();
 DECAPx1_ASAP7_75t_R FILLER_24_654 ();
 DECAPx2_ASAP7_75t_R FILLER_24_664 ();
 FILLER_ASAP7_75t_R FILLER_24_670 ();
 DECAPx2_ASAP7_75t_R FILLER_24_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_693 ();
 DECAPx10_ASAP7_75t_R FILLER_24_697 ();
 DECAPx1_ASAP7_75t_R FILLER_24_731 ();
 DECAPx10_ASAP7_75t_R FILLER_24_741 ();
 DECAPx6_ASAP7_75t_R FILLER_24_763 ();
 DECAPx2_ASAP7_75t_R FILLER_24_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_783 ();
 DECAPx10_ASAP7_75t_R FILLER_24_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_812 ();
 DECAPx10_ASAP7_75t_R FILLER_24_833 ();
 DECAPx10_ASAP7_75t_R FILLER_24_855 ();
 DECAPx10_ASAP7_75t_R FILLER_24_877 ();
 DECAPx1_ASAP7_75t_R FILLER_24_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_903 ();
 DECAPx4_ASAP7_75t_R FILLER_24_910 ();
 FILLER_ASAP7_75t_R FILLER_24_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_943 ();
 DECAPx1_ASAP7_75t_R FILLER_24_968 ();
 DECAPx4_ASAP7_75t_R FILLER_24_974 ();
 FILLER_ASAP7_75t_R FILLER_24_984 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1014 ();
 FILLER_ASAP7_75t_R FILLER_24_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1069 ();
 FILLER_ASAP7_75t_R FILLER_24_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1109 ();
 FILLER_ASAP7_75t_R FILLER_24_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1171 ();
 FILLER_ASAP7_75t_R FILLER_24_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_24_1280 ();
 FILLER_ASAP7_75t_R FILLER_24_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_25_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_534 ();
 DECAPx10_ASAP7_75t_R FILLER_25_548 ();
 DECAPx10_ASAP7_75t_R FILLER_25_570 ();
 FILLER_ASAP7_75t_R FILLER_25_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_594 ();
 DECAPx10_ASAP7_75t_R FILLER_25_601 ();
 DECAPx6_ASAP7_75t_R FILLER_25_623 ();
 FILLER_ASAP7_75t_R FILLER_25_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_639 ();
 DECAPx4_ASAP7_75t_R FILLER_25_650 ();
 FILLER_ASAP7_75t_R FILLER_25_660 ();
 DECAPx10_ASAP7_75t_R FILLER_25_692 ();
 DECAPx10_ASAP7_75t_R FILLER_25_714 ();
 DECAPx6_ASAP7_75t_R FILLER_25_736 ();
 DECAPx2_ASAP7_75t_R FILLER_25_768 ();
 FILLER_ASAP7_75t_R FILLER_25_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_776 ();
 FILLER_ASAP7_75t_R FILLER_25_783 ();
 DECAPx10_ASAP7_75t_R FILLER_25_794 ();
 DECAPx1_ASAP7_75t_R FILLER_25_816 ();
 DECAPx1_ASAP7_75t_R FILLER_25_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_830 ();
 DECAPx10_ASAP7_75t_R FILLER_25_851 ();
 DECAPx10_ASAP7_75t_R FILLER_25_873 ();
 DECAPx2_ASAP7_75t_R FILLER_25_895 ();
 FILLER_ASAP7_75t_R FILLER_25_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_903 ();
 DECAPx10_ASAP7_75t_R FILLER_25_931 ();
 DECAPx10_ASAP7_75t_R FILLER_25_953 ();
 FILLER_ASAP7_75t_R FILLER_25_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_977 ();
 DECAPx1_ASAP7_75t_R FILLER_25_984 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1020 ();
 FILLER_ASAP7_75t_R FILLER_25_1034 ();
 FILLER_ASAP7_75t_R FILLER_25_1042 ();
 FILLER_ASAP7_75t_R FILLER_25_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1052 ();
 FILLER_ASAP7_75t_R FILLER_25_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_25_1103 ();
 FILLER_ASAP7_75t_R FILLER_25_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_25_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_26_512 ();
 DECAPx4_ASAP7_75t_R FILLER_26_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_544 ();
 DECAPx2_ASAP7_75t_R FILLER_26_552 ();
 FILLER_ASAP7_75t_R FILLER_26_558 ();
 DECAPx2_ASAP7_75t_R FILLER_26_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_587 ();
 DECAPx2_ASAP7_75t_R FILLER_26_614 ();
 FILLER_ASAP7_75t_R FILLER_26_620 ();
 DECAPx4_ASAP7_75t_R FILLER_26_643 ();
 FILLER_ASAP7_75t_R FILLER_26_653 ();
 DECAPx6_ASAP7_75t_R FILLER_26_669 ();
 DECAPx1_ASAP7_75t_R FILLER_26_683 ();
 DECAPx6_ASAP7_75t_R FILLER_26_697 ();
 DECAPx1_ASAP7_75t_R FILLER_26_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_715 ();
 DECAPx2_ASAP7_75t_R FILLER_26_722 ();
 FILLER_ASAP7_75t_R FILLER_26_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_730 ();
 DECAPx4_ASAP7_75t_R FILLER_26_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_792 ();
 DECAPx1_ASAP7_75t_R FILLER_26_801 ();
 DECAPx1_ASAP7_75t_R FILLER_26_814 ();
 DECAPx6_ASAP7_75t_R FILLER_26_824 ();
 DECAPx1_ASAP7_75t_R FILLER_26_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_842 ();
 DECAPx10_ASAP7_75t_R FILLER_26_849 ();
 DECAPx10_ASAP7_75t_R FILLER_26_871 ();
 DECAPx2_ASAP7_75t_R FILLER_26_893 ();
 FILLER_ASAP7_75t_R FILLER_26_899 ();
 DECAPx6_ASAP7_75t_R FILLER_26_907 ();
 DECAPx2_ASAP7_75t_R FILLER_26_921 ();
 DECAPx6_ASAP7_75t_R FILLER_26_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_947 ();
 DECAPx1_ASAP7_75t_R FILLER_26_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_971 ();
 DECAPx1_ASAP7_75t_R FILLER_26_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_978 ();
 DECAPx4_ASAP7_75t_R FILLER_26_985 ();
 FILLER_ASAP7_75t_R FILLER_26_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1003 ();
 FILLER_ASAP7_75t_R FILLER_26_1014 ();
 FILLER_ASAP7_75t_R FILLER_26_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1100 ();
 DECAPx4_ASAP7_75t_R FILLER_26_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_26_1146 ();
 FILLER_ASAP7_75t_R FILLER_26_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1181 ();
 FILLER_ASAP7_75t_R FILLER_26_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_26_1281 ();
 FILLER_ASAP7_75t_R FILLER_26_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_27_512 ();
 DECAPx2_ASAP7_75t_R FILLER_27_534 ();
 FILLER_ASAP7_75t_R FILLER_27_540 ();
 FILLER_ASAP7_75t_R FILLER_27_563 ();
 FILLER_ASAP7_75t_R FILLER_27_572 ();
 FILLER_ASAP7_75t_R FILLER_27_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_597 ();
 DECAPx6_ASAP7_75t_R FILLER_27_635 ();
 DECAPx2_ASAP7_75t_R FILLER_27_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_655 ();
 DECAPx4_ASAP7_75t_R FILLER_27_670 ();
 FILLER_ASAP7_75t_R FILLER_27_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_688 ();
 DECAPx2_ASAP7_75t_R FILLER_27_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_711 ();
 DECAPx2_ASAP7_75t_R FILLER_27_735 ();
 FILLER_ASAP7_75t_R FILLER_27_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_753 ();
 DECAPx2_ASAP7_75t_R FILLER_27_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_775 ();
 DECAPx1_ASAP7_75t_R FILLER_27_779 ();
 DECAPx10_ASAP7_75t_R FILLER_27_803 ();
 DECAPx6_ASAP7_75t_R FILLER_27_825 ();
 FILLER_ASAP7_75t_R FILLER_27_839 ();
 DECAPx10_ASAP7_75t_R FILLER_27_851 ();
 DECAPx6_ASAP7_75t_R FILLER_27_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_901 ();
 DECAPx10_ASAP7_75t_R FILLER_27_908 ();
 DECAPx2_ASAP7_75t_R FILLER_27_930 ();
 FILLER_ASAP7_75t_R FILLER_27_936 ();
 DECAPx6_ASAP7_75t_R FILLER_27_965 ();
 FILLER_ASAP7_75t_R FILLER_27_979 ();
 DECAPx2_ASAP7_75t_R FILLER_27_988 ();
 FILLER_ASAP7_75t_R FILLER_27_994 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_27_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_27_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1153 ();
 FILLER_ASAP7_75t_R FILLER_27_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1184 ();
 FILLER_ASAP7_75t_R FILLER_27_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1281 ();
 FILLER_ASAP7_75t_R FILLER_27_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_28_512 ();
 FILLER_ASAP7_75t_R FILLER_28_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_536 ();
 DECAPx4_ASAP7_75t_R FILLER_28_556 ();
 FILLER_ASAP7_75t_R FILLER_28_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_568 ();
 DECAPx6_ASAP7_75t_R FILLER_28_575 ();
 DECAPx1_ASAP7_75t_R FILLER_28_589 ();
 DECAPx10_ASAP7_75t_R FILLER_28_625 ();
 DECAPx1_ASAP7_75t_R FILLER_28_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_651 ();
 FILLER_ASAP7_75t_R FILLER_28_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_666 ();
 DECAPx4_ASAP7_75t_R FILLER_28_673 ();
 FILLER_ASAP7_75t_R FILLER_28_683 ();
 DECAPx4_ASAP7_75t_R FILLER_28_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_723 ();
 DECAPx10_ASAP7_75t_R FILLER_28_730 ();
 DECAPx10_ASAP7_75t_R FILLER_28_752 ();
 DECAPx2_ASAP7_75t_R FILLER_28_774 ();
 FILLER_ASAP7_75t_R FILLER_28_780 ();
 DECAPx4_ASAP7_75t_R FILLER_28_798 ();
 FILLER_ASAP7_75t_R FILLER_28_808 ();
 FILLER_ASAP7_75t_R FILLER_28_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_819 ();
 DECAPx1_ASAP7_75t_R FILLER_28_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_827 ();
 FILLER_ASAP7_75t_R FILLER_28_834 ();
 DECAPx1_ASAP7_75t_R FILLER_28_842 ();
 FILLER_ASAP7_75t_R FILLER_28_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_858 ();
 DECAPx2_ASAP7_75t_R FILLER_28_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_871 ();
 DECAPx4_ASAP7_75t_R FILLER_28_883 ();
 FILLER_ASAP7_75t_R FILLER_28_893 ();
 DECAPx4_ASAP7_75t_R FILLER_28_901 ();
 FILLER_ASAP7_75t_R FILLER_28_911 ();
 DECAPx10_ASAP7_75t_R FILLER_28_933 ();
 DECAPx6_ASAP7_75t_R FILLER_28_955 ();
 FILLER_ASAP7_75t_R FILLER_28_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_974 ();
 FILLER_ASAP7_75t_R FILLER_28_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1001 ();
 FILLER_ASAP7_75t_R FILLER_28_1008 ();
 FILLER_ASAP7_75t_R FILLER_28_1016 ();
 FILLER_ASAP7_75t_R FILLER_28_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_28_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1169 ();
 FILLER_ASAP7_75t_R FILLER_28_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_28_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_29_512 ();
 DECAPx1_ASAP7_75t_R FILLER_29_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_530 ();
 DECAPx10_ASAP7_75t_R FILLER_29_552 ();
 DECAPx10_ASAP7_75t_R FILLER_29_574 ();
 DECAPx10_ASAP7_75t_R FILLER_29_596 ();
 DECAPx10_ASAP7_75t_R FILLER_29_618 ();
 DECAPx10_ASAP7_75t_R FILLER_29_640 ();
 DECAPx1_ASAP7_75t_R FILLER_29_662 ();
 DECAPx10_ASAP7_75t_R FILLER_29_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_700 ();
 DECAPx6_ASAP7_75t_R FILLER_29_714 ();
 FILLER_ASAP7_75t_R FILLER_29_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_730 ();
 DECAPx2_ASAP7_75t_R FILLER_29_737 ();
 FILLER_ASAP7_75t_R FILLER_29_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_745 ();
 DECAPx6_ASAP7_75t_R FILLER_29_752 ();
 DECAPx2_ASAP7_75t_R FILLER_29_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_772 ();
 DECAPx4_ASAP7_75t_R FILLER_29_779 ();
 FILLER_ASAP7_75t_R FILLER_29_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_791 ();
 DECAPx2_ASAP7_75t_R FILLER_29_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_806 ();
 FILLER_ASAP7_75t_R FILLER_29_828 ();
 DECAPx2_ASAP7_75t_R FILLER_29_842 ();
 FILLER_ASAP7_75t_R FILLER_29_848 ();
 FILLER_ASAP7_75t_R FILLER_29_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_859 ();
 DECAPx10_ASAP7_75t_R FILLER_29_882 ();
 DECAPx2_ASAP7_75t_R FILLER_29_904 ();
 FILLER_ASAP7_75t_R FILLER_29_910 ();
 DECAPx4_ASAP7_75t_R FILLER_29_920 ();
 DECAPx10_ASAP7_75t_R FILLER_29_936 ();
 DECAPx10_ASAP7_75t_R FILLER_29_958 ();
 FILLER_ASAP7_75t_R FILLER_29_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_982 ();
 DECAPx6_ASAP7_75t_R FILLER_29_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_29_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_29_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1066 ();
 FILLER_ASAP7_75t_R FILLER_29_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1277 ();
 FILLER_ASAP7_75t_R FILLER_29_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_30_512 ();
 DECAPx6_ASAP7_75t_R FILLER_30_534 ();
 FILLER_ASAP7_75t_R FILLER_30_548 ();
 DECAPx6_ASAP7_75t_R FILLER_30_568 ();
 DECAPx1_ASAP7_75t_R FILLER_30_582 ();
 DECAPx10_ASAP7_75t_R FILLER_30_599 ();
 DECAPx4_ASAP7_75t_R FILLER_30_621 ();
 DECAPx10_ASAP7_75t_R FILLER_30_659 ();
 DECAPx10_ASAP7_75t_R FILLER_30_687 ();
 DECAPx4_ASAP7_75t_R FILLER_30_709 ();
 FILLER_ASAP7_75t_R FILLER_30_719 ();
 DECAPx4_ASAP7_75t_R FILLER_30_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_769 ();
 DECAPx6_ASAP7_75t_R FILLER_30_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_791 ();
 DECAPx6_ASAP7_75t_R FILLER_30_798 ();
 FILLER_ASAP7_75t_R FILLER_30_812 ();
 DECAPx10_ASAP7_75t_R FILLER_30_820 ();
 DECAPx2_ASAP7_75t_R FILLER_30_842 ();
 FILLER_ASAP7_75t_R FILLER_30_848 ();
 DECAPx2_ASAP7_75t_R FILLER_30_875 ();
 FILLER_ASAP7_75t_R FILLER_30_881 ();
 DECAPx2_ASAP7_75t_R FILLER_30_889 ();
 DECAPx1_ASAP7_75t_R FILLER_30_915 ();
 DECAPx2_ASAP7_75t_R FILLER_30_939 ();
 DECAPx2_ASAP7_75t_R FILLER_30_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_961 ();
 DECAPx2_ASAP7_75t_R FILLER_30_974 ();
 DECAPx6_ASAP7_75t_R FILLER_30_990 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1010 ();
 FILLER_ASAP7_75t_R FILLER_30_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1060 ();
 FILLER_ASAP7_75t_R FILLER_30_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_30_1281 ();
 FILLER_ASAP7_75t_R FILLER_30_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_31_512 ();
 DECAPx10_ASAP7_75t_R FILLER_31_534 ();
 FILLER_ASAP7_75t_R FILLER_31_556 ();
 DECAPx1_ASAP7_75t_R FILLER_31_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_584 ();
 DECAPx2_ASAP7_75t_R FILLER_31_606 ();
 FILLER_ASAP7_75t_R FILLER_31_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_614 ();
 DECAPx10_ASAP7_75t_R FILLER_31_621 ();
 DECAPx2_ASAP7_75t_R FILLER_31_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_674 ();
 FILLER_ASAP7_75t_R FILLER_31_693 ();
 DECAPx10_ASAP7_75t_R FILLER_31_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_723 ();
 DECAPx10_ASAP7_75t_R FILLER_31_742 ();
 FILLER_ASAP7_75t_R FILLER_31_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_766 ();
 DECAPx6_ASAP7_75t_R FILLER_31_794 ();
 DECAPx2_ASAP7_75t_R FILLER_31_808 ();
 DECAPx10_ASAP7_75t_R FILLER_31_820 ();
 DECAPx4_ASAP7_75t_R FILLER_31_842 ();
 FILLER_ASAP7_75t_R FILLER_31_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_854 ();
 DECAPx10_ASAP7_75t_R FILLER_31_861 ();
 DECAPx6_ASAP7_75t_R FILLER_31_897 ();
 FILLER_ASAP7_75t_R FILLER_31_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_913 ();
 DECAPx2_ASAP7_75t_R FILLER_31_920 ();
 FILLER_ASAP7_75t_R FILLER_31_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_928 ();
 DECAPx4_ASAP7_75t_R FILLER_31_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_945 ();
 DECAPx2_ASAP7_75t_R FILLER_31_955 ();
 FILLER_ASAP7_75t_R FILLER_31_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_963 ();
 FILLER_ASAP7_75t_R FILLER_31_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_972 ();
 DECAPx10_ASAP7_75t_R FILLER_31_981 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1003 ();
 FILLER_ASAP7_75t_R FILLER_31_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1075 ();
 FILLER_ASAP7_75t_R FILLER_31_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1090 ();
 FILLER_ASAP7_75t_R FILLER_31_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_31_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1149 ();
 FILLER_ASAP7_75t_R FILLER_31_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_31_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_31_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_32_512 ();
 DECAPx4_ASAP7_75t_R FILLER_32_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_544 ();
 DECAPx10_ASAP7_75t_R FILLER_32_587 ();
 DECAPx10_ASAP7_75t_R FILLER_32_609 ();
 DECAPx6_ASAP7_75t_R FILLER_32_631 ();
 DECAPx1_ASAP7_75t_R FILLER_32_645 ();
 DECAPx10_ASAP7_75t_R FILLER_32_661 ();
 DECAPx10_ASAP7_75t_R FILLER_32_683 ();
 FILLER_ASAP7_75t_R FILLER_32_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_707 ();
 DECAPx10_ASAP7_75t_R FILLER_32_717 ();
 DECAPx4_ASAP7_75t_R FILLER_32_739 ();
 FILLER_ASAP7_75t_R FILLER_32_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_751 ();
 DECAPx6_ASAP7_75t_R FILLER_32_781 ();
 DECAPx2_ASAP7_75t_R FILLER_32_795 ();
 DECAPx4_ASAP7_75t_R FILLER_32_815 ();
 FILLER_ASAP7_75t_R FILLER_32_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_827 ();
 DECAPx1_ASAP7_75t_R FILLER_32_855 ();
 DECAPx2_ASAP7_75t_R FILLER_32_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_874 ();
 DECAPx10_ASAP7_75t_R FILLER_32_889 ();
 DECAPx1_ASAP7_75t_R FILLER_32_911 ();
 DECAPx10_ASAP7_75t_R FILLER_32_921 ();
 DECAPx2_ASAP7_75t_R FILLER_32_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_961 ();
 DECAPx1_ASAP7_75t_R FILLER_32_968 ();
 DECAPx6_ASAP7_75t_R FILLER_32_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_988 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1112 ();
 FILLER_ASAP7_75t_R FILLER_32_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1171 ();
 FILLER_ASAP7_75t_R FILLER_32_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1207 ();
 FILLER_ASAP7_75t_R FILLER_32_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1280 ();
 FILLER_ASAP7_75t_R FILLER_32_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_33_512 ();
 DECAPx6_ASAP7_75t_R FILLER_33_534 ();
 DECAPx2_ASAP7_75t_R FILLER_33_548 ();
 DECAPx2_ASAP7_75t_R FILLER_33_557 ();
 FILLER_ASAP7_75t_R FILLER_33_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_565 ();
 DECAPx10_ASAP7_75t_R FILLER_33_579 ();
 DECAPx1_ASAP7_75t_R FILLER_33_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_605 ();
 FILLER_ASAP7_75t_R FILLER_33_634 ();
 DECAPx2_ASAP7_75t_R FILLER_33_664 ();
 FILLER_ASAP7_75t_R FILLER_33_670 ();
 DECAPx10_ASAP7_75t_R FILLER_33_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_718 ();
 DECAPx10_ASAP7_75t_R FILLER_33_761 ();
 DECAPx10_ASAP7_75t_R FILLER_33_783 ();
 DECAPx2_ASAP7_75t_R FILLER_33_805 ();
 DECAPx4_ASAP7_75t_R FILLER_33_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_827 ();
 DECAPx10_ASAP7_75t_R FILLER_33_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_863 ();
 DECAPx2_ASAP7_75t_R FILLER_33_871 ();
 FILLER_ASAP7_75t_R FILLER_33_907 ();
 DECAPx2_ASAP7_75t_R FILLER_33_937 ();
 DECAPx10_ASAP7_75t_R FILLER_33_949 ();
 DECAPx1_ASAP7_75t_R FILLER_33_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1098 ();
 FILLER_ASAP7_75t_R FILLER_33_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1164 ();
 FILLER_ASAP7_75t_R FILLER_33_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_34_512 ();
 DECAPx10_ASAP7_75t_R FILLER_34_534 ();
 DECAPx2_ASAP7_75t_R FILLER_34_556 ();
 FILLER_ASAP7_75t_R FILLER_34_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_564 ();
 DECAPx6_ASAP7_75t_R FILLER_34_572 ();
 FILLER_ASAP7_75t_R FILLER_34_586 ();
 DECAPx10_ASAP7_75t_R FILLER_34_609 ();
 DECAPx10_ASAP7_75t_R FILLER_34_631 ();
 DECAPx10_ASAP7_75t_R FILLER_34_653 ();
 DECAPx1_ASAP7_75t_R FILLER_34_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_679 ();
 DECAPx2_ASAP7_75t_R FILLER_34_692 ();
 FILLER_ASAP7_75t_R FILLER_34_698 ();
 DECAPx10_ASAP7_75t_R FILLER_34_714 ();
 DECAPx10_ASAP7_75t_R FILLER_34_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_758 ();
 DECAPx2_ASAP7_75t_R FILLER_34_773 ();
 FILLER_ASAP7_75t_R FILLER_34_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_793 ();
 DECAPx10_ASAP7_75t_R FILLER_34_816 ();
 DECAPx10_ASAP7_75t_R FILLER_34_838 ();
 DECAPx1_ASAP7_75t_R FILLER_34_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_888 ();
 FILLER_ASAP7_75t_R FILLER_34_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_907 ();
 FILLER_ASAP7_75t_R FILLER_34_914 ();
 DECAPx1_ASAP7_75t_R FILLER_34_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_926 ();
 DECAPx1_ASAP7_75t_R FILLER_34_938 ();
 DECAPx2_ASAP7_75t_R FILLER_34_951 ();
 FILLER_ASAP7_75t_R FILLER_34_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_965 ();
 FILLER_ASAP7_75t_R FILLER_34_980 ();
 DECAPx6_ASAP7_75t_R FILLER_34_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1015 ();
 FILLER_ASAP7_75t_R FILLER_34_1032 ();
 FILLER_ASAP7_75t_R FILLER_34_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1113 ();
 FILLER_ASAP7_75t_R FILLER_34_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_34_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_35_512 ();
 DECAPx10_ASAP7_75t_R FILLER_35_534 ();
 DECAPx2_ASAP7_75t_R FILLER_35_556 ();
 FILLER_ASAP7_75t_R FILLER_35_562 ();
 FILLER_ASAP7_75t_R FILLER_35_585 ();
 DECAPx10_ASAP7_75t_R FILLER_35_600 ();
 DECAPx6_ASAP7_75t_R FILLER_35_622 ();
 DECAPx2_ASAP7_75t_R FILLER_35_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_664 ();
 DECAPx2_ASAP7_75t_R FILLER_35_683 ();
 FILLER_ASAP7_75t_R FILLER_35_689 ();
 FILLER_ASAP7_75t_R FILLER_35_699 ();
 DECAPx10_ASAP7_75t_R FILLER_35_714 ();
 DECAPx1_ASAP7_75t_R FILLER_35_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_740 ();
 DECAPx4_ASAP7_75t_R FILLER_35_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_761 ();
 DECAPx10_ASAP7_75t_R FILLER_35_768 ();
 DECAPx6_ASAP7_75t_R FILLER_35_790 ();
 DECAPx2_ASAP7_75t_R FILLER_35_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_838 ();
 FILLER_ASAP7_75t_R FILLER_35_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_848 ();
 FILLER_ASAP7_75t_R FILLER_35_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_857 ();
 DECAPx2_ASAP7_75t_R FILLER_35_861 ();
 FILLER_ASAP7_75t_R FILLER_35_867 ();
 DECAPx4_ASAP7_75t_R FILLER_35_875 ();
 FILLER_ASAP7_75t_R FILLER_35_885 ();
 DECAPx6_ASAP7_75t_R FILLER_35_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_925 ();
 FILLER_ASAP7_75t_R FILLER_35_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_936 ();
 DECAPx4_ASAP7_75t_R FILLER_35_949 ();
 FILLER_ASAP7_75t_R FILLER_35_959 ();
 DECAPx2_ASAP7_75t_R FILLER_35_969 ();
 FILLER_ASAP7_75t_R FILLER_35_996 ();
 FILLER_ASAP7_75t_R FILLER_35_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1043 ();
 FILLER_ASAP7_75t_R FILLER_35_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1089 ();
 FILLER_ASAP7_75t_R FILLER_35_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1140 ();
 FILLER_ASAP7_75t_R FILLER_35_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1154 ();
 FILLER_ASAP7_75t_R FILLER_35_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_36_512 ();
 DECAPx10_ASAP7_75t_R FILLER_36_534 ();
 DECAPx2_ASAP7_75t_R FILLER_36_556 ();
 FILLER_ASAP7_75t_R FILLER_36_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_564 ();
 DECAPx10_ASAP7_75t_R FILLER_36_571 ();
 DECAPx10_ASAP7_75t_R FILLER_36_593 ();
 DECAPx4_ASAP7_75t_R FILLER_36_615 ();
 FILLER_ASAP7_75t_R FILLER_36_625 ();
 FILLER_ASAP7_75t_R FILLER_36_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_651 ();
 FILLER_ASAP7_75t_R FILLER_36_688 ();
 DECAPx2_ASAP7_75t_R FILLER_36_696 ();
 DECAPx2_ASAP7_75t_R FILLER_36_714 ();
 FILLER_ASAP7_75t_R FILLER_36_720 ();
 DECAPx2_ASAP7_75t_R FILLER_36_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_742 ();
 DECAPx10_ASAP7_75t_R FILLER_36_757 ();
 DECAPx4_ASAP7_75t_R FILLER_36_779 ();
 FILLER_ASAP7_75t_R FILLER_36_789 ();
 DECAPx2_ASAP7_75t_R FILLER_36_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_821 ();
 DECAPx2_ASAP7_75t_R FILLER_36_829 ();
 FILLER_ASAP7_75t_R FILLER_36_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_837 ();
 DECAPx10_ASAP7_75t_R FILLER_36_880 ();
 FILLER_ASAP7_75t_R FILLER_36_902 ();
 DECAPx10_ASAP7_75t_R FILLER_36_910 ();
 DECAPx4_ASAP7_75t_R FILLER_36_932 ();
 DECAPx6_ASAP7_75t_R FILLER_36_956 ();
 FILLER_ASAP7_75t_R FILLER_36_970 ();
 DECAPx10_ASAP7_75t_R FILLER_36_974 ();
 DECAPx10_ASAP7_75t_R FILLER_36_996 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1040 ();
 DECAPx4_ASAP7_75t_R FILLER_36_1062 ();
 FILLER_ASAP7_75t_R FILLER_36_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_36_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1168 ();
 FILLER_ASAP7_75t_R FILLER_36_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_37_512 ();
 DECAPx10_ASAP7_75t_R FILLER_37_534 ();
 DECAPx6_ASAP7_75t_R FILLER_37_556 ();
 DECAPx2_ASAP7_75t_R FILLER_37_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_576 ();
 DECAPx2_ASAP7_75t_R FILLER_37_584 ();
 DECAPx10_ASAP7_75t_R FILLER_37_596 ();
 DECAPx4_ASAP7_75t_R FILLER_37_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_628 ();
 DECAPx10_ASAP7_75t_R FILLER_37_651 ();
 FILLER_ASAP7_75t_R FILLER_37_679 ();
 DECAPx4_ASAP7_75t_R FILLER_37_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_700 ();
 DECAPx2_ASAP7_75t_R FILLER_37_719 ();
 FILLER_ASAP7_75t_R FILLER_37_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_727 ();
 FILLER_ASAP7_75t_R FILLER_37_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_744 ();
 DECAPx6_ASAP7_75t_R FILLER_37_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_765 ();
 FILLER_ASAP7_75t_R FILLER_37_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_774 ();
 FILLER_ASAP7_75t_R FILLER_37_788 ();
 DECAPx1_ASAP7_75t_R FILLER_37_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_802 ();
 DECAPx4_ASAP7_75t_R FILLER_37_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_827 ();
 DECAPx2_ASAP7_75t_R FILLER_37_838 ();
 DECAPx10_ASAP7_75t_R FILLER_37_850 ();
 DECAPx2_ASAP7_75t_R FILLER_37_872 ();
 FILLER_ASAP7_75t_R FILLER_37_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_880 ();
 DECAPx2_ASAP7_75t_R FILLER_37_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_895 ();
 DECAPx1_ASAP7_75t_R FILLER_37_904 ();
 DECAPx10_ASAP7_75t_R FILLER_37_916 ();
 DECAPx6_ASAP7_75t_R FILLER_37_938 ();
 DECAPx6_ASAP7_75t_R FILLER_37_958 ();
 DECAPx1_ASAP7_75t_R FILLER_37_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_976 ();
 DECAPx10_ASAP7_75t_R FILLER_37_983 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1078 ();
 FILLER_ASAP7_75t_R FILLER_37_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1175 ();
 FILLER_ASAP7_75t_R FILLER_37_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1281 ();
 FILLER_ASAP7_75t_R FILLER_37_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_38_512 ();
 DECAPx10_ASAP7_75t_R FILLER_38_534 ();
 DECAPx2_ASAP7_75t_R FILLER_38_556 ();
 DECAPx2_ASAP7_75t_R FILLER_38_569 ();
 DECAPx10_ASAP7_75t_R FILLER_38_596 ();
 DECAPx10_ASAP7_75t_R FILLER_38_618 ();
 DECAPx1_ASAP7_75t_R FILLER_38_640 ();
 DECAPx1_ASAP7_75t_R FILLER_38_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_676 ();
 DECAPx2_ASAP7_75t_R FILLER_38_680 ();
 FILLER_ASAP7_75t_R FILLER_38_686 ();
 FILLER_ASAP7_75t_R FILLER_38_694 ();
 DECAPx10_ASAP7_75t_R FILLER_38_710 ();
 DECAPx6_ASAP7_75t_R FILLER_38_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_746 ();
 DECAPx2_ASAP7_75t_R FILLER_38_763 ();
 DECAPx6_ASAP7_75t_R FILLER_38_775 ();
 DECAPx1_ASAP7_75t_R FILLER_38_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_793 ();
 DECAPx4_ASAP7_75t_R FILLER_38_800 ();
 DECAPx10_ASAP7_75t_R FILLER_38_837 ();
 DECAPx6_ASAP7_75t_R FILLER_38_859 ();
 FILLER_ASAP7_75t_R FILLER_38_873 ();
 DECAPx2_ASAP7_75t_R FILLER_38_889 ();
 DECAPx2_ASAP7_75t_R FILLER_38_901 ();
 DECAPx2_ASAP7_75t_R FILLER_38_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_955 ();
 DECAPx4_ASAP7_75t_R FILLER_38_962 ();
 DECAPx2_ASAP7_75t_R FILLER_38_994 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1269 ();
 FILLER_ASAP7_75t_R FILLER_38_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_39_512 ();
 DECAPx10_ASAP7_75t_R FILLER_39_534 ();
 DECAPx10_ASAP7_75t_R FILLER_39_556 ();
 DECAPx4_ASAP7_75t_R FILLER_39_578 ();
 DECAPx10_ASAP7_75t_R FILLER_39_595 ();
 DECAPx4_ASAP7_75t_R FILLER_39_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_627 ();
 DECAPx6_ASAP7_75t_R FILLER_39_646 ();
 FILLER_ASAP7_75t_R FILLER_39_660 ();
 DECAPx10_ASAP7_75t_R FILLER_39_682 ();
 DECAPx10_ASAP7_75t_R FILLER_39_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_726 ();
 DECAPx1_ASAP7_75t_R FILLER_39_758 ();
 DECAPx6_ASAP7_75t_R FILLER_39_772 ();
 DECAPx2_ASAP7_75t_R FILLER_39_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_792 ();
 DECAPx4_ASAP7_75t_R FILLER_39_799 ();
 FILLER_ASAP7_75t_R FILLER_39_809 ();
 DECAPx6_ASAP7_75t_R FILLER_39_824 ();
 DECAPx2_ASAP7_75t_R FILLER_39_838 ();
 DECAPx2_ASAP7_75t_R FILLER_39_865 ();
 FILLER_ASAP7_75t_R FILLER_39_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_873 ();
 DECAPx2_ASAP7_75t_R FILLER_39_880 ();
 FILLER_ASAP7_75t_R FILLER_39_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_895 ();
 FILLER_ASAP7_75t_R FILLER_39_903 ();
 DECAPx2_ASAP7_75t_R FILLER_39_908 ();
 FILLER_ASAP7_75t_R FILLER_39_914 ();
 FILLER_ASAP7_75t_R FILLER_39_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_928 ();
 DECAPx1_ASAP7_75t_R FILLER_39_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_939 ();
 DECAPx6_ASAP7_75t_R FILLER_39_947 ();
 DECAPx2_ASAP7_75t_R FILLER_39_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_967 ();
 DECAPx4_ASAP7_75t_R FILLER_39_989 ();
 DECAPx4_ASAP7_75t_R FILLER_39_1005 ();
 FILLER_ASAP7_75t_R FILLER_39_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1285 ();
 FILLER_ASAP7_75t_R FILLER_39_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_40_512 ();
 DECAPx10_ASAP7_75t_R FILLER_40_534 ();
 DECAPx4_ASAP7_75t_R FILLER_40_556 ();
 DECAPx4_ASAP7_75t_R FILLER_40_573 ();
 FILLER_ASAP7_75t_R FILLER_40_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_585 ();
 DECAPx10_ASAP7_75t_R FILLER_40_607 ();
 DECAPx6_ASAP7_75t_R FILLER_40_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_643 ();
 DECAPx10_ASAP7_75t_R FILLER_40_662 ();
 DECAPx2_ASAP7_75t_R FILLER_40_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_690 ();
 DECAPx10_ASAP7_75t_R FILLER_40_699 ();
 DECAPx6_ASAP7_75t_R FILLER_40_721 ();
 FILLER_ASAP7_75t_R FILLER_40_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_737 ();
 DECAPx6_ASAP7_75t_R FILLER_40_775 ();
 FILLER_ASAP7_75t_R FILLER_40_789 ();
 DECAPx10_ASAP7_75t_R FILLER_40_799 ();
 DECAPx4_ASAP7_75t_R FILLER_40_821 ();
 FILLER_ASAP7_75t_R FILLER_40_831 ();
 DECAPx10_ASAP7_75t_R FILLER_40_857 ();
 DECAPx2_ASAP7_75t_R FILLER_40_886 ();
 DECAPx6_ASAP7_75t_R FILLER_40_898 ();
 DECAPx2_ASAP7_75t_R FILLER_40_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_918 ();
 DECAPx10_ASAP7_75t_R FILLER_40_925 ();
 DECAPx4_ASAP7_75t_R FILLER_40_947 ();
 DECAPx2_ASAP7_75t_R FILLER_40_964 ();
 FILLER_ASAP7_75t_R FILLER_40_970 ();
 FILLER_ASAP7_75t_R FILLER_40_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_976 ();
 DECAPx2_ASAP7_75t_R FILLER_40_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_993 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_40_1163 ();
 FILLER_ASAP7_75t_R FILLER_40_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1186 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_41_516 ();
 DECAPx10_ASAP7_75t_R FILLER_41_538 ();
 DECAPx1_ASAP7_75t_R FILLER_41_560 ();
 DECAPx2_ASAP7_75t_R FILLER_41_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_591 ();
 DECAPx2_ASAP7_75t_R FILLER_41_598 ();
 FILLER_ASAP7_75t_R FILLER_41_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_606 ();
 DECAPx10_ASAP7_75t_R FILLER_41_628 ();
 DECAPx2_ASAP7_75t_R FILLER_41_650 ();
 FILLER_ASAP7_75t_R FILLER_41_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_686 ();
 DECAPx4_ASAP7_75t_R FILLER_41_697 ();
 DECAPx10_ASAP7_75t_R FILLER_41_729 ();
 DECAPx4_ASAP7_75t_R FILLER_41_751 ();
 FILLER_ASAP7_75t_R FILLER_41_761 ();
 DECAPx6_ASAP7_75t_R FILLER_41_771 ();
 DECAPx1_ASAP7_75t_R FILLER_41_785 ();
 DECAPx10_ASAP7_75t_R FILLER_41_807 ();
 FILLER_ASAP7_75t_R FILLER_41_829 ();
 DECAPx6_ASAP7_75t_R FILLER_41_845 ();
 DECAPx2_ASAP7_75t_R FILLER_41_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_865 ();
 DECAPx1_ASAP7_75t_R FILLER_41_872 ();
 DECAPx4_ASAP7_75t_R FILLER_41_884 ();
 FILLER_ASAP7_75t_R FILLER_41_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_896 ();
 DECAPx2_ASAP7_75t_R FILLER_41_904 ();
 DECAPx10_ASAP7_75t_R FILLER_41_916 ();
 DECAPx6_ASAP7_75t_R FILLER_41_938 ();
 DECAPx1_ASAP7_75t_R FILLER_41_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_956 ();
 DECAPx6_ASAP7_75t_R FILLER_41_964 ();
 DECAPx10_ASAP7_75t_R FILLER_41_986 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1075 ();
 FILLER_ASAP7_75t_R FILLER_41_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1128 ();
 FILLER_ASAP7_75t_R FILLER_41_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1158 ();
 FILLER_ASAP7_75t_R FILLER_41_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_41_1181 ();
 FILLER_ASAP7_75t_R FILLER_41_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_41_1283 ();
 DECAPx6_ASAP7_75t_R FILLER_42_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_532 ();
 DECAPx10_ASAP7_75t_R FILLER_42_539 ();
 DECAPx2_ASAP7_75t_R FILLER_42_561 ();
 FILLER_ASAP7_75t_R FILLER_42_567 ();
 DECAPx10_ASAP7_75t_R FILLER_42_575 ();
 DECAPx4_ASAP7_75t_R FILLER_42_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_607 ();
 DECAPx6_ASAP7_75t_R FILLER_42_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_635 ();
 DECAPx10_ASAP7_75t_R FILLER_42_682 ();
 DECAPx6_ASAP7_75t_R FILLER_42_704 ();
 FILLER_ASAP7_75t_R FILLER_42_718 ();
 DECAPx10_ASAP7_75t_R FILLER_42_736 ();
 DECAPx10_ASAP7_75t_R FILLER_42_758 ();
 DECAPx4_ASAP7_75t_R FILLER_42_780 ();
 FILLER_ASAP7_75t_R FILLER_42_790 ();
 DECAPx2_ASAP7_75t_R FILLER_42_799 ();
 FILLER_ASAP7_75t_R FILLER_42_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_807 ();
 DECAPx10_ASAP7_75t_R FILLER_42_815 ();
 DECAPx10_ASAP7_75t_R FILLER_42_837 ();
 FILLER_ASAP7_75t_R FILLER_42_859 ();
 DECAPx4_ASAP7_75t_R FILLER_42_873 ();
 FILLER_ASAP7_75t_R FILLER_42_883 ();
 DECAPx1_ASAP7_75t_R FILLER_42_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_895 ();
 DECAPx10_ASAP7_75t_R FILLER_42_902 ();
 DECAPx10_ASAP7_75t_R FILLER_42_924 ();
 FILLER_ASAP7_75t_R FILLER_42_946 ();
 FILLER_ASAP7_75t_R FILLER_42_956 ();
 DECAPx2_ASAP7_75t_R FILLER_42_966 ();
 DECAPx10_ASAP7_75t_R FILLER_42_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_996 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1025 ();
 FILLER_ASAP7_75t_R FILLER_42_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1140 ();
 FILLER_ASAP7_75t_R FILLER_42_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1285 ();
 FILLER_ASAP7_75t_R FILLER_42_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_43_512 ();
 FILLER_ASAP7_75t_R FILLER_43_526 ();
 DECAPx6_ASAP7_75t_R FILLER_43_544 ();
 DECAPx1_ASAP7_75t_R FILLER_43_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_562 ();
 DECAPx4_ASAP7_75t_R FILLER_43_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_590 ();
 DECAPx10_ASAP7_75t_R FILLER_43_598 ();
 DECAPx10_ASAP7_75t_R FILLER_43_620 ();
 DECAPx2_ASAP7_75t_R FILLER_43_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_648 ();
 DECAPx10_ASAP7_75t_R FILLER_43_671 ();
 DECAPx10_ASAP7_75t_R FILLER_43_693 ();
 DECAPx2_ASAP7_75t_R FILLER_43_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_777 ();
 DECAPx2_ASAP7_75t_R FILLER_43_784 ();
 FILLER_ASAP7_75t_R FILLER_43_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_792 ();
 DECAPx2_ASAP7_75t_R FILLER_43_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_807 ();
 DECAPx10_ASAP7_75t_R FILLER_43_829 ();
 DECAPx6_ASAP7_75t_R FILLER_43_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_865 ();
 DECAPx4_ASAP7_75t_R FILLER_43_872 ();
 FILLER_ASAP7_75t_R FILLER_43_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_884 ();
 DECAPx1_ASAP7_75t_R FILLER_43_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_952 ();
 DECAPx1_ASAP7_75t_R FILLER_43_979 ();
 DECAPx1_ASAP7_75t_R FILLER_43_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_994 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_43_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_43_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1268 ();
 FILLER_ASAP7_75t_R FILLER_43_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_44_512 ();
 FILLER_ASAP7_75t_R FILLER_44_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_524 ();
 DECAPx2_ASAP7_75t_R FILLER_44_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_547 ();
 FILLER_ASAP7_75t_R FILLER_44_558 ();
 FILLER_ASAP7_75t_R FILLER_44_591 ();
 DECAPx10_ASAP7_75t_R FILLER_44_599 ();
 DECAPx6_ASAP7_75t_R FILLER_44_621 ();
 FILLER_ASAP7_75t_R FILLER_44_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_637 ();
 DECAPx2_ASAP7_75t_R FILLER_44_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_656 ();
 FILLER_ASAP7_75t_R FILLER_44_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_683 ();
 DECAPx6_ASAP7_75t_R FILLER_44_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_712 ();
 DECAPx1_ASAP7_75t_R FILLER_44_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_733 ();
 DECAPx10_ASAP7_75t_R FILLER_44_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_793 ();
 DECAPx4_ASAP7_75t_R FILLER_44_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_819 ();
 DECAPx6_ASAP7_75t_R FILLER_44_823 ();
 DECAPx4_ASAP7_75t_R FILLER_44_855 ();
 DECAPx6_ASAP7_75t_R FILLER_44_875 ();
 FILLER_ASAP7_75t_R FILLER_44_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_891 ();
 DECAPx4_ASAP7_75t_R FILLER_44_899 ();
 FILLER_ASAP7_75t_R FILLER_44_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_911 ();
 DECAPx6_ASAP7_75t_R FILLER_44_932 ();
 DECAPx1_ASAP7_75t_R FILLER_44_946 ();
 DECAPx6_ASAP7_75t_R FILLER_44_958 ();
 FILLER_ASAP7_75t_R FILLER_44_974 ();
 DECAPx2_ASAP7_75t_R FILLER_44_982 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_45_512 ();
 DECAPx10_ASAP7_75t_R FILLER_45_534 ();
 DECAPx1_ASAP7_75t_R FILLER_45_556 ();
 DECAPx1_ASAP7_75t_R FILLER_45_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_577 ();
 DECAPx2_ASAP7_75t_R FILLER_45_584 ();
 FILLER_ASAP7_75t_R FILLER_45_590 ();
 DECAPx4_ASAP7_75t_R FILLER_45_613 ();
 FILLER_ASAP7_75t_R FILLER_45_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_625 ();
 FILLER_ASAP7_75t_R FILLER_45_644 ();
 DECAPx2_ASAP7_75t_R FILLER_45_666 ();
 DECAPx1_ASAP7_75t_R FILLER_45_678 ();
 DECAPx2_ASAP7_75t_R FILLER_45_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_702 ();
 DECAPx2_ASAP7_75t_R FILLER_45_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_724 ();
 DECAPx10_ASAP7_75t_R FILLER_45_756 ();
 FILLER_ASAP7_75t_R FILLER_45_778 ();
 DECAPx10_ASAP7_75t_R FILLER_45_801 ();
 DECAPx1_ASAP7_75t_R FILLER_45_823 ();
 DECAPx4_ASAP7_75t_R FILLER_45_834 ();
 FILLER_ASAP7_75t_R FILLER_45_844 ();
 FILLER_ASAP7_75t_R FILLER_45_862 ();
 FILLER_ASAP7_75t_R FILLER_45_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_876 ();
 DECAPx4_ASAP7_75t_R FILLER_45_890 ();
 FILLER_ASAP7_75t_R FILLER_45_900 ();
 DECAPx6_ASAP7_75t_R FILLER_45_917 ();
 FILLER_ASAP7_75t_R FILLER_45_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_933 ();
 DECAPx2_ASAP7_75t_R FILLER_45_940 ();
 DECAPx2_ASAP7_75t_R FILLER_45_954 ();
 FILLER_ASAP7_75t_R FILLER_45_960 ();
 DECAPx2_ASAP7_75t_R FILLER_45_968 ();
 DECAPx4_ASAP7_75t_R FILLER_45_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_996 ();
 FILLER_ASAP7_75t_R FILLER_45_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1029 ();
 FILLER_ASAP7_75t_R FILLER_45_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1074 ();
 FILLER_ASAP7_75t_R FILLER_45_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1202 ();
 FILLER_ASAP7_75t_R FILLER_45_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_46_512 ();
 DECAPx1_ASAP7_75t_R FILLER_46_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_538 ();
 DECAPx6_ASAP7_75t_R FILLER_46_549 ();
 DECAPx2_ASAP7_75t_R FILLER_46_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_569 ();
 DECAPx10_ASAP7_75t_R FILLER_46_591 ();
 DECAPx10_ASAP7_75t_R FILLER_46_613 ();
 DECAPx10_ASAP7_75t_R FILLER_46_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_657 ();
 DECAPx10_ASAP7_75t_R FILLER_46_672 ();
 DECAPx1_ASAP7_75t_R FILLER_46_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_698 ();
 DECAPx2_ASAP7_75t_R FILLER_46_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_716 ();
 DECAPx2_ASAP7_75t_R FILLER_46_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_730 ();
 DECAPx10_ASAP7_75t_R FILLER_46_737 ();
 DECAPx2_ASAP7_75t_R FILLER_46_759 ();
 DECAPx2_ASAP7_75t_R FILLER_46_772 ();
 FILLER_ASAP7_75t_R FILLER_46_778 ();
 DECAPx4_ASAP7_75t_R FILLER_46_787 ();
 FILLER_ASAP7_75t_R FILLER_46_797 ();
 DECAPx6_ASAP7_75t_R FILLER_46_813 ();
 DECAPx10_ASAP7_75t_R FILLER_46_833 ();
 DECAPx6_ASAP7_75t_R FILLER_46_855 ();
 FILLER_ASAP7_75t_R FILLER_46_869 ();
 FILLER_ASAP7_75t_R FILLER_46_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_889 ();
 DECAPx10_ASAP7_75t_R FILLER_46_919 ();
 DECAPx2_ASAP7_75t_R FILLER_46_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_947 ();
 DECAPx2_ASAP7_75t_R FILLER_46_964 ();
 FILLER_ASAP7_75t_R FILLER_46_970 ();
 DECAPx2_ASAP7_75t_R FILLER_46_981 ();
 FILLER_ASAP7_75t_R FILLER_46_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_989 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1038 ();
 FILLER_ASAP7_75t_R FILLER_46_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1084 ();
 FILLER_ASAP7_75t_R FILLER_46_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1243 ();
 FILLER_ASAP7_75t_R FILLER_46_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1276 ();
 FILLER_ASAP7_75t_R FILLER_46_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_47_512 ();
 DECAPx10_ASAP7_75t_R FILLER_47_534 ();
 DECAPx6_ASAP7_75t_R FILLER_47_556 ();
 FILLER_ASAP7_75t_R FILLER_47_570 ();
 DECAPx6_ASAP7_75t_R FILLER_47_579 ();
 DECAPx1_ASAP7_75t_R FILLER_47_593 ();
 DECAPx4_ASAP7_75t_R FILLER_47_618 ();
 FILLER_ASAP7_75t_R FILLER_47_628 ();
 DECAPx10_ASAP7_75t_R FILLER_47_633 ();
 DECAPx6_ASAP7_75t_R FILLER_47_655 ();
 DECAPx1_ASAP7_75t_R FILLER_47_669 ();
 DECAPx1_ASAP7_75t_R FILLER_47_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_700 ();
 DECAPx10_ASAP7_75t_R FILLER_47_708 ();
 DECAPx6_ASAP7_75t_R FILLER_47_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_751 ();
 FILLER_ASAP7_75t_R FILLER_47_779 ();
 DECAPx4_ASAP7_75t_R FILLER_47_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_805 ();
 DECAPx4_ASAP7_75t_R FILLER_47_819 ();
 DECAPx10_ASAP7_75t_R FILLER_47_892 ();
 DECAPx10_ASAP7_75t_R FILLER_47_914 ();
 DECAPx10_ASAP7_75t_R FILLER_47_936 ();
 DECAPx4_ASAP7_75t_R FILLER_47_958 ();
 FILLER_ASAP7_75t_R FILLER_47_968 ();
 FILLER_ASAP7_75t_R FILLER_47_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_993 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1118 ();
 FILLER_ASAP7_75t_R FILLER_47_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_48_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_522 ();
 DECAPx1_ASAP7_75t_R FILLER_48_547 ();
 DECAPx1_ASAP7_75t_R FILLER_48_593 ();
 DECAPx1_ASAP7_75t_R FILLER_48_604 ();
 DECAPx2_ASAP7_75t_R FILLER_48_614 ();
 DECAPx4_ASAP7_75t_R FILLER_48_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_636 ();
 DECAPx10_ASAP7_75t_R FILLER_48_643 ();
 DECAPx1_ASAP7_75t_R FILLER_48_665 ();
 DECAPx6_ASAP7_75t_R FILLER_48_687 ();
 DECAPx6_ASAP7_75t_R FILLER_48_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_728 ();
 DECAPx6_ASAP7_75t_R FILLER_48_750 ();
 DECAPx1_ASAP7_75t_R FILLER_48_764 ();
 DECAPx2_ASAP7_75t_R FILLER_48_795 ();
 FILLER_ASAP7_75t_R FILLER_48_801 ();
 FILLER_ASAP7_75t_R FILLER_48_824 ();
 DECAPx1_ASAP7_75t_R FILLER_48_832 ();
 DECAPx10_ASAP7_75t_R FILLER_48_842 ();
 DECAPx10_ASAP7_75t_R FILLER_48_864 ();
 DECAPx4_ASAP7_75t_R FILLER_48_886 ();
 FILLER_ASAP7_75t_R FILLER_48_896 ();
 DECAPx10_ASAP7_75t_R FILLER_48_904 ();
 DECAPx10_ASAP7_75t_R FILLER_48_926 ();
 DECAPx10_ASAP7_75t_R FILLER_48_948 ();
 FILLER_ASAP7_75t_R FILLER_48_970 ();
 FILLER_ASAP7_75t_R FILLER_48_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_976 ();
 DECAPx4_ASAP7_75t_R FILLER_48_983 ();
 FILLER_ASAP7_75t_R FILLER_48_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_995 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1017 ();
 FILLER_ASAP7_75t_R FILLER_48_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1042 ();
 FILLER_ASAP7_75t_R FILLER_48_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1066 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1099 ();
 FILLER_ASAP7_75t_R FILLER_48_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1148 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1281 ();
 FILLER_ASAP7_75t_R FILLER_48_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_49_512 ();
 FILLER_ASAP7_75t_R FILLER_49_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_528 ();
 DECAPx2_ASAP7_75t_R FILLER_49_550 ();
 DECAPx4_ASAP7_75t_R FILLER_49_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_573 ();
 DECAPx10_ASAP7_75t_R FILLER_49_580 ();
 FILLER_ASAP7_75t_R FILLER_49_602 ();
 DECAPx2_ASAP7_75t_R FILLER_49_625 ();
 DECAPx2_ASAP7_75t_R FILLER_49_649 ();
 DECAPx10_ASAP7_75t_R FILLER_49_662 ();
 FILLER_ASAP7_75t_R FILLER_49_684 ();
 DECAPx6_ASAP7_75t_R FILLER_49_707 ();
 DECAPx1_ASAP7_75t_R FILLER_49_728 ();
 DECAPx10_ASAP7_75t_R FILLER_49_738 ();
 DECAPx1_ASAP7_75t_R FILLER_49_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_764 ();
 DECAPx2_ASAP7_75t_R FILLER_49_768 ();
 DECAPx10_ASAP7_75t_R FILLER_49_807 ();
 DECAPx4_ASAP7_75t_R FILLER_49_835 ();
 FILLER_ASAP7_75t_R FILLER_49_845 ();
 DECAPx10_ASAP7_75t_R FILLER_49_854 ();
 DECAPx6_ASAP7_75t_R FILLER_49_876 ();
 DECAPx2_ASAP7_75t_R FILLER_49_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_896 ();
 DECAPx2_ASAP7_75t_R FILLER_49_905 ();
 FILLER_ASAP7_75t_R FILLER_49_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_934 ();
 DECAPx1_ASAP7_75t_R FILLER_49_953 ();
 DECAPx10_ASAP7_75t_R FILLER_49_978 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1000 ();
 FILLER_ASAP7_75t_R FILLER_49_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1081 ();
 FILLER_ASAP7_75t_R FILLER_49_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1089 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1100 ();
 FILLER_ASAP7_75t_R FILLER_49_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_49_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1199 ();
 FILLER_ASAP7_75t_R FILLER_49_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_50_512 ();
 FILLER_ASAP7_75t_R FILLER_50_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_536 ();
 DECAPx6_ASAP7_75t_R FILLER_50_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_557 ();
 DECAPx10_ASAP7_75t_R FILLER_50_564 ();
 DECAPx10_ASAP7_75t_R FILLER_50_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_608 ();
 DECAPx10_ASAP7_75t_R FILLER_50_615 ();
 DECAPx4_ASAP7_75t_R FILLER_50_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_647 ();
 DECAPx2_ASAP7_75t_R FILLER_50_654 ();
 DECAPx6_ASAP7_75t_R FILLER_50_666 ();
 DECAPx1_ASAP7_75t_R FILLER_50_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_684 ();
 DECAPx6_ASAP7_75t_R FILLER_50_692 ();
 DECAPx10_ASAP7_75t_R FILLER_50_733 ();
 DECAPx6_ASAP7_75t_R FILLER_50_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_769 ();
 DECAPx4_ASAP7_75t_R FILLER_50_796 ();
 FILLER_ASAP7_75t_R FILLER_50_806 ();
 DECAPx10_ASAP7_75t_R FILLER_50_818 ();
 DECAPx2_ASAP7_75t_R FILLER_50_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_846 ();
 DECAPx6_ASAP7_75t_R FILLER_50_853 ();
 DECAPx4_ASAP7_75t_R FILLER_50_880 ();
 DECAPx2_ASAP7_75t_R FILLER_50_904 ();
 FILLER_ASAP7_75t_R FILLER_50_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_919 ();
 DECAPx4_ASAP7_75t_R FILLER_50_929 ();
 FILLER_ASAP7_75t_R FILLER_50_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_941 ();
 DECAPx1_ASAP7_75t_R FILLER_50_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_974 ();
 DECAPx6_ASAP7_75t_R FILLER_50_996 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1014 ();
 FILLER_ASAP7_75t_R FILLER_50_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1047 ();
 FILLER_ASAP7_75t_R FILLER_50_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1067 ();
 FILLER_ASAP7_75t_R FILLER_50_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1217 ();
 FILLER_ASAP7_75t_R FILLER_50_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1236 ();
 FILLER_ASAP7_75t_R FILLER_50_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1244 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_51_512 ();
 DECAPx6_ASAP7_75t_R FILLER_51_534 ();
 FILLER_ASAP7_75t_R FILLER_51_548 ();
 DECAPx10_ASAP7_75t_R FILLER_51_560 ();
 DECAPx10_ASAP7_75t_R FILLER_51_582 ();
 DECAPx10_ASAP7_75t_R FILLER_51_604 ();
 DECAPx6_ASAP7_75t_R FILLER_51_626 ();
 DECAPx2_ASAP7_75t_R FILLER_51_640 ();
 DECAPx6_ASAP7_75t_R FILLER_51_654 ();
 DECAPx4_ASAP7_75t_R FILLER_51_692 ();
 FILLER_ASAP7_75t_R FILLER_51_702 ();
 DECAPx2_ASAP7_75t_R FILLER_51_718 ();
 DECAPx2_ASAP7_75t_R FILLER_51_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_742 ();
 FILLER_ASAP7_75t_R FILLER_51_767 ();
 DECAPx10_ASAP7_75t_R FILLER_51_775 ();
 DECAPx4_ASAP7_75t_R FILLER_51_797 ();
 FILLER_ASAP7_75t_R FILLER_51_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_809 ();
 DECAPx10_ASAP7_75t_R FILLER_51_818 ();
 DECAPx2_ASAP7_75t_R FILLER_51_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_846 ();
 DECAPx6_ASAP7_75t_R FILLER_51_889 ();
 DECAPx1_ASAP7_75t_R FILLER_51_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_907 ();
 DECAPx2_ASAP7_75t_R FILLER_51_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_921 ();
 DECAPx10_ASAP7_75t_R FILLER_51_928 ();
 DECAPx10_ASAP7_75t_R FILLER_51_950 ();
 DECAPx6_ASAP7_75t_R FILLER_51_972 ();
 DECAPx1_ASAP7_75t_R FILLER_51_986 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1008 ();
 FILLER_ASAP7_75t_R FILLER_51_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1029 ();
 FILLER_ASAP7_75t_R FILLER_51_1051 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1061 ();
 FILLER_ASAP7_75t_R FILLER_51_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1122 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1129 ();
 FILLER_ASAP7_75t_R FILLER_51_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_51_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1265 ();
 DECAPx6_ASAP7_75t_R FILLER_51_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_512 ();
 DECAPx10_ASAP7_75t_R FILLER_52_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_547 ();
 DECAPx2_ASAP7_75t_R FILLER_52_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_560 ();
 DECAPx2_ASAP7_75t_R FILLER_52_582 ();
 FILLER_ASAP7_75t_R FILLER_52_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_590 ();
 FILLER_ASAP7_75t_R FILLER_52_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_600 ();
 DECAPx10_ASAP7_75t_R FILLER_52_622 ();
 DECAPx10_ASAP7_75t_R FILLER_52_644 ();
 DECAPx10_ASAP7_75t_R FILLER_52_666 ();
 DECAPx10_ASAP7_75t_R FILLER_52_688 ();
 DECAPx10_ASAP7_75t_R FILLER_52_710 ();
 DECAPx2_ASAP7_75t_R FILLER_52_748 ();
 FILLER_ASAP7_75t_R FILLER_52_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_756 ();
 DECAPx4_ASAP7_75t_R FILLER_52_764 ();
 FILLER_ASAP7_75t_R FILLER_52_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_776 ();
 DECAPx10_ASAP7_75t_R FILLER_52_784 ();
 DECAPx6_ASAP7_75t_R FILLER_52_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_820 ();
 DECAPx10_ASAP7_75t_R FILLER_52_827 ();
 DECAPx10_ASAP7_75t_R FILLER_52_849 ();
 DECAPx10_ASAP7_75t_R FILLER_52_871 ();
 DECAPx6_ASAP7_75t_R FILLER_52_893 ();
 DECAPx1_ASAP7_75t_R FILLER_52_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_911 ();
 DECAPx4_ASAP7_75t_R FILLER_52_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_928 ();
 DECAPx6_ASAP7_75t_R FILLER_52_935 ();
 FILLER_ASAP7_75t_R FILLER_52_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_951 ();
 FILLER_ASAP7_75t_R FILLER_52_959 ();
 DECAPx1_ASAP7_75t_R FILLER_52_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_971 ();
 DECAPx10_ASAP7_75t_R FILLER_52_974 ();
 FILLER_ASAP7_75t_R FILLER_52_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_998 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1053 ();
 FILLER_ASAP7_75t_R FILLER_52_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1128 ();
 FILLER_ASAP7_75t_R FILLER_52_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1173 ();
 FILLER_ASAP7_75t_R FILLER_52_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_53_512 ();
 FILLER_ASAP7_75t_R FILLER_53_526 ();
 DECAPx1_ASAP7_75t_R FILLER_53_557 ();
 FILLER_ASAP7_75t_R FILLER_53_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_572 ();
 FILLER_ASAP7_75t_R FILLER_53_576 ();
 FILLER_ASAP7_75t_R FILLER_53_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_588 ();
 DECAPx10_ASAP7_75t_R FILLER_53_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_623 ();
 DECAPx6_ASAP7_75t_R FILLER_53_660 ();
 DECAPx2_ASAP7_75t_R FILLER_53_674 ();
 DECAPx1_ASAP7_75t_R FILLER_53_724 ();
 DECAPx1_ASAP7_75t_R FILLER_53_734 ();
 DECAPx2_ASAP7_75t_R FILLER_53_744 ();
 FILLER_ASAP7_75t_R FILLER_53_750 ();
 FILLER_ASAP7_75t_R FILLER_53_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_775 ();
 DECAPx6_ASAP7_75t_R FILLER_53_803 ();
 DECAPx1_ASAP7_75t_R FILLER_53_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_821 ();
 DECAPx6_ASAP7_75t_R FILLER_53_828 ();
 DECAPx1_ASAP7_75t_R FILLER_53_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_846 ();
 DECAPx10_ASAP7_75t_R FILLER_53_854 ();
 DECAPx6_ASAP7_75t_R FILLER_53_876 ();
 DECAPx2_ASAP7_75t_R FILLER_53_890 ();
 DECAPx1_ASAP7_75t_R FILLER_53_931 ();
 DECAPx1_ASAP7_75t_R FILLER_53_949 ();
 DECAPx4_ASAP7_75t_R FILLER_53_974 ();
 FILLER_ASAP7_75t_R FILLER_53_984 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1016 ();
 FILLER_ASAP7_75t_R FILLER_53_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1069 ();
 FILLER_ASAP7_75t_R FILLER_53_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1083 ();
 FILLER_ASAP7_75t_R FILLER_53_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1160 ();
 FILLER_ASAP7_75t_R FILLER_53_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1176 ();
 FILLER_ASAP7_75t_R FILLER_53_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1221 ();
 FILLER_ASAP7_75t_R FILLER_53_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_54_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_534 ();
 DECAPx2_ASAP7_75t_R FILLER_54_552 ();
 FILLER_ASAP7_75t_R FILLER_54_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_560 ();
 DECAPx2_ASAP7_75t_R FILLER_54_567 ();
 FILLER_ASAP7_75t_R FILLER_54_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_575 ();
 DECAPx10_ASAP7_75t_R FILLER_54_597 ();
 DECAPx10_ASAP7_75t_R FILLER_54_619 ();
 FILLER_ASAP7_75t_R FILLER_54_641 ();
 DECAPx6_ASAP7_75t_R FILLER_54_653 ();
 DECAPx2_ASAP7_75t_R FILLER_54_667 ();
 DECAPx2_ASAP7_75t_R FILLER_54_682 ();
 FILLER_ASAP7_75t_R FILLER_54_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_690 ();
 DECAPx1_ASAP7_75t_R FILLER_54_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_715 ();
 FILLER_ASAP7_75t_R FILLER_54_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_728 ();
 DECAPx10_ASAP7_75t_R FILLER_54_735 ();
 DECAPx4_ASAP7_75t_R FILLER_54_757 ();
 FILLER_ASAP7_75t_R FILLER_54_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_769 ();
 DECAPx10_ASAP7_75t_R FILLER_54_783 ();
 DECAPx10_ASAP7_75t_R FILLER_54_805 ();
 FILLER_ASAP7_75t_R FILLER_54_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_829 ();
 DECAPx2_ASAP7_75t_R FILLER_54_837 ();
 FILLER_ASAP7_75t_R FILLER_54_843 ();
 DECAPx4_ASAP7_75t_R FILLER_54_866 ();
 FILLER_ASAP7_75t_R FILLER_54_876 ();
 DECAPx10_ASAP7_75t_R FILLER_54_888 ();
 DECAPx10_ASAP7_75t_R FILLER_54_910 ();
 DECAPx4_ASAP7_75t_R FILLER_54_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_942 ();
 DECAPx10_ASAP7_75t_R FILLER_54_950 ();
 DECAPx2_ASAP7_75t_R FILLER_54_974 ();
 FILLER_ASAP7_75t_R FILLER_54_980 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1132 ();
 FILLER_ASAP7_75t_R FILLER_54_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1209 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_55_512 ();
 DECAPx10_ASAP7_75t_R FILLER_55_534 ();
 DECAPx6_ASAP7_75t_R FILLER_55_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_570 ();
 DECAPx10_ASAP7_75t_R FILLER_55_604 ();
 DECAPx6_ASAP7_75t_R FILLER_55_626 ();
 DECAPx2_ASAP7_75t_R FILLER_55_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_646 ();
 DECAPx10_ASAP7_75t_R FILLER_55_656 ();
 DECAPx10_ASAP7_75t_R FILLER_55_678 ();
 DECAPx6_ASAP7_75t_R FILLER_55_700 ();
 FILLER_ASAP7_75t_R FILLER_55_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_716 ();
 DECAPx10_ASAP7_75t_R FILLER_55_737 ();
 DECAPx2_ASAP7_75t_R FILLER_55_759 ();
 FILLER_ASAP7_75t_R FILLER_55_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_767 ();
 DECAPx6_ASAP7_75t_R FILLER_55_796 ();
 DECAPx4_ASAP7_75t_R FILLER_55_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_856 ();
 DECAPx10_ASAP7_75t_R FILLER_55_863 ();
 DECAPx2_ASAP7_75t_R FILLER_55_885 ();
 FILLER_ASAP7_75t_R FILLER_55_891 ();
 DECAPx10_ASAP7_75t_R FILLER_55_914 ();
 DECAPx2_ASAP7_75t_R FILLER_55_936 ();
 FILLER_ASAP7_75t_R FILLER_55_942 ();
 DECAPx10_ASAP7_75t_R FILLER_55_965 ();
 DECAPx4_ASAP7_75t_R FILLER_55_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1080 ();
 FILLER_ASAP7_75t_R FILLER_55_1091 ();
 FILLER_ASAP7_75t_R FILLER_55_1099 ();
 FILLER_ASAP7_75t_R FILLER_55_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_55_1126 ();
 FILLER_ASAP7_75t_R FILLER_55_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_55_1191 ();
 FILLER_ASAP7_75t_R FILLER_55_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1256 ();
 FILLER_ASAP7_75t_R FILLER_55_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_56_512 ();
 DECAPx1_ASAP7_75t_R FILLER_56_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_549 ();
 DECAPx4_ASAP7_75t_R FILLER_56_571 ();
 FILLER_ASAP7_75t_R FILLER_56_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_583 ();
 DECAPx6_ASAP7_75t_R FILLER_56_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_605 ();
 DECAPx2_ASAP7_75t_R FILLER_56_613 ();
 FILLER_ASAP7_75t_R FILLER_56_619 ();
 DECAPx10_ASAP7_75t_R FILLER_56_627 ();
 DECAPx2_ASAP7_75t_R FILLER_56_649 ();
 DECAPx10_ASAP7_75t_R FILLER_56_661 ();
 DECAPx2_ASAP7_75t_R FILLER_56_683 ();
 DECAPx10_ASAP7_75t_R FILLER_56_705 ();
 DECAPx1_ASAP7_75t_R FILLER_56_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_744 ();
 DECAPx2_ASAP7_75t_R FILLER_56_752 ();
 FILLER_ASAP7_75t_R FILLER_56_758 ();
 DECAPx1_ASAP7_75t_R FILLER_56_767 ();
 DECAPx2_ASAP7_75t_R FILLER_56_783 ();
 FILLER_ASAP7_75t_R FILLER_56_831 ();
 DECAPx6_ASAP7_75t_R FILLER_56_839 ();
 DECAPx1_ASAP7_75t_R FILLER_56_853 ();
 DECAPx2_ASAP7_75t_R FILLER_56_885 ();
 FILLER_ASAP7_75t_R FILLER_56_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_893 ();
 FILLER_ASAP7_75t_R FILLER_56_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_909 ();
 FILLER_ASAP7_75t_R FILLER_56_920 ();
 FILLER_ASAP7_75t_R FILLER_56_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_932 ();
 DECAPx6_ASAP7_75t_R FILLER_56_936 ();
 DECAPx1_ASAP7_75t_R FILLER_56_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_954 ();
 DECAPx2_ASAP7_75t_R FILLER_56_964 ();
 FILLER_ASAP7_75t_R FILLER_56_970 ();
 DECAPx10_ASAP7_75t_R FILLER_56_974 ();
 DECAPx1_ASAP7_75t_R FILLER_56_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1076 ();
 FILLER_ASAP7_75t_R FILLER_56_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1230 ();
 FILLER_ASAP7_75t_R FILLER_56_1236 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1244 ();
 FILLER_ASAP7_75t_R FILLER_56_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_57_512 ();
 FILLER_ASAP7_75t_R FILLER_57_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_528 ();
 FILLER_ASAP7_75t_R FILLER_57_547 ();
 DECAPx4_ASAP7_75t_R FILLER_57_562 ();
 DECAPx1_ASAP7_75t_R FILLER_57_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_628 ();
 DECAPx2_ASAP7_75t_R FILLER_57_647 ();
 FILLER_ASAP7_75t_R FILLER_57_653 ();
 DECAPx1_ASAP7_75t_R FILLER_57_669 ();
 FILLER_ASAP7_75t_R FILLER_57_691 ();
 DECAPx2_ASAP7_75t_R FILLER_57_701 ();
 FILLER_ASAP7_75t_R FILLER_57_707 ();
 FILLER_ASAP7_75t_R FILLER_57_737 ();
 DECAPx2_ASAP7_75t_R FILLER_57_755 ();
 DECAPx10_ASAP7_75t_R FILLER_57_767 ();
 DECAPx2_ASAP7_75t_R FILLER_57_789 ();
 DECAPx4_ASAP7_75t_R FILLER_57_801 ();
 FILLER_ASAP7_75t_R FILLER_57_811 ();
 DECAPx10_ASAP7_75t_R FILLER_57_819 ();
 DECAPx10_ASAP7_75t_R FILLER_57_841 ();
 DECAPx6_ASAP7_75t_R FILLER_57_863 ();
 DECAPx1_ASAP7_75t_R FILLER_57_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_881 ();
 DECAPx2_ASAP7_75t_R FILLER_57_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_912 ();
 DECAPx6_ASAP7_75t_R FILLER_57_940 ();
 DECAPx1_ASAP7_75t_R FILLER_57_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_958 ();
 DECAPx2_ASAP7_75t_R FILLER_57_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_979 ();
 DECAPx4_ASAP7_75t_R FILLER_57_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1232 ();
 FILLER_ASAP7_75t_R FILLER_57_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1269 ();
 FILLER_ASAP7_75t_R FILLER_57_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_58_512 ();
 DECAPx1_ASAP7_75t_R FILLER_58_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_530 ();
 FILLER_ASAP7_75t_R FILLER_58_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_543 ();
 DECAPx6_ASAP7_75t_R FILLER_58_554 ();
 FILLER_ASAP7_75t_R FILLER_58_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_570 ();
 DECAPx4_ASAP7_75t_R FILLER_58_578 ();
 FILLER_ASAP7_75t_R FILLER_58_588 ();
 DECAPx10_ASAP7_75t_R FILLER_58_596 ();
 DECAPx6_ASAP7_75t_R FILLER_58_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_632 ();
 DECAPx10_ASAP7_75t_R FILLER_58_673 ();
 DECAPx4_ASAP7_75t_R FILLER_58_695 ();
 FILLER_ASAP7_75t_R FILLER_58_705 ();
 DECAPx2_ASAP7_75t_R FILLER_58_719 ();
 FILLER_ASAP7_75t_R FILLER_58_725 ();
 DECAPx6_ASAP7_75t_R FILLER_58_741 ();
 DECAPx1_ASAP7_75t_R FILLER_58_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_759 ();
 DECAPx10_ASAP7_75t_R FILLER_58_788 ();
 DECAPx6_ASAP7_75t_R FILLER_58_810 ();
 DECAPx1_ASAP7_75t_R FILLER_58_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_828 ();
 DECAPx6_ASAP7_75t_R FILLER_58_836 ();
 DECAPx10_ASAP7_75t_R FILLER_58_862 ();
 DECAPx4_ASAP7_75t_R FILLER_58_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_894 ();
 DECAPx2_ASAP7_75t_R FILLER_58_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_931 ();
 DECAPx10_ASAP7_75t_R FILLER_58_938 ();
 DECAPx4_ASAP7_75t_R FILLER_58_960 ();
 FILLER_ASAP7_75t_R FILLER_58_970 ();
 FILLER_ASAP7_75t_R FILLER_58_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_990 ();
 FILLER_ASAP7_75t_R FILLER_58_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_58_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1079 ();
 FILLER_ASAP7_75t_R FILLER_58_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1149 ();
 FILLER_ASAP7_75t_R FILLER_58_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1202 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1238 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_59_512 ();
 DECAPx10_ASAP7_75t_R FILLER_59_534 ();
 DECAPx6_ASAP7_75t_R FILLER_59_556 ();
 FILLER_ASAP7_75t_R FILLER_59_570 ();
 DECAPx10_ASAP7_75t_R FILLER_59_600 ();
 DECAPx6_ASAP7_75t_R FILLER_59_622 ();
 DECAPx2_ASAP7_75t_R FILLER_59_658 ();
 FILLER_ASAP7_75t_R FILLER_59_664 ();
 DECAPx4_ASAP7_75t_R FILLER_59_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_684 ();
 DECAPx10_ASAP7_75t_R FILLER_59_691 ();
 DECAPx4_ASAP7_75t_R FILLER_59_713 ();
 FILLER_ASAP7_75t_R FILLER_59_723 ();
 DECAPx10_ASAP7_75t_R FILLER_59_741 ();
 DECAPx6_ASAP7_75t_R FILLER_59_763 ();
 DECAPx10_ASAP7_75t_R FILLER_59_798 ();
 DECAPx2_ASAP7_75t_R FILLER_59_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_826 ();
 FILLER_ASAP7_75t_R FILLER_59_854 ();
 DECAPx10_ASAP7_75t_R FILLER_59_865 ();
 DECAPx2_ASAP7_75t_R FILLER_59_887 ();
 FILLER_ASAP7_75t_R FILLER_59_893 ();
 DECAPx4_ASAP7_75t_R FILLER_59_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_913 ();
 DECAPx6_ASAP7_75t_R FILLER_59_921 ();
 DECAPx1_ASAP7_75t_R FILLER_59_935 ();
 FILLER_ASAP7_75t_R FILLER_59_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_954 ();
 DECAPx6_ASAP7_75t_R FILLER_59_966 ();
 DECAPx2_ASAP7_75t_R FILLER_59_996 ();
 FILLER_ASAP7_75t_R FILLER_59_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1013 ();
 FILLER_ASAP7_75t_R FILLER_59_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1048 ();
 FILLER_ASAP7_75t_R FILLER_59_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1060 ();
 FILLER_ASAP7_75t_R FILLER_59_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1080 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1098 ();
 FILLER_ASAP7_75t_R FILLER_59_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1116 ();
 FILLER_ASAP7_75t_R FILLER_59_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1127 ();
 FILLER_ASAP7_75t_R FILLER_59_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1140 ();
 FILLER_ASAP7_75t_R FILLER_59_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1280 ();
 FILLER_ASAP7_75t_R FILLER_59_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_60_512 ();
 DECAPx6_ASAP7_75t_R FILLER_60_534 ();
 DECAPx1_ASAP7_75t_R FILLER_60_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_552 ();
 DECAPx4_ASAP7_75t_R FILLER_60_559 ();
 FILLER_ASAP7_75t_R FILLER_60_569 ();
 DECAPx2_ASAP7_75t_R FILLER_60_577 ();
 DECAPx10_ASAP7_75t_R FILLER_60_612 ();
 DECAPx4_ASAP7_75t_R FILLER_60_634 ();
 FILLER_ASAP7_75t_R FILLER_60_644 ();
 DECAPx2_ASAP7_75t_R FILLER_60_691 ();
 FILLER_ASAP7_75t_R FILLER_60_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_699 ();
 FILLER_ASAP7_75t_R FILLER_60_715 ();
 DECAPx4_ASAP7_75t_R FILLER_60_723 ();
 FILLER_ASAP7_75t_R FILLER_60_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_735 ();
 DECAPx2_ASAP7_75t_R FILLER_60_750 ();
 DECAPx10_ASAP7_75t_R FILLER_60_762 ();
 FILLER_ASAP7_75t_R FILLER_60_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_786 ();
 DECAPx6_ASAP7_75t_R FILLER_60_793 ();
 DECAPx1_ASAP7_75t_R FILLER_60_807 ();
 DECAPx2_ASAP7_75t_R FILLER_60_821 ();
 FILLER_ASAP7_75t_R FILLER_60_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_829 ();
 DECAPx4_ASAP7_75t_R FILLER_60_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_846 ();
 DECAPx1_ASAP7_75t_R FILLER_60_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_857 ();
 DECAPx6_ASAP7_75t_R FILLER_60_864 ();
 FILLER_ASAP7_75t_R FILLER_60_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_880 ();
 DECAPx6_ASAP7_75t_R FILLER_60_887 ();
 FILLER_ASAP7_75t_R FILLER_60_901 ();
 DECAPx4_ASAP7_75t_R FILLER_60_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_921 ();
 DECAPx4_ASAP7_75t_R FILLER_60_928 ();
 DECAPx2_ASAP7_75t_R FILLER_60_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_971 ();
 DECAPx10_ASAP7_75t_R FILLER_60_974 ();
 DECAPx6_ASAP7_75t_R FILLER_60_996 ();
 FILLER_ASAP7_75t_R FILLER_60_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1063 ();
 FILLER_ASAP7_75t_R FILLER_60_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1079 ();
 FILLER_ASAP7_75t_R FILLER_60_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1088 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1166 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1201 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1215 ();
 FILLER_ASAP7_75t_R FILLER_60_1229 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_61_512 ();
 DECAPx10_ASAP7_75t_R FILLER_61_534 ();
 DECAPx4_ASAP7_75t_R FILLER_61_556 ();
 DECAPx6_ASAP7_75t_R FILLER_61_574 ();
 DECAPx2_ASAP7_75t_R FILLER_61_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_604 ();
 DECAPx10_ASAP7_75t_R FILLER_61_611 ();
 DECAPx10_ASAP7_75t_R FILLER_61_633 ();
 DECAPx1_ASAP7_75t_R FILLER_61_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_659 ();
 DECAPx4_ASAP7_75t_R FILLER_61_678 ();
 FILLER_ASAP7_75t_R FILLER_61_702 ();
 DECAPx6_ASAP7_75t_R FILLER_61_722 ();
 DECAPx1_ASAP7_75t_R FILLER_61_736 ();
 DECAPx10_ASAP7_75t_R FILLER_61_746 ();
 DECAPx1_ASAP7_75t_R FILLER_61_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_772 ();
 DECAPx2_ASAP7_75t_R FILLER_61_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_795 ();
 DECAPx10_ASAP7_75t_R FILLER_61_808 ();
 DECAPx10_ASAP7_75t_R FILLER_61_830 ();
 DECAPx10_ASAP7_75t_R FILLER_61_852 ();
 DECAPx2_ASAP7_75t_R FILLER_61_874 ();
 DECAPx2_ASAP7_75t_R FILLER_61_892 ();
 FILLER_ASAP7_75t_R FILLER_61_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_900 ();
 DECAPx10_ASAP7_75t_R FILLER_61_929 ();
 DECAPx2_ASAP7_75t_R FILLER_61_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_957 ();
 DECAPx10_ASAP7_75t_R FILLER_61_972 ();
 DECAPx2_ASAP7_75t_R FILLER_61_994 ();
 FILLER_ASAP7_75t_R FILLER_61_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1015 ();
 FILLER_ASAP7_75t_R FILLER_61_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1195 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1281 ();
 FILLER_ASAP7_75t_R FILLER_61_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_62_512 ();
 DECAPx10_ASAP7_75t_R FILLER_62_534 ();
 FILLER_ASAP7_75t_R FILLER_62_556 ();
 DECAPx10_ASAP7_75t_R FILLER_62_578 ();
 DECAPx10_ASAP7_75t_R FILLER_62_600 ();
 DECAPx2_ASAP7_75t_R FILLER_62_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_628 ();
 DECAPx2_ASAP7_75t_R FILLER_62_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_651 ();
 DECAPx10_ASAP7_75t_R FILLER_62_659 ();
 DECAPx10_ASAP7_75t_R FILLER_62_681 ();
 DECAPx10_ASAP7_75t_R FILLER_62_703 ();
 DECAPx1_ASAP7_75t_R FILLER_62_725 ();
 DECAPx1_ASAP7_75t_R FILLER_62_739 ();
 DECAPx6_ASAP7_75t_R FILLER_62_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_767 ();
 DECAPx1_ASAP7_75t_R FILLER_62_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_793 ();
 FILLER_ASAP7_75t_R FILLER_62_800 ();
 DECAPx10_ASAP7_75t_R FILLER_62_808 ();
 DECAPx10_ASAP7_75t_R FILLER_62_830 ();
 DECAPx4_ASAP7_75t_R FILLER_62_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_862 ();
 DECAPx10_ASAP7_75t_R FILLER_62_882 ();
 DECAPx10_ASAP7_75t_R FILLER_62_904 ();
 FILLER_ASAP7_75t_R FILLER_62_926 ();
 DECAPx1_ASAP7_75t_R FILLER_62_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_944 ();
 DECAPx4_ASAP7_75t_R FILLER_62_959 ();
 FILLER_ASAP7_75t_R FILLER_62_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_971 ();
 DECAPx2_ASAP7_75t_R FILLER_62_984 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1013 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1046 ();
 FILLER_ASAP7_75t_R FILLER_62_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1060 ();
 FILLER_ASAP7_75t_R FILLER_62_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1122 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1144 ();
 FILLER_ASAP7_75t_R FILLER_62_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1166 ();
 FILLER_ASAP7_75t_R FILLER_62_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1218 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_63_512 ();
 DECAPx10_ASAP7_75t_R FILLER_63_534 ();
 DECAPx10_ASAP7_75t_R FILLER_63_556 ();
 DECAPx2_ASAP7_75t_R FILLER_63_578 ();
 FILLER_ASAP7_75t_R FILLER_63_584 ();
 DECAPx10_ASAP7_75t_R FILLER_63_594 ();
 DECAPx10_ASAP7_75t_R FILLER_63_640 ();
 DECAPx10_ASAP7_75t_R FILLER_63_662 ();
 FILLER_ASAP7_75t_R FILLER_63_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_686 ();
 FILLER_ASAP7_75t_R FILLER_63_693 ();
 FILLER_ASAP7_75t_R FILLER_63_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_725 ();
 DECAPx10_ASAP7_75t_R FILLER_63_732 ();
 DECAPx6_ASAP7_75t_R FILLER_63_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_782 ();
 DECAPx10_ASAP7_75t_R FILLER_63_793 ();
 DECAPx4_ASAP7_75t_R FILLER_63_822 ();
 FILLER_ASAP7_75t_R FILLER_63_838 ();
 DECAPx6_ASAP7_75t_R FILLER_63_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_860 ();
 DECAPx1_ASAP7_75t_R FILLER_63_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_877 ();
 DECAPx10_ASAP7_75t_R FILLER_63_884 ();
 DECAPx10_ASAP7_75t_R FILLER_63_906 ();
 DECAPx1_ASAP7_75t_R FILLER_63_928 ();
 DECAPx2_ASAP7_75t_R FILLER_63_939 ();
 DECAPx6_ASAP7_75t_R FILLER_63_966 ();
 DECAPx2_ASAP7_75t_R FILLER_63_986 ();
 FILLER_ASAP7_75t_R FILLER_63_992 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1027 ();
 FILLER_ASAP7_75t_R FILLER_63_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_63_1103 ();
 FILLER_ASAP7_75t_R FILLER_63_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1115 ();
 FILLER_ASAP7_75t_R FILLER_63_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1148 ();
 FILLER_ASAP7_75t_R FILLER_63_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1252 ();
 DECAPx4_ASAP7_75t_R FILLER_63_1259 ();
 FILLER_ASAP7_75t_R FILLER_63_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_64_512 ();
 DECAPx6_ASAP7_75t_R FILLER_64_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_548 ();
 DECAPx1_ASAP7_75t_R FILLER_64_561 ();
 DECAPx1_ASAP7_75t_R FILLER_64_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_584 ();
 FILLER_ASAP7_75t_R FILLER_64_588 ();
 DECAPx10_ASAP7_75t_R FILLER_64_599 ();
 DECAPx2_ASAP7_75t_R FILLER_64_621 ();
 FILLER_ASAP7_75t_R FILLER_64_627 ();
 DECAPx6_ASAP7_75t_R FILLER_64_647 ();
 FILLER_ASAP7_75t_R FILLER_64_661 ();
 DECAPx6_ASAP7_75t_R FILLER_64_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_688 ();
 FILLER_ASAP7_75t_R FILLER_64_704 ();
 DECAPx2_ASAP7_75t_R FILLER_64_724 ();
 DECAPx10_ASAP7_75t_R FILLER_64_736 ();
 FILLER_ASAP7_75t_R FILLER_64_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_760 ();
 DECAPx10_ASAP7_75t_R FILLER_64_767 ();
 DECAPx10_ASAP7_75t_R FILLER_64_789 ();
 FILLER_ASAP7_75t_R FILLER_64_811 ();
 DECAPx2_ASAP7_75t_R FILLER_64_834 ();
 FILLER_ASAP7_75t_R FILLER_64_840 ();
 DECAPx6_ASAP7_75t_R FILLER_64_848 ();
 DECAPx2_ASAP7_75t_R FILLER_64_862 ();
 DECAPx2_ASAP7_75t_R FILLER_64_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_899 ();
 DECAPx10_ASAP7_75t_R FILLER_64_906 ();
 DECAPx6_ASAP7_75t_R FILLER_64_928 ();
 DECAPx1_ASAP7_75t_R FILLER_64_942 ();
 DECAPx1_ASAP7_75t_R FILLER_64_953 ();
 DECAPx2_ASAP7_75t_R FILLER_64_963 ();
 FILLER_ASAP7_75t_R FILLER_64_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_971 ();
 FILLER_ASAP7_75t_R FILLER_64_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_976 ();
 DECAPx2_ASAP7_75t_R FILLER_64_984 ();
 FILLER_ASAP7_75t_R FILLER_64_996 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1028 ();
 FILLER_ASAP7_75t_R FILLER_64_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1050 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1107 ();
 FILLER_ASAP7_75t_R FILLER_64_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1150 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1195 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_65_512 ();
 DECAPx1_ASAP7_75t_R FILLER_65_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_538 ();
 DECAPx2_ASAP7_75t_R FILLER_65_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_588 ();
 DECAPx4_ASAP7_75t_R FILLER_65_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_623 ();
 DECAPx4_ASAP7_75t_R FILLER_65_629 ();
 FILLER_ASAP7_75t_R FILLER_65_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_641 ();
 DECAPx1_ASAP7_75t_R FILLER_65_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_689 ();
 DECAPx1_ASAP7_75t_R FILLER_65_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_707 ();
 DECAPx6_ASAP7_75t_R FILLER_65_720 ();
 FILLER_ASAP7_75t_R FILLER_65_744 ();
 DECAPx10_ASAP7_75t_R FILLER_65_768 ();
 DECAPx6_ASAP7_75t_R FILLER_65_790 ();
 DECAPx2_ASAP7_75t_R FILLER_65_810 ();
 DECAPx10_ASAP7_75t_R FILLER_65_822 ();
 FILLER_ASAP7_75t_R FILLER_65_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_846 ();
 DECAPx10_ASAP7_75t_R FILLER_65_857 ();
 DECAPx4_ASAP7_75t_R FILLER_65_879 ();
 FILLER_ASAP7_75t_R FILLER_65_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_891 ();
 FILLER_ASAP7_75t_R FILLER_65_898 ();
 FILLER_ASAP7_75t_R FILLER_65_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_916 ();
 DECAPx10_ASAP7_75t_R FILLER_65_952 ();
 DECAPx2_ASAP7_75t_R FILLER_65_974 ();
 DECAPx1_ASAP7_75t_R FILLER_65_995 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1130 ();
 FILLER_ASAP7_75t_R FILLER_65_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1202 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1237 ();
 FILLER_ASAP7_75t_R FILLER_65_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_66_512 ();
 DECAPx10_ASAP7_75t_R FILLER_66_534 ();
 DECAPx10_ASAP7_75t_R FILLER_66_556 ();
 FILLER_ASAP7_75t_R FILLER_66_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_587 ();
 DECAPx10_ASAP7_75t_R FILLER_66_594 ();
 DECAPx6_ASAP7_75t_R FILLER_66_616 ();
 DECAPx1_ASAP7_75t_R FILLER_66_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_634 ();
 DECAPx2_ASAP7_75t_R FILLER_66_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_647 ();
 DECAPx10_ASAP7_75t_R FILLER_66_654 ();
 DECAPx6_ASAP7_75t_R FILLER_66_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_690 ();
 DECAPx4_ASAP7_75t_R FILLER_66_707 ();
 FILLER_ASAP7_75t_R FILLER_66_717 ();
 DECAPx4_ASAP7_75t_R FILLER_66_725 ();
 DECAPx4_ASAP7_75t_R FILLER_66_745 ();
 FILLER_ASAP7_75t_R FILLER_66_755 ();
 DECAPx2_ASAP7_75t_R FILLER_66_763 ();
 FILLER_ASAP7_75t_R FILLER_66_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_771 ();
 FILLER_ASAP7_75t_R FILLER_66_788 ();
 DECAPx6_ASAP7_75t_R FILLER_66_808 ();
 DECAPx2_ASAP7_75t_R FILLER_66_822 ();
 DECAPx10_ASAP7_75t_R FILLER_66_834 ();
 DECAPx6_ASAP7_75t_R FILLER_66_856 ();
 DECAPx1_ASAP7_75t_R FILLER_66_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_874 ();
 DECAPx1_ASAP7_75t_R FILLER_66_881 ();
 FILLER_ASAP7_75t_R FILLER_66_895 ();
 DECAPx6_ASAP7_75t_R FILLER_66_909 ();
 FILLER_ASAP7_75t_R FILLER_66_923 ();
 DECAPx6_ASAP7_75t_R FILLER_66_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_958 ();
 DECAPx1_ASAP7_75t_R FILLER_66_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_971 ();
 DECAPx6_ASAP7_75t_R FILLER_66_974 ();
 DECAPx2_ASAP7_75t_R FILLER_66_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_994 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1077 ();
 FILLER_ASAP7_75t_R FILLER_66_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1167 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1240 ();
 FILLER_ASAP7_75t_R FILLER_66_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1283 ();
 DECAPx4_ASAP7_75t_R FILLER_67_512 ();
 FILLER_ASAP7_75t_R FILLER_67_522 ();
 DECAPx4_ASAP7_75t_R FILLER_67_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_571 ();
 DECAPx10_ASAP7_75t_R FILLER_67_593 ();
 DECAPx6_ASAP7_75t_R FILLER_67_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_629 ();
 DECAPx10_ASAP7_75t_R FILLER_67_643 ();
 DECAPx1_ASAP7_75t_R FILLER_67_665 ();
 DECAPx10_ASAP7_75t_R FILLER_67_703 ();
 DECAPx1_ASAP7_75t_R FILLER_67_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_729 ();
 DECAPx6_ASAP7_75t_R FILLER_67_740 ();
 FILLER_ASAP7_75t_R FILLER_67_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_756 ();
 DECAPx10_ASAP7_75t_R FILLER_67_763 ();
 DECAPx10_ASAP7_75t_R FILLER_67_791 ();
 DECAPx6_ASAP7_75t_R FILLER_67_813 ();
 DECAPx1_ASAP7_75t_R FILLER_67_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_831 ();
 DECAPx10_ASAP7_75t_R FILLER_67_838 ();
 DECAPx10_ASAP7_75t_R FILLER_67_860 ();
 DECAPx10_ASAP7_75t_R FILLER_67_882 ();
 DECAPx1_ASAP7_75t_R FILLER_67_904 ();
 DECAPx2_ASAP7_75t_R FILLER_67_919 ();
 FILLER_ASAP7_75t_R FILLER_67_925 ();
 DECAPx10_ASAP7_75t_R FILLER_67_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_955 ();
 DECAPx10_ASAP7_75t_R FILLER_67_987 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1130 ();
 FILLER_ASAP7_75t_R FILLER_67_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1175 ();
 FILLER_ASAP7_75t_R FILLER_67_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1280 ();
 FILLER_ASAP7_75t_R FILLER_67_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_68_512 ();
 DECAPx2_ASAP7_75t_R FILLER_68_555 ();
 FILLER_ASAP7_75t_R FILLER_68_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_575 ();
 DECAPx10_ASAP7_75t_R FILLER_68_582 ();
 DECAPx10_ASAP7_75t_R FILLER_68_604 ();
 DECAPx4_ASAP7_75t_R FILLER_68_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_636 ();
 DECAPx1_ASAP7_75t_R FILLER_68_657 ();
 FILLER_ASAP7_75t_R FILLER_68_671 ();
 DECAPx2_ASAP7_75t_R FILLER_68_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_695 ();
 DECAPx10_ASAP7_75t_R FILLER_68_710 ();
 FILLER_ASAP7_75t_R FILLER_68_732 ();
 DECAPx4_ASAP7_75t_R FILLER_68_748 ();
 DECAPx10_ASAP7_75t_R FILLER_68_764 ();
 DECAPx10_ASAP7_75t_R FILLER_68_786 ();
 DECAPx10_ASAP7_75t_R FILLER_68_808 ();
 DECAPx10_ASAP7_75t_R FILLER_68_830 ();
 DECAPx10_ASAP7_75t_R FILLER_68_852 ();
 DECAPx10_ASAP7_75t_R FILLER_68_874 ();
 DECAPx10_ASAP7_75t_R FILLER_68_896 ();
 DECAPx10_ASAP7_75t_R FILLER_68_918 ();
 DECAPx10_ASAP7_75t_R FILLER_68_940 ();
 DECAPx4_ASAP7_75t_R FILLER_68_962 ();
 DECAPx10_ASAP7_75t_R FILLER_68_974 ();
 DECAPx10_ASAP7_75t_R FILLER_68_996 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1105 ();
 FILLER_ASAP7_75t_R FILLER_68_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1135 ();
 FILLER_ASAP7_75t_R FILLER_68_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1170 ();
 FILLER_ASAP7_75t_R FILLER_68_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1207 ();
 FILLER_ASAP7_75t_R FILLER_68_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_69_512 ();
 DECAPx10_ASAP7_75t_R FILLER_69_534 ();
 DECAPx1_ASAP7_75t_R FILLER_69_556 ();
 DECAPx10_ASAP7_75t_R FILLER_69_581 ();
 DECAPx10_ASAP7_75t_R FILLER_69_603 ();
 FILLER_ASAP7_75t_R FILLER_69_625 ();
 DECAPx10_ASAP7_75t_R FILLER_69_651 ();
 DECAPx4_ASAP7_75t_R FILLER_69_673 ();
 DECAPx2_ASAP7_75t_R FILLER_69_689 ();
 FILLER_ASAP7_75t_R FILLER_69_695 ();
 DECAPx10_ASAP7_75t_R FILLER_69_717 ();
 DECAPx10_ASAP7_75t_R FILLER_69_739 ();
 DECAPx4_ASAP7_75t_R FILLER_69_761 ();
 FILLER_ASAP7_75t_R FILLER_69_771 ();
 DECAPx6_ASAP7_75t_R FILLER_69_783 ();
 FILLER_ASAP7_75t_R FILLER_69_797 ();
 DECAPx6_ASAP7_75t_R FILLER_69_806 ();
 DECAPx1_ASAP7_75t_R FILLER_69_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_824 ();
 FILLER_ASAP7_75t_R FILLER_69_832 ();
 DECAPx6_ASAP7_75t_R FILLER_69_840 ();
 DECAPx1_ASAP7_75t_R FILLER_69_854 ();
 DECAPx2_ASAP7_75t_R FILLER_69_868 ();
 FILLER_ASAP7_75t_R FILLER_69_874 ();
 DECAPx10_ASAP7_75t_R FILLER_69_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_912 ();
 DECAPx2_ASAP7_75t_R FILLER_69_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_931 ();
 DECAPx10_ASAP7_75t_R FILLER_69_940 ();
 DECAPx10_ASAP7_75t_R FILLER_69_962 ();
 DECAPx10_ASAP7_75t_R FILLER_69_984 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1093 ();
 FILLER_ASAP7_75t_R FILLER_69_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1150 ();
 FILLER_ASAP7_75t_R FILLER_69_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1277 ();
 FILLER_ASAP7_75t_R FILLER_69_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_512 ();
 DECAPx6_ASAP7_75t_R FILLER_70_523 ();
 DECAPx4_ASAP7_75t_R FILLER_70_547 ();
 FILLER_ASAP7_75t_R FILLER_70_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_559 ();
 DECAPx10_ASAP7_75t_R FILLER_70_566 ();
 DECAPx10_ASAP7_75t_R FILLER_70_588 ();
 DECAPx4_ASAP7_75t_R FILLER_70_610 ();
 DECAPx10_ASAP7_75t_R FILLER_70_654 ();
 DECAPx10_ASAP7_75t_R FILLER_70_676 ();
 DECAPx1_ASAP7_75t_R FILLER_70_698 ();
 DECAPx4_ASAP7_75t_R FILLER_70_753 ();
 FILLER_ASAP7_75t_R FILLER_70_763 ();
 DECAPx10_ASAP7_75t_R FILLER_70_775 ();
 FILLER_ASAP7_75t_R FILLER_70_797 ();
 DECAPx6_ASAP7_75t_R FILLER_70_815 ();
 DECAPx2_ASAP7_75t_R FILLER_70_840 ();
 FILLER_ASAP7_75t_R FILLER_70_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_865 ();
 DECAPx1_ASAP7_75t_R FILLER_70_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_876 ();
 DECAPx1_ASAP7_75t_R FILLER_70_883 ();
 DECAPx10_ASAP7_75t_R FILLER_70_917 ();
 FILLER_ASAP7_75t_R FILLER_70_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_941 ();
 FILLER_ASAP7_75t_R FILLER_70_949 ();
 DECAPx10_ASAP7_75t_R FILLER_70_974 ();
 DECAPx2_ASAP7_75t_R FILLER_70_996 ();
 FILLER_ASAP7_75t_R FILLER_70_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1134 ();
 FILLER_ASAP7_75t_R FILLER_70_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1180 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1208 ();
 FILLER_ASAP7_75t_R FILLER_70_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1241 ();
 FILLER_ASAP7_75t_R FILLER_70_1247 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1255 ();
 FILLER_ASAP7_75t_R FILLER_70_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_71_512 ();
 DECAPx4_ASAP7_75t_R FILLER_71_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_544 ();
 DECAPx2_ASAP7_75t_R FILLER_71_551 ();
 DECAPx4_ASAP7_75t_R FILLER_71_563 ();
 FILLER_ASAP7_75t_R FILLER_71_573 ();
 DECAPx10_ASAP7_75t_R FILLER_71_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_618 ();
 DECAPx6_ASAP7_75t_R FILLER_71_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_651 ();
 DECAPx10_ASAP7_75t_R FILLER_71_662 ();
 DECAPx6_ASAP7_75t_R FILLER_71_684 ();
 DECAPx1_ASAP7_75t_R FILLER_71_698 ();
 DECAPx4_ASAP7_75t_R FILLER_71_732 ();
 FILLER_ASAP7_75t_R FILLER_71_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_756 ();
 DECAPx2_ASAP7_75t_R FILLER_71_764 ();
 FILLER_ASAP7_75t_R FILLER_71_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_772 ();
 FILLER_ASAP7_75t_R FILLER_71_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_785 ();
 DECAPx10_ASAP7_75t_R FILLER_71_794 ();
 DECAPx10_ASAP7_75t_R FILLER_71_816 ();
 DECAPx10_ASAP7_75t_R FILLER_71_838 ();
 DECAPx10_ASAP7_75t_R FILLER_71_860 ();
 DECAPx10_ASAP7_75t_R FILLER_71_882 ();
 DECAPx10_ASAP7_75t_R FILLER_71_904 ();
 DECAPx1_ASAP7_75t_R FILLER_71_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_930 ();
 DECAPx6_ASAP7_75t_R FILLER_71_973 ();
 FILLER_ASAP7_75t_R FILLER_71_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_989 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1004 ();
 FILLER_ASAP7_75t_R FILLER_71_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1035 ();
 FILLER_ASAP7_75t_R FILLER_71_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1055 ();
 FILLER_ASAP7_75t_R FILLER_71_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1127 ();
 FILLER_ASAP7_75t_R FILLER_71_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1151 ();
 FILLER_ASAP7_75t_R FILLER_71_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_72_512 ();
 FILLER_ASAP7_75t_R FILLER_72_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_524 ();
 DECAPx2_ASAP7_75t_R FILLER_72_564 ();
 FILLER_ASAP7_75t_R FILLER_72_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_572 ();
 DECAPx10_ASAP7_75t_R FILLER_72_581 ();
 DECAPx10_ASAP7_75t_R FILLER_72_603 ();
 DECAPx1_ASAP7_75t_R FILLER_72_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_629 ();
 DECAPx2_ASAP7_75t_R FILLER_72_636 ();
 FILLER_ASAP7_75t_R FILLER_72_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_668 ();
 DECAPx2_ASAP7_75t_R FILLER_72_699 ();
 DECAPx4_ASAP7_75t_R FILLER_72_712 ();
 DECAPx10_ASAP7_75t_R FILLER_72_729 ();
 DECAPx2_ASAP7_75t_R FILLER_72_751 ();
 FILLER_ASAP7_75t_R FILLER_72_757 ();
 DECAPx2_ASAP7_75t_R FILLER_72_775 ();
 FILLER_ASAP7_75t_R FILLER_72_781 ();
 DECAPx10_ASAP7_75t_R FILLER_72_789 ();
 DECAPx10_ASAP7_75t_R FILLER_72_811 ();
 DECAPx10_ASAP7_75t_R FILLER_72_833 ();
 DECAPx10_ASAP7_75t_R FILLER_72_855 ();
 DECAPx10_ASAP7_75t_R FILLER_72_877 ();
 DECAPx4_ASAP7_75t_R FILLER_72_899 ();
 DECAPx2_ASAP7_75t_R FILLER_72_915 ();
 FILLER_ASAP7_75t_R FILLER_72_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_923 ();
 DECAPx4_ASAP7_75t_R FILLER_72_934 ();
 DECAPx10_ASAP7_75t_R FILLER_72_950 ();
 DECAPx10_ASAP7_75t_R FILLER_72_974 ();
 DECAPx6_ASAP7_75t_R FILLER_72_996 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1076 ();
 FILLER_ASAP7_75t_R FILLER_72_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1092 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_73_512 ();
 DECAPx10_ASAP7_75t_R FILLER_73_534 ();
 DECAPx1_ASAP7_75t_R FILLER_73_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_560 ();
 DECAPx2_ASAP7_75t_R FILLER_73_582 ();
 FILLER_ASAP7_75t_R FILLER_73_588 ();
 DECAPx10_ASAP7_75t_R FILLER_73_596 ();
 DECAPx10_ASAP7_75t_R FILLER_73_618 ();
 DECAPx10_ASAP7_75t_R FILLER_73_658 ();
 DECAPx10_ASAP7_75t_R FILLER_73_680 ();
 DECAPx10_ASAP7_75t_R FILLER_73_702 ();
 DECAPx6_ASAP7_75t_R FILLER_73_724 ();
 DECAPx1_ASAP7_75t_R FILLER_73_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_742 ();
 DECAPx10_ASAP7_75t_R FILLER_73_746 ();
 DECAPx10_ASAP7_75t_R FILLER_73_768 ();
 DECAPx10_ASAP7_75t_R FILLER_73_790 ();
 DECAPx10_ASAP7_75t_R FILLER_73_812 ();
 DECAPx6_ASAP7_75t_R FILLER_73_834 ();
 FILLER_ASAP7_75t_R FILLER_73_848 ();
 DECAPx4_ASAP7_75t_R FILLER_73_858 ();
 FILLER_ASAP7_75t_R FILLER_73_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_870 ();
 DECAPx10_ASAP7_75t_R FILLER_73_893 ();
 DECAPx4_ASAP7_75t_R FILLER_73_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_925 ();
 DECAPx2_ASAP7_75t_R FILLER_73_956 ();
 FILLER_ASAP7_75t_R FILLER_73_962 ();
 DECAPx6_ASAP7_75t_R FILLER_73_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_996 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1007 ();
 FILLER_ASAP7_75t_R FILLER_73_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1139 ();
 FILLER_ASAP7_75t_R FILLER_73_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1175 ();
 FILLER_ASAP7_75t_R FILLER_73_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1201 ();
 FILLER_ASAP7_75t_R FILLER_73_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1216 ();
 FILLER_ASAP7_75t_R FILLER_73_1225 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1242 ();
 FILLER_ASAP7_75t_R FILLER_73_1252 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1281 ();
 FILLER_ASAP7_75t_R FILLER_73_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_74_512 ();
 DECAPx6_ASAP7_75t_R FILLER_74_534 ();
 DECAPx1_ASAP7_75t_R FILLER_74_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_560 ();
 DECAPx10_ASAP7_75t_R FILLER_74_575 ();
 DECAPx6_ASAP7_75t_R FILLER_74_597 ();
 DECAPx2_ASAP7_75t_R FILLER_74_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_633 ();
 DECAPx2_ASAP7_75t_R FILLER_74_644 ();
 FILLER_ASAP7_75t_R FILLER_74_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_652 ();
 DECAPx2_ASAP7_75t_R FILLER_74_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_677 ();
 FILLER_ASAP7_75t_R FILLER_74_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_709 ();
 DECAPx1_ASAP7_75t_R FILLER_74_716 ();
 DECAPx4_ASAP7_75t_R FILLER_74_726 ();
 FILLER_ASAP7_75t_R FILLER_74_736 ();
 DECAPx6_ASAP7_75t_R FILLER_74_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_773 ();
 DECAPx6_ASAP7_75t_R FILLER_74_780 ();
 DECAPx2_ASAP7_75t_R FILLER_74_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_800 ();
 DECAPx4_ASAP7_75t_R FILLER_74_813 ();
 FILLER_ASAP7_75t_R FILLER_74_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_825 ();
 DECAPx10_ASAP7_75t_R FILLER_74_838 ();
 DECAPx10_ASAP7_75t_R FILLER_74_860 ();
 DECAPx2_ASAP7_75t_R FILLER_74_882 ();
 DECAPx10_ASAP7_75t_R FILLER_74_894 ();
 DECAPx2_ASAP7_75t_R FILLER_74_916 ();
 DECAPx2_ASAP7_75t_R FILLER_74_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_937 ();
 DECAPx2_ASAP7_75t_R FILLER_74_952 ();
 DECAPx10_ASAP7_75t_R FILLER_74_974 ();
 DECAPx10_ASAP7_75t_R FILLER_74_996 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1018 ();
 FILLER_ASAP7_75t_R FILLER_74_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1071 ();
 FILLER_ASAP7_75t_R FILLER_74_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1161 ();
 FILLER_ASAP7_75t_R FILLER_74_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1190 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1232 ();
 DECAPx6_ASAP7_75t_R FILLER_75_512 ();
 FILLER_ASAP7_75t_R FILLER_75_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_528 ();
 DECAPx2_ASAP7_75t_R FILLER_75_551 ();
 DECAPx10_ASAP7_75t_R FILLER_75_563 ();
 DECAPx10_ASAP7_75t_R FILLER_75_585 ();
 DECAPx4_ASAP7_75t_R FILLER_75_607 ();
 FILLER_ASAP7_75t_R FILLER_75_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_626 ();
 DECAPx10_ASAP7_75t_R FILLER_75_645 ();
 DECAPx6_ASAP7_75t_R FILLER_75_667 ();
 DECAPx10_ASAP7_75t_R FILLER_75_697 ();
 DECAPx1_ASAP7_75t_R FILLER_75_719 ();
 DECAPx10_ASAP7_75t_R FILLER_75_733 ();
 DECAPx6_ASAP7_75t_R FILLER_75_755 ();
 DECAPx2_ASAP7_75t_R FILLER_75_769 ();
 DECAPx6_ASAP7_75t_R FILLER_75_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_795 ();
 DECAPx10_ASAP7_75t_R FILLER_75_802 ();
 DECAPx10_ASAP7_75t_R FILLER_75_824 ();
 DECAPx6_ASAP7_75t_R FILLER_75_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_860 ();
 DECAPx10_ASAP7_75t_R FILLER_75_867 ();
 DECAPx4_ASAP7_75t_R FILLER_75_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_899 ();
 DECAPx10_ASAP7_75t_R FILLER_75_914 ();
 DECAPx6_ASAP7_75t_R FILLER_75_936 ();
 DECAPx1_ASAP7_75t_R FILLER_75_950 ();
 DECAPx10_ASAP7_75t_R FILLER_75_964 ();
 DECAPx1_ASAP7_75t_R FILLER_75_986 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1058 ();
 FILLER_ASAP7_75t_R FILLER_75_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1096 ();
 FILLER_ASAP7_75t_R FILLER_75_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1132 ();
 FILLER_ASAP7_75t_R FILLER_75_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1181 ();
 FILLER_ASAP7_75t_R FILLER_75_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_76_512 ();
 DECAPx6_ASAP7_75t_R FILLER_76_534 ();
 FILLER_ASAP7_75t_R FILLER_76_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_550 ();
 DECAPx4_ASAP7_75t_R FILLER_76_559 ();
 FILLER_ASAP7_75t_R FILLER_76_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_571 ();
 DECAPx6_ASAP7_75t_R FILLER_76_598 ();
 DECAPx1_ASAP7_75t_R FILLER_76_612 ();
 DECAPx6_ASAP7_75t_R FILLER_76_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_652 ();
 FILLER_ASAP7_75t_R FILLER_76_659 ();
 DECAPx1_ASAP7_75t_R FILLER_76_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_671 ();
 DECAPx10_ASAP7_75t_R FILLER_76_681 ();
 DECAPx1_ASAP7_75t_R FILLER_76_703 ();
 DECAPx6_ASAP7_75t_R FILLER_76_733 ();
 DECAPx4_ASAP7_75t_R FILLER_76_765 ();
 FILLER_ASAP7_75t_R FILLER_76_775 ();
 DECAPx6_ASAP7_75t_R FILLER_76_783 ();
 DECAPx10_ASAP7_75t_R FILLER_76_803 ();
 DECAPx10_ASAP7_75t_R FILLER_76_825 ();
 DECAPx4_ASAP7_75t_R FILLER_76_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_857 ();
 DECAPx10_ASAP7_75t_R FILLER_76_886 ();
 DECAPx10_ASAP7_75t_R FILLER_76_908 ();
 DECAPx10_ASAP7_75t_R FILLER_76_930 ();
 DECAPx6_ASAP7_75t_R FILLER_76_952 ();
 DECAPx2_ASAP7_75t_R FILLER_76_966 ();
 DECAPx10_ASAP7_75t_R FILLER_76_974 ();
 DECAPx10_ASAP7_75t_R FILLER_76_996 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1065 ();
 FILLER_ASAP7_75t_R FILLER_76_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1136 ();
 FILLER_ASAP7_75t_R FILLER_76_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1161 ();
 FILLER_ASAP7_75t_R FILLER_76_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1181 ();
 FILLER_ASAP7_75t_R FILLER_76_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1244 ();
 FILLER_ASAP7_75t_R FILLER_76_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_77_512 ();
 FILLER_ASAP7_75t_R FILLER_77_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_546 ();
 DECAPx10_ASAP7_75t_R FILLER_77_568 ();
 DECAPx10_ASAP7_75t_R FILLER_77_590 ();
 DECAPx4_ASAP7_75t_R FILLER_77_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_622 ();
 DECAPx4_ASAP7_75t_R FILLER_77_639 ();
 DECAPx2_ASAP7_75t_R FILLER_77_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_668 ();
 DECAPx6_ASAP7_75t_R FILLER_77_676 ();
 FILLER_ASAP7_75t_R FILLER_77_690 ();
 DECAPx4_ASAP7_75t_R FILLER_77_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_710 ();
 DECAPx6_ASAP7_75t_R FILLER_77_746 ();
 DECAPx2_ASAP7_75t_R FILLER_77_766 ();
 FILLER_ASAP7_75t_R FILLER_77_772 ();
 DECAPx10_ASAP7_75t_R FILLER_77_786 ();
 DECAPx10_ASAP7_75t_R FILLER_77_808 ();
 DECAPx6_ASAP7_75t_R FILLER_77_830 ();
 DECAPx2_ASAP7_75t_R FILLER_77_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_850 ();
 DECAPx2_ASAP7_75t_R FILLER_77_861 ();
 FILLER_ASAP7_75t_R FILLER_77_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_869 ();
 DECAPx10_ASAP7_75t_R FILLER_77_886 ();
 DECAPx6_ASAP7_75t_R FILLER_77_908 ();
 FILLER_ASAP7_75t_R FILLER_77_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_924 ();
 DECAPx4_ASAP7_75t_R FILLER_77_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_963 ();
 DECAPx2_ASAP7_75t_R FILLER_77_974 ();
 FILLER_ASAP7_75t_R FILLER_77_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_982 ();
 DECAPx2_ASAP7_75t_R FILLER_77_993 ();
 FILLER_ASAP7_75t_R FILLER_77_999 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1037 ();
 FILLER_ASAP7_75t_R FILLER_77_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1081 ();
 FILLER_ASAP7_75t_R FILLER_77_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1136 ();
 FILLER_ASAP7_75t_R FILLER_77_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1162 ();
 FILLER_ASAP7_75t_R FILLER_77_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1179 ();
 FILLER_ASAP7_75t_R FILLER_77_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_78_512 ();
 DECAPx4_ASAP7_75t_R FILLER_78_534 ();
 FILLER_ASAP7_75t_R FILLER_78_544 ();
 DECAPx1_ASAP7_75t_R FILLER_78_554 ();
 DECAPx10_ASAP7_75t_R FILLER_78_566 ();
 DECAPx10_ASAP7_75t_R FILLER_78_588 ();
 DECAPx10_ASAP7_75t_R FILLER_78_610 ();
 DECAPx2_ASAP7_75t_R FILLER_78_632 ();
 FILLER_ASAP7_75t_R FILLER_78_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_640 ();
 DECAPx10_ASAP7_75t_R FILLER_78_663 ();
 DECAPx10_ASAP7_75t_R FILLER_78_685 ();
 DECAPx1_ASAP7_75t_R FILLER_78_707 ();
 FILLER_ASAP7_75t_R FILLER_78_735 ();
 DECAPx2_ASAP7_75t_R FILLER_78_743 ();
 FILLER_ASAP7_75t_R FILLER_78_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_751 ();
 DECAPx4_ASAP7_75t_R FILLER_78_758 ();
 FILLER_ASAP7_75t_R FILLER_78_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_770 ();
 DECAPx6_ASAP7_75t_R FILLER_78_787 ();
 FILLER_ASAP7_75t_R FILLER_78_801 ();
 DECAPx1_ASAP7_75t_R FILLER_78_820 ();
 DECAPx6_ASAP7_75t_R FILLER_78_830 ();
 DECAPx2_ASAP7_75t_R FILLER_78_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_850 ();
 DECAPx1_ASAP7_75t_R FILLER_78_867 ();
 DECAPx10_ASAP7_75t_R FILLER_78_899 ();
 FILLER_ASAP7_75t_R FILLER_78_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_923 ();
 DECAPx10_ASAP7_75t_R FILLER_78_942 ();
 DECAPx2_ASAP7_75t_R FILLER_78_964 ();
 FILLER_ASAP7_75t_R FILLER_78_970 ();
 DECAPx10_ASAP7_75t_R FILLER_78_974 ();
 DECAPx2_ASAP7_75t_R FILLER_78_996 ();
 DECAPx4_ASAP7_75t_R FILLER_78_1018 ();
 FILLER_ASAP7_75t_R FILLER_78_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1059 ();
 FILLER_ASAP7_75t_R FILLER_78_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1091 ();
 FILLER_ASAP7_75t_R FILLER_78_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1200 ();
 FILLER_ASAP7_75t_R FILLER_78_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1243 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1276 ();
 FILLER_ASAP7_75t_R FILLER_78_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_79_512 ();
 FILLER_ASAP7_75t_R FILLER_79_526 ();
 DECAPx2_ASAP7_75t_R FILLER_79_538 ();
 DECAPx2_ASAP7_75t_R FILLER_79_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_556 ();
 FILLER_ASAP7_75t_R FILLER_79_578 ();
 DECAPx10_ASAP7_75t_R FILLER_79_588 ();
 DECAPx6_ASAP7_75t_R FILLER_79_610 ();
 DECAPx2_ASAP7_75t_R FILLER_79_624 ();
 DECAPx10_ASAP7_75t_R FILLER_79_654 ();
 DECAPx10_ASAP7_75t_R FILLER_79_676 ();
 DECAPx10_ASAP7_75t_R FILLER_79_698 ();
 DECAPx2_ASAP7_75t_R FILLER_79_720 ();
 DECAPx6_ASAP7_75t_R FILLER_79_746 ();
 FILLER_ASAP7_75t_R FILLER_79_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_762 ();
 FILLER_ASAP7_75t_R FILLER_79_775 ();
 DECAPx10_ASAP7_75t_R FILLER_79_783 ();
 FILLER_ASAP7_75t_R FILLER_79_805 ();
 DECAPx10_ASAP7_75t_R FILLER_79_834 ();
 DECAPx10_ASAP7_75t_R FILLER_79_856 ();
 DECAPx6_ASAP7_75t_R FILLER_79_878 ();
 DECAPx10_ASAP7_75t_R FILLER_79_898 ();
 DECAPx2_ASAP7_75t_R FILLER_79_920 ();
 FILLER_ASAP7_75t_R FILLER_79_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_928 ();
 DECAPx10_ASAP7_75t_R FILLER_79_937 ();
 DECAPx4_ASAP7_75t_R FILLER_79_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_969 ();
 DECAPx6_ASAP7_75t_R FILLER_79_988 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1016 ();
 FILLER_ASAP7_75t_R FILLER_79_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1039 ();
 FILLER_ASAP7_75t_R FILLER_79_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1225 ();
 FILLER_ASAP7_75t_R FILLER_79_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1277 ();
 FILLER_ASAP7_75t_R FILLER_79_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_80_512 ();
 DECAPx2_ASAP7_75t_R FILLER_80_534 ();
 FILLER_ASAP7_75t_R FILLER_80_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_542 ();
 DECAPx4_ASAP7_75t_R FILLER_80_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_569 ();
 DECAPx6_ASAP7_75t_R FILLER_80_576 ();
 DECAPx2_ASAP7_75t_R FILLER_80_590 ();
 DECAPx6_ASAP7_75t_R FILLER_80_602 ();
 FILLER_ASAP7_75t_R FILLER_80_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_618 ();
 DECAPx4_ASAP7_75t_R FILLER_80_635 ();
 FILLER_ASAP7_75t_R FILLER_80_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_647 ();
 FILLER_ASAP7_75t_R FILLER_80_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_660 ();
 DECAPx4_ASAP7_75t_R FILLER_80_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_677 ();
 DECAPx10_ASAP7_75t_R FILLER_80_690 ();
 DECAPx4_ASAP7_75t_R FILLER_80_712 ();
 DECAPx10_ASAP7_75t_R FILLER_80_736 ();
 DECAPx2_ASAP7_75t_R FILLER_80_758 ();
 FILLER_ASAP7_75t_R FILLER_80_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_766 ();
 DECAPx10_ASAP7_75t_R FILLER_80_785 ();
 DECAPx10_ASAP7_75t_R FILLER_80_807 ();
 DECAPx6_ASAP7_75t_R FILLER_80_829 ();
 DECAPx2_ASAP7_75t_R FILLER_80_843 ();
 DECAPx6_ASAP7_75t_R FILLER_80_867 ();
 DECAPx10_ASAP7_75t_R FILLER_80_892 ();
 DECAPx6_ASAP7_75t_R FILLER_80_914 ();
 FILLER_ASAP7_75t_R FILLER_80_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_930 ();
 DECAPx2_ASAP7_75t_R FILLER_80_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_943 ();
 DECAPx6_ASAP7_75t_R FILLER_80_958 ();
 DECAPx10_ASAP7_75t_R FILLER_80_974 ();
 DECAPx6_ASAP7_75t_R FILLER_80_996 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1042 ();
 FILLER_ASAP7_75t_R FILLER_80_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1109 ();
 FILLER_ASAP7_75t_R FILLER_80_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1213 ();
 FILLER_ASAP7_75t_R FILLER_80_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1245 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_81_512 ();
 FILLER_ASAP7_75t_R FILLER_81_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_524 ();
 DECAPx6_ASAP7_75t_R FILLER_81_567 ();
 DECAPx10_ASAP7_75t_R FILLER_81_602 ();
 DECAPx2_ASAP7_75t_R FILLER_81_624 ();
 DECAPx10_ASAP7_75t_R FILLER_81_636 ();
 FILLER_ASAP7_75t_R FILLER_81_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_679 ();
 FILLER_ASAP7_75t_R FILLER_81_686 ();
 DECAPx10_ASAP7_75t_R FILLER_81_694 ();
 DECAPx1_ASAP7_75t_R FILLER_81_716 ();
 DECAPx2_ASAP7_75t_R FILLER_81_745 ();
 FILLER_ASAP7_75t_R FILLER_81_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_753 ();
 DECAPx10_ASAP7_75t_R FILLER_81_761 ();
 DECAPx10_ASAP7_75t_R FILLER_81_783 ();
 DECAPx6_ASAP7_75t_R FILLER_81_805 ();
 DECAPx10_ASAP7_75t_R FILLER_81_835 ();
 DECAPx10_ASAP7_75t_R FILLER_81_857 ();
 DECAPx10_ASAP7_75t_R FILLER_81_879 ();
 DECAPx10_ASAP7_75t_R FILLER_81_901 ();
 DECAPx10_ASAP7_75t_R FILLER_81_923 ();
 DECAPx10_ASAP7_75t_R FILLER_81_945 ();
 DECAPx10_ASAP7_75t_R FILLER_81_967 ();
 DECAPx6_ASAP7_75t_R FILLER_81_989 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1150 ();
 FILLER_ASAP7_75t_R FILLER_81_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1251 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1281 ();
 FILLER_ASAP7_75t_R FILLER_81_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_82_512 ();
 DECAPx6_ASAP7_75t_R FILLER_82_534 ();
 DECAPx1_ASAP7_75t_R FILLER_82_548 ();
 DECAPx4_ASAP7_75t_R FILLER_82_558 ();
 FILLER_ASAP7_75t_R FILLER_82_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_570 ();
 DECAPx10_ASAP7_75t_R FILLER_82_581 ();
 DECAPx1_ASAP7_75t_R FILLER_82_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_607 ();
 DECAPx10_ASAP7_75t_R FILLER_82_630 ();
 DECAPx10_ASAP7_75t_R FILLER_82_652 ();
 DECAPx10_ASAP7_75t_R FILLER_82_674 ();
 DECAPx10_ASAP7_75t_R FILLER_82_696 ();
 DECAPx2_ASAP7_75t_R FILLER_82_718 ();
 FILLER_ASAP7_75t_R FILLER_82_724 ();
 DECAPx10_ASAP7_75t_R FILLER_82_768 ();
 DECAPx2_ASAP7_75t_R FILLER_82_790 ();
 DECAPx10_ASAP7_75t_R FILLER_82_809 ();
 DECAPx4_ASAP7_75t_R FILLER_82_831 ();
 FILLER_ASAP7_75t_R FILLER_82_841 ();
 DECAPx6_ASAP7_75t_R FILLER_82_853 ();
 DECAPx1_ASAP7_75t_R FILLER_82_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_885 ();
 DECAPx10_ASAP7_75t_R FILLER_82_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_918 ();
 DECAPx2_ASAP7_75t_R FILLER_82_937 ();
 FILLER_ASAP7_75t_R FILLER_82_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_952 ();
 DECAPx4_ASAP7_75t_R FILLER_82_959 ();
 FILLER_ASAP7_75t_R FILLER_82_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_971 ();
 DECAPx6_ASAP7_75t_R FILLER_82_974 ();
 DECAPx1_ASAP7_75t_R FILLER_82_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1041 ();
 FILLER_ASAP7_75t_R FILLER_82_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1111 ();
 DECAPx4_ASAP7_75t_R FILLER_82_1133 ();
 FILLER_ASAP7_75t_R FILLER_82_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1200 ();
 FILLER_ASAP7_75t_R FILLER_82_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1260 ();
 FILLER_ASAP7_75t_R FILLER_82_1291 ();
 DECAPx4_ASAP7_75t_R FILLER_83_512 ();
 DECAPx1_ASAP7_75t_R FILLER_83_557 ();
 DECAPx4_ASAP7_75t_R FILLER_83_569 ();
 FILLER_ASAP7_75t_R FILLER_83_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_581 ();
 DECAPx2_ASAP7_75t_R FILLER_83_603 ();
 FILLER_ASAP7_75t_R FILLER_83_609 ();
 DECAPx10_ASAP7_75t_R FILLER_83_633 ();
 DECAPx4_ASAP7_75t_R FILLER_83_655 ();
 DECAPx1_ASAP7_75t_R FILLER_83_681 ();
 DECAPx10_ASAP7_75t_R FILLER_83_699 ();
 DECAPx6_ASAP7_75t_R FILLER_83_721 ();
 DECAPx1_ASAP7_75t_R FILLER_83_735 ();
 DECAPx10_ASAP7_75t_R FILLER_83_745 ();
 DECAPx10_ASAP7_75t_R FILLER_83_767 ();
 DECAPx1_ASAP7_75t_R FILLER_83_789 ();
 DECAPx1_ASAP7_75t_R FILLER_83_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_818 ();
 DECAPx10_ASAP7_75t_R FILLER_83_831 ();
 DECAPx6_ASAP7_75t_R FILLER_83_853 ();
 FILLER_ASAP7_75t_R FILLER_83_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_869 ();
 DECAPx4_ASAP7_75t_R FILLER_83_884 ();
 DECAPx10_ASAP7_75t_R FILLER_83_900 ();
 DECAPx6_ASAP7_75t_R FILLER_83_922 ();
 DECAPx2_ASAP7_75t_R FILLER_83_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_942 ();
 DECAPx4_ASAP7_75t_R FILLER_83_964 ();
 FILLER_ASAP7_75t_R FILLER_83_974 ();
 DECAPx6_ASAP7_75t_R FILLER_83_988 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1140 ();
 FILLER_ASAP7_75t_R FILLER_83_1146 ();
 FILLER_ASAP7_75t_R FILLER_83_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1242 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1276 ();
 FILLER_ASAP7_75t_R FILLER_83_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_84_512 ();
 DECAPx1_ASAP7_75t_R FILLER_84_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_538 ();
 FILLER_ASAP7_75t_R FILLER_84_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_568 ();
 DECAPx4_ASAP7_75t_R FILLER_84_575 ();
 DECAPx2_ASAP7_75t_R FILLER_84_593 ();
 DECAPx6_ASAP7_75t_R FILLER_84_605 ();
 DECAPx2_ASAP7_75t_R FILLER_84_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_625 ();
 DECAPx4_ASAP7_75t_R FILLER_84_632 ();
 DECAPx10_ASAP7_75t_R FILLER_84_648 ();
 DECAPx10_ASAP7_75t_R FILLER_84_670 ();
 DECAPx10_ASAP7_75t_R FILLER_84_692 ();
 DECAPx10_ASAP7_75t_R FILLER_84_714 ();
 DECAPx6_ASAP7_75t_R FILLER_84_736 ();
 DECAPx2_ASAP7_75t_R FILLER_84_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_756 ();
 DECAPx6_ASAP7_75t_R FILLER_84_763 ();
 DECAPx6_ASAP7_75t_R FILLER_84_787 ();
 DECAPx4_ASAP7_75t_R FILLER_84_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_817 ();
 DECAPx10_ASAP7_75t_R FILLER_84_824 ();
 FILLER_ASAP7_75t_R FILLER_84_846 ();
 DECAPx10_ASAP7_75t_R FILLER_84_862 ();
 FILLER_ASAP7_75t_R FILLER_84_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_886 ();
 DECAPx10_ASAP7_75t_R FILLER_84_917 ();
 DECAPx1_ASAP7_75t_R FILLER_84_939 ();
 DECAPx10_ASAP7_75t_R FILLER_84_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_971 ();
 DECAPx2_ASAP7_75t_R FILLER_84_974 ();
 FILLER_ASAP7_75t_R FILLER_84_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_982 ();
 DECAPx10_ASAP7_75t_R FILLER_84_999 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1131 ();
 FILLER_ASAP7_75t_R FILLER_84_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1140 ();
 FILLER_ASAP7_75t_R FILLER_84_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1159 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1166 ();
 FILLER_ASAP7_75t_R FILLER_84_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1269 ();
 FILLER_ASAP7_75t_R FILLER_84_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_85_512 ();
 DECAPx1_ASAP7_75t_R FILLER_85_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_530 ();
 DECAPx4_ASAP7_75t_R FILLER_85_539 ();
 FILLER_ASAP7_75t_R FILLER_85_549 ();
 DECAPx1_ASAP7_75t_R FILLER_85_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_591 ();
 DECAPx10_ASAP7_75t_R FILLER_85_600 ();
 DECAPx10_ASAP7_75t_R FILLER_85_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_644 ();
 DECAPx2_ASAP7_75t_R FILLER_85_655 ();
 FILLER_ASAP7_75t_R FILLER_85_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_663 ();
 DECAPx4_ASAP7_75t_R FILLER_85_697 ();
 FILLER_ASAP7_75t_R FILLER_85_707 ();
 DECAPx4_ASAP7_75t_R FILLER_85_715 ();
 FILLER_ASAP7_75t_R FILLER_85_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_727 ();
 DECAPx10_ASAP7_75t_R FILLER_85_734 ();
 DECAPx2_ASAP7_75t_R FILLER_85_756 ();
 FILLER_ASAP7_75t_R FILLER_85_762 ();
 DECAPx10_ASAP7_75t_R FILLER_85_770 ();
 FILLER_ASAP7_75t_R FILLER_85_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_794 ();
 DECAPx2_ASAP7_75t_R FILLER_85_803 ();
 DECAPx10_ASAP7_75t_R FILLER_85_816 ();
 DECAPx10_ASAP7_75t_R FILLER_85_838 ();
 DECAPx10_ASAP7_75t_R FILLER_85_860 ();
 DECAPx10_ASAP7_75t_R FILLER_85_882 ();
 DECAPx10_ASAP7_75t_R FILLER_85_904 ();
 DECAPx4_ASAP7_75t_R FILLER_85_926 ();
 FILLER_ASAP7_75t_R FILLER_85_936 ();
 DECAPx6_ASAP7_75t_R FILLER_85_944 ();
 DECAPx10_ASAP7_75t_R FILLER_85_968 ();
 DECAPx10_ASAP7_75t_R FILLER_85_990 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1084 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1159 ();
 FILLER_ASAP7_75t_R FILLER_85_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1245 ();
 FILLER_ASAP7_75t_R FILLER_85_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_86_512 ();
 DECAPx6_ASAP7_75t_R FILLER_86_534 ();
 FILLER_ASAP7_75t_R FILLER_86_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_550 ();
 FILLER_ASAP7_75t_R FILLER_86_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_566 ();
 DECAPx10_ASAP7_75t_R FILLER_86_588 ();
 DECAPx6_ASAP7_75t_R FILLER_86_610 ();
 DECAPx1_ASAP7_75t_R FILLER_86_624 ();
 DECAPx4_ASAP7_75t_R FILLER_86_646 ();
 DECAPx4_ASAP7_75t_R FILLER_86_662 ();
 DECAPx2_ASAP7_75t_R FILLER_86_678 ();
 FILLER_ASAP7_75t_R FILLER_86_684 ();
 DECAPx1_ASAP7_75t_R FILLER_86_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_696 ();
 DECAPx2_ASAP7_75t_R FILLER_86_703 ();
 DECAPx2_ASAP7_75t_R FILLER_86_719 ();
 FILLER_ASAP7_75t_R FILLER_86_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_727 ();
 DECAPx10_ASAP7_75t_R FILLER_86_734 ();
 DECAPx1_ASAP7_75t_R FILLER_86_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_760 ();
 DECAPx10_ASAP7_75t_R FILLER_86_767 ();
 DECAPx6_ASAP7_75t_R FILLER_86_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_803 ();
 FILLER_ASAP7_75t_R FILLER_86_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_819 ();
 DECAPx10_ASAP7_75t_R FILLER_86_832 ();
 DECAPx10_ASAP7_75t_R FILLER_86_854 ();
 DECAPx10_ASAP7_75t_R FILLER_86_876 ();
 DECAPx4_ASAP7_75t_R FILLER_86_907 ();
 FILLER_ASAP7_75t_R FILLER_86_917 ();
 DECAPx10_ASAP7_75t_R FILLER_86_940 ();
 DECAPx4_ASAP7_75t_R FILLER_86_962 ();
 DECAPx10_ASAP7_75t_R FILLER_86_974 ();
 DECAPx10_ASAP7_75t_R FILLER_86_996 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1049 ();
 FILLER_ASAP7_75t_R FILLER_86_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1224 ();
 FILLER_ASAP7_75t_R FILLER_86_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1236 ();
 FILLER_ASAP7_75t_R FILLER_86_1243 ();
 FILLER_ASAP7_75t_R FILLER_86_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1265 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_87_512 ();
 DECAPx1_ASAP7_75t_R FILLER_87_534 ();
 DECAPx6_ASAP7_75t_R FILLER_87_559 ();
 FILLER_ASAP7_75t_R FILLER_87_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_575 ();
 DECAPx10_ASAP7_75t_R FILLER_87_586 ();
 DECAPx10_ASAP7_75t_R FILLER_87_608 ();
 FILLER_ASAP7_75t_R FILLER_87_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_632 ();
 DECAPx4_ASAP7_75t_R FILLER_87_643 ();
 FILLER_ASAP7_75t_R FILLER_87_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_655 ();
 DECAPx10_ASAP7_75t_R FILLER_87_666 ();
 DECAPx10_ASAP7_75t_R FILLER_87_688 ();
 DECAPx2_ASAP7_75t_R FILLER_87_710 ();
 DECAPx10_ASAP7_75t_R FILLER_87_722 ();
 DECAPx10_ASAP7_75t_R FILLER_87_756 ();
 DECAPx10_ASAP7_75t_R FILLER_87_778 ();
 DECAPx4_ASAP7_75t_R FILLER_87_810 ();
 FILLER_ASAP7_75t_R FILLER_87_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_822 ();
 DECAPx10_ASAP7_75t_R FILLER_87_835 ();
 DECAPx10_ASAP7_75t_R FILLER_87_857 ();
 DECAPx10_ASAP7_75t_R FILLER_87_879 ();
 DECAPx10_ASAP7_75t_R FILLER_87_901 ();
 FILLER_ASAP7_75t_R FILLER_87_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_938 ();
 DECAPx2_ASAP7_75t_R FILLER_87_945 ();
 FILLER_ASAP7_75t_R FILLER_87_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_966 ();
 FILLER_ASAP7_75t_R FILLER_87_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_975 ();
 DECAPx4_ASAP7_75t_R FILLER_87_991 ();
 FILLER_ASAP7_75t_R FILLER_87_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1019 ();
 FILLER_ASAP7_75t_R FILLER_87_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1204 ();
 FILLER_ASAP7_75t_R FILLER_87_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1222 ();
 FILLER_ASAP7_75t_R FILLER_87_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_88_512 ();
 DECAPx1_ASAP7_75t_R FILLER_88_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_544 ();
 DECAPx1_ASAP7_75t_R FILLER_88_551 ();
 DECAPx4_ASAP7_75t_R FILLER_88_576 ();
 FILLER_ASAP7_75t_R FILLER_88_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_594 ();
 FILLER_ASAP7_75t_R FILLER_88_607 ();
 DECAPx2_ASAP7_75t_R FILLER_88_615 ();
 FILLER_ASAP7_75t_R FILLER_88_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_623 ();
 DECAPx2_ASAP7_75t_R FILLER_88_646 ();
 FILLER_ASAP7_75t_R FILLER_88_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_654 ();
 DECAPx10_ASAP7_75t_R FILLER_88_662 ();
 DECAPx10_ASAP7_75t_R FILLER_88_690 ();
 DECAPx10_ASAP7_75t_R FILLER_88_712 ();
 DECAPx6_ASAP7_75t_R FILLER_88_734 ();
 DECAPx1_ASAP7_75t_R FILLER_88_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_752 ();
 DECAPx1_ASAP7_75t_R FILLER_88_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_765 ();
 DECAPx4_ASAP7_75t_R FILLER_88_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_782 ();
 DECAPx10_ASAP7_75t_R FILLER_88_789 ();
 DECAPx10_ASAP7_75t_R FILLER_88_811 ();
 DECAPx10_ASAP7_75t_R FILLER_88_833 ();
 DECAPx4_ASAP7_75t_R FILLER_88_855 ();
 DECAPx10_ASAP7_75t_R FILLER_88_881 ();
 DECAPx1_ASAP7_75t_R FILLER_88_903 ();
 DECAPx10_ASAP7_75t_R FILLER_88_913 ();
 DECAPx2_ASAP7_75t_R FILLER_88_935 ();
 FILLER_ASAP7_75t_R FILLER_88_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_971 ();
 DECAPx10_ASAP7_75t_R FILLER_88_974 ();
 DECAPx4_ASAP7_75t_R FILLER_88_996 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1094 ();
 FILLER_ASAP7_75t_R FILLER_88_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1118 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1140 ();
 FILLER_ASAP7_75t_R FILLER_88_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1201 ();
 FILLER_ASAP7_75t_R FILLER_88_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1241 ();
 FILLER_ASAP7_75t_R FILLER_88_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1277 ();
 FILLER_ASAP7_75t_R FILLER_88_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_89_512 ();
 DECAPx6_ASAP7_75t_R FILLER_89_534 ();
 DECAPx1_ASAP7_75t_R FILLER_89_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_559 ();
 DECAPx4_ASAP7_75t_R FILLER_89_566 ();
 FILLER_ASAP7_75t_R FILLER_89_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_578 ();
 DECAPx6_ASAP7_75t_R FILLER_89_621 ();
 DECAPx2_ASAP7_75t_R FILLER_89_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_641 ();
 DECAPx10_ASAP7_75t_R FILLER_89_657 ();
 DECAPx2_ASAP7_75t_R FILLER_89_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_685 ();
 DECAPx4_ASAP7_75t_R FILLER_89_692 ();
 DECAPx6_ASAP7_75t_R FILLER_89_708 ();
 DECAPx1_ASAP7_75t_R FILLER_89_722 ();
 DECAPx10_ASAP7_75t_R FILLER_89_740 ();
 DECAPx10_ASAP7_75t_R FILLER_89_762 ();
 DECAPx10_ASAP7_75t_R FILLER_89_792 ();
 DECAPx2_ASAP7_75t_R FILLER_89_814 ();
 FILLER_ASAP7_75t_R FILLER_89_820 ();
 DECAPx6_ASAP7_75t_R FILLER_89_828 ();
 FILLER_ASAP7_75t_R FILLER_89_842 ();
 DECAPx10_ASAP7_75t_R FILLER_89_854 ();
 DECAPx10_ASAP7_75t_R FILLER_89_876 ();
 DECAPx10_ASAP7_75t_R FILLER_89_898 ();
 DECAPx10_ASAP7_75t_R FILLER_89_920 ();
 DECAPx10_ASAP7_75t_R FILLER_89_942 ();
 DECAPx10_ASAP7_75t_R FILLER_89_964 ();
 DECAPx10_ASAP7_75t_R FILLER_89_986 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1062 ();
 FILLER_ASAP7_75t_R FILLER_89_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1078 ();
 FILLER_ASAP7_75t_R FILLER_89_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_90_512 ();
 DECAPx10_ASAP7_75t_R FILLER_90_534 ();
 DECAPx4_ASAP7_75t_R FILLER_90_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_566 ();
 DECAPx2_ASAP7_75t_R FILLER_90_573 ();
 FILLER_ASAP7_75t_R FILLER_90_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_581 ();
 DECAPx10_ASAP7_75t_R FILLER_90_588 ();
 DECAPx10_ASAP7_75t_R FILLER_90_610 ();
 DECAPx10_ASAP7_75t_R FILLER_90_632 ();
 DECAPx6_ASAP7_75t_R FILLER_90_654 ();
 DECAPx1_ASAP7_75t_R FILLER_90_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_672 ();
 FILLER_ASAP7_75t_R FILLER_90_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_687 ();
 DECAPx4_ASAP7_75t_R FILLER_90_694 ();
 DECAPx10_ASAP7_75t_R FILLER_90_710 ();
 DECAPx2_ASAP7_75t_R FILLER_90_732 ();
 DECAPx10_ASAP7_75t_R FILLER_90_750 ();
 DECAPx1_ASAP7_75t_R FILLER_90_772 ();
 DECAPx10_ASAP7_75t_R FILLER_90_782 ();
 DECAPx6_ASAP7_75t_R FILLER_90_804 ();
 DECAPx1_ASAP7_75t_R FILLER_90_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_822 ();
 FILLER_ASAP7_75t_R FILLER_90_829 ();
 DECAPx10_ASAP7_75t_R FILLER_90_837 ();
 DECAPx10_ASAP7_75t_R FILLER_90_859 ();
 DECAPx2_ASAP7_75t_R FILLER_90_881 ();
 DECAPx10_ASAP7_75t_R FILLER_90_914 ();
 DECAPx10_ASAP7_75t_R FILLER_90_936 ();
 DECAPx6_ASAP7_75t_R FILLER_90_958 ();
 DECAPx6_ASAP7_75t_R FILLER_90_974 ();
 FILLER_ASAP7_75t_R FILLER_90_988 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1131 ();
 FILLER_ASAP7_75t_R FILLER_90_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1191 ();
 FILLER_ASAP7_75t_R FILLER_90_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1215 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_91_512 ();
 FILLER_ASAP7_75t_R FILLER_91_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_536 ();
 FILLER_ASAP7_75t_R FILLER_91_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_566 ();
 DECAPx10_ASAP7_75t_R FILLER_91_594 ();
 DECAPx10_ASAP7_75t_R FILLER_91_616 ();
 DECAPx2_ASAP7_75t_R FILLER_91_638 ();
 FILLER_ASAP7_75t_R FILLER_91_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_646 ();
 DECAPx2_ASAP7_75t_R FILLER_91_669 ();
 FILLER_ASAP7_75t_R FILLER_91_687 ();
 DECAPx10_ASAP7_75t_R FILLER_91_701 ();
 DECAPx2_ASAP7_75t_R FILLER_91_723 ();
 DECAPx6_ASAP7_75t_R FILLER_91_759 ();
 DECAPx1_ASAP7_75t_R FILLER_91_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_777 ();
 DECAPx10_ASAP7_75t_R FILLER_91_786 ();
 DECAPx6_ASAP7_75t_R FILLER_91_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_822 ();
 DECAPx4_ASAP7_75t_R FILLER_91_833 ();
 DECAPx4_ASAP7_75t_R FILLER_91_859 ();
 FILLER_ASAP7_75t_R FILLER_91_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_871 ();
 DECAPx1_ASAP7_75t_R FILLER_91_886 ();
 FILLER_ASAP7_75t_R FILLER_91_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_898 ();
 FILLER_ASAP7_75t_R FILLER_91_905 ();
 DECAPx2_ASAP7_75t_R FILLER_91_915 ();
 FILLER_ASAP7_75t_R FILLER_91_921 ();
 DECAPx2_ASAP7_75t_R FILLER_91_950 ();
 DECAPx10_ASAP7_75t_R FILLER_91_964 ();
 DECAPx10_ASAP7_75t_R FILLER_91_986 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1032 ();
 FILLER_ASAP7_75t_R FILLER_91_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1088 ();
 FILLER_ASAP7_75t_R FILLER_91_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1147 ();
 FILLER_ASAP7_75t_R FILLER_91_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1178 ();
 FILLER_ASAP7_75t_R FILLER_91_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1248 ();
 FILLER_ASAP7_75t_R FILLER_91_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_92_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_526 ();
 DECAPx2_ASAP7_75t_R FILLER_92_545 ();
 DECAPx4_ASAP7_75t_R FILLER_92_572 ();
 FILLER_ASAP7_75t_R FILLER_92_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_584 ();
 DECAPx10_ASAP7_75t_R FILLER_92_606 ();
 DECAPx4_ASAP7_75t_R FILLER_92_628 ();
 DECAPx10_ASAP7_75t_R FILLER_92_648 ();
 DECAPx4_ASAP7_75t_R FILLER_92_670 ();
 FILLER_ASAP7_75t_R FILLER_92_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_682 ();
 FILLER_ASAP7_75t_R FILLER_92_689 ();
 DECAPx6_ASAP7_75t_R FILLER_92_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_715 ();
 DECAPx2_ASAP7_75t_R FILLER_92_726 ();
 FILLER_ASAP7_75t_R FILLER_92_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_734 ();
 DECAPx6_ASAP7_75t_R FILLER_92_741 ();
 FILLER_ASAP7_75t_R FILLER_92_755 ();
 DECAPx10_ASAP7_75t_R FILLER_92_763 ();
 DECAPx4_ASAP7_75t_R FILLER_92_785 ();
 FILLER_ASAP7_75t_R FILLER_92_795 ();
 DECAPx10_ASAP7_75t_R FILLER_92_803 ();
 DECAPx10_ASAP7_75t_R FILLER_92_825 ();
 DECAPx10_ASAP7_75t_R FILLER_92_847 ();
 DECAPx10_ASAP7_75t_R FILLER_92_869 ();
 DECAPx10_ASAP7_75t_R FILLER_92_891 ();
 DECAPx4_ASAP7_75t_R FILLER_92_913 ();
 FILLER_ASAP7_75t_R FILLER_92_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_933 ();
 DECAPx4_ASAP7_75t_R FILLER_92_940 ();
 FILLER_ASAP7_75t_R FILLER_92_950 ();
 DECAPx6_ASAP7_75t_R FILLER_92_958 ();
 DECAPx10_ASAP7_75t_R FILLER_92_974 ();
 DECAPx4_ASAP7_75t_R FILLER_92_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1094 ();
 FILLER_ASAP7_75t_R FILLER_92_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1140 ();
 FILLER_ASAP7_75t_R FILLER_92_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_93_512 ();
 FILLER_ASAP7_75t_R FILLER_93_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_542 ();
 FILLER_ASAP7_75t_R FILLER_93_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_553 ();
 DECAPx10_ASAP7_75t_R FILLER_93_560 ();
 DECAPx1_ASAP7_75t_R FILLER_93_582 ();
 DECAPx10_ASAP7_75t_R FILLER_93_592 ();
 DECAPx6_ASAP7_75t_R FILLER_93_614 ();
 DECAPx1_ASAP7_75t_R FILLER_93_628 ();
 DECAPx10_ASAP7_75t_R FILLER_93_662 ();
 FILLER_ASAP7_75t_R FILLER_93_684 ();
 DECAPx10_ASAP7_75t_R FILLER_93_692 ();
 DECAPx10_ASAP7_75t_R FILLER_93_714 ();
 DECAPx6_ASAP7_75t_R FILLER_93_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_753 ();
 DECAPx10_ASAP7_75t_R FILLER_93_779 ();
 DECAPx10_ASAP7_75t_R FILLER_93_801 ();
 DECAPx10_ASAP7_75t_R FILLER_93_823 ();
 DECAPx6_ASAP7_75t_R FILLER_93_845 ();
 FILLER_ASAP7_75t_R FILLER_93_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_861 ();
 DECAPx10_ASAP7_75t_R FILLER_93_874 ();
 DECAPx10_ASAP7_75t_R FILLER_93_896 ();
 DECAPx1_ASAP7_75t_R FILLER_93_918 ();
 FILLER_ASAP7_75t_R FILLER_93_948 ();
 DECAPx1_ASAP7_75t_R FILLER_93_957 ();
 DECAPx10_ASAP7_75t_R FILLER_93_971 ();
 FILLER_ASAP7_75t_R FILLER_93_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_995 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_93_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1045 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1054 ();
 FILLER_ASAP7_75t_R FILLER_93_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1079 ();
 FILLER_ASAP7_75t_R FILLER_93_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_94_512 ();
 DECAPx1_ASAP7_75t_R FILLER_94_534 ();
 DECAPx4_ASAP7_75t_R FILLER_94_565 ();
 DECAPx10_ASAP7_75t_R FILLER_94_587 ();
 DECAPx10_ASAP7_75t_R FILLER_94_609 ();
 DECAPx10_ASAP7_75t_R FILLER_94_631 ();
 DECAPx2_ASAP7_75t_R FILLER_94_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_659 ();
 FILLER_ASAP7_75t_R FILLER_94_683 ();
 DECAPx2_ASAP7_75t_R FILLER_94_696 ();
 FILLER_ASAP7_75t_R FILLER_94_702 ();
 DECAPx2_ASAP7_75t_R FILLER_94_713 ();
 FILLER_ASAP7_75t_R FILLER_94_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_721 ();
 DECAPx1_ASAP7_75t_R FILLER_94_729 ();
 DECAPx10_ASAP7_75t_R FILLER_94_784 ();
 DECAPx10_ASAP7_75t_R FILLER_94_806 ();
 DECAPx1_ASAP7_75t_R FILLER_94_828 ();
 DECAPx2_ASAP7_75t_R FILLER_94_850 ();
 FILLER_ASAP7_75t_R FILLER_94_856 ();
 DECAPx10_ASAP7_75t_R FILLER_94_864 ();
 DECAPx10_ASAP7_75t_R FILLER_94_886 ();
 DECAPx10_ASAP7_75t_R FILLER_94_908 ();
 DECAPx10_ASAP7_75t_R FILLER_94_930 ();
 DECAPx6_ASAP7_75t_R FILLER_94_952 ();
 DECAPx2_ASAP7_75t_R FILLER_94_966 ();
 DECAPx6_ASAP7_75t_R FILLER_94_974 ();
 FILLER_ASAP7_75t_R FILLER_94_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_990 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1043 ();
 FILLER_ASAP7_75t_R FILLER_94_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1091 ();
 FILLER_ASAP7_75t_R FILLER_94_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1120 ();
 FILLER_ASAP7_75t_R FILLER_94_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1128 ();
 FILLER_ASAP7_75t_R FILLER_94_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1146 ();
 FILLER_ASAP7_75t_R FILLER_94_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1218 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1240 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_95_512 ();
 DECAPx1_ASAP7_75t_R FILLER_95_534 ();
 DECAPx1_ASAP7_75t_R FILLER_95_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_552 ();
 DECAPx4_ASAP7_75t_R FILLER_95_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_571 ();
 DECAPx10_ASAP7_75t_R FILLER_95_593 ();
 DECAPx6_ASAP7_75t_R FILLER_95_615 ();
 FILLER_ASAP7_75t_R FILLER_95_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_631 ();
 DECAPx2_ASAP7_75t_R FILLER_95_638 ();
 FILLER_ASAP7_75t_R FILLER_95_644 ();
 FILLER_ASAP7_75t_R FILLER_95_668 ();
 DECAPx6_ASAP7_75t_R FILLER_95_684 ();
 DECAPx1_ASAP7_75t_R FILLER_95_698 ();
 DECAPx1_ASAP7_75t_R FILLER_95_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_716 ();
 DECAPx2_ASAP7_75t_R FILLER_95_744 ();
 FILLER_ASAP7_75t_R FILLER_95_750 ();
 DECAPx2_ASAP7_75t_R FILLER_95_768 ();
 FILLER_ASAP7_75t_R FILLER_95_774 ();
 DECAPx2_ASAP7_75t_R FILLER_95_788 ();
 FILLER_ASAP7_75t_R FILLER_95_794 ();
 DECAPx2_ASAP7_75t_R FILLER_95_816 ();
 FILLER_ASAP7_75t_R FILLER_95_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_824 ();
 DECAPx10_ASAP7_75t_R FILLER_95_839 ();
 DECAPx10_ASAP7_75t_R FILLER_95_861 ();
 DECAPx10_ASAP7_75t_R FILLER_95_883 ();
 DECAPx4_ASAP7_75t_R FILLER_95_905 ();
 FILLER_ASAP7_75t_R FILLER_95_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_917 ();
 DECAPx10_ASAP7_75t_R FILLER_95_932 ();
 DECAPx10_ASAP7_75t_R FILLER_95_954 ();
 DECAPx4_ASAP7_75t_R FILLER_95_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_986 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1001 ();
 FILLER_ASAP7_75t_R FILLER_95_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_95_1113 ();
 FILLER_ASAP7_75t_R FILLER_95_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1125 ();
 DECAPx4_ASAP7_75t_R FILLER_95_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1221 ();
 FILLER_ASAP7_75t_R FILLER_95_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_96_512 ();
 DECAPx2_ASAP7_75t_R FILLER_96_534 ();
 DECAPx10_ASAP7_75t_R FILLER_96_550 ();
 DECAPx4_ASAP7_75t_R FILLER_96_572 ();
 DECAPx10_ASAP7_75t_R FILLER_96_590 ();
 DECAPx2_ASAP7_75t_R FILLER_96_612 ();
 DECAPx1_ASAP7_75t_R FILLER_96_650 ();
 DECAPx6_ASAP7_75t_R FILLER_96_660 ();
 FILLER_ASAP7_75t_R FILLER_96_674 ();
 DECAPx2_ASAP7_75t_R FILLER_96_683 ();
 DECAPx4_ASAP7_75t_R FILLER_96_703 ();
 FILLER_ASAP7_75t_R FILLER_96_713 ();
 DECAPx10_ASAP7_75t_R FILLER_96_724 ();
 DECAPx10_ASAP7_75t_R FILLER_96_746 ();
 DECAPx4_ASAP7_75t_R FILLER_96_768 ();
 FILLER_ASAP7_75t_R FILLER_96_778 ();
 DECAPx10_ASAP7_75t_R FILLER_96_786 ();
 DECAPx1_ASAP7_75t_R FILLER_96_818 ();
 DECAPx10_ASAP7_75t_R FILLER_96_860 ();
 FILLER_ASAP7_75t_R FILLER_96_882 ();
 DECAPx1_ASAP7_75t_R FILLER_96_893 ();
 DECAPx6_ASAP7_75t_R FILLER_96_917 ();
 FILLER_ASAP7_75t_R FILLER_96_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_952 ();
 DECAPx1_ASAP7_75t_R FILLER_96_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_971 ();
 DECAPx6_ASAP7_75t_R FILLER_96_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_988 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1075 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1097 ();
 FILLER_ASAP7_75t_R FILLER_96_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_96_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_96_1256 ();
 FILLER_ASAP7_75t_R FILLER_96_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1268 ();
 DECAPx2_ASAP7_75t_R FILLER_97_512 ();
 FILLER_ASAP7_75t_R FILLER_97_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_520 ();
 DECAPx6_ASAP7_75t_R FILLER_97_527 ();
 FILLER_ASAP7_75t_R FILLER_97_541 ();
 DECAPx2_ASAP7_75t_R FILLER_97_551 ();
 FILLER_ASAP7_75t_R FILLER_97_557 ();
 DECAPx6_ASAP7_75t_R FILLER_97_565 ();
 DECAPx10_ASAP7_75t_R FILLER_97_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_628 ();
 DECAPx2_ASAP7_75t_R FILLER_97_647 ();
 DECAPx2_ASAP7_75t_R FILLER_97_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_670 ();
 DECAPx6_ASAP7_75t_R FILLER_97_689 ();
 FILLER_ASAP7_75t_R FILLER_97_703 ();
 DECAPx6_ASAP7_75t_R FILLER_97_713 ();
 FILLER_ASAP7_75t_R FILLER_97_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_729 ();
 DECAPx4_ASAP7_75t_R FILLER_97_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_746 ();
 DECAPx10_ASAP7_75t_R FILLER_97_759 ();
 DECAPx6_ASAP7_75t_R FILLER_97_781 ();
 FILLER_ASAP7_75t_R FILLER_97_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_797 ();
 DECAPx6_ASAP7_75t_R FILLER_97_816 ();
 DECAPx1_ASAP7_75t_R FILLER_97_830 ();
 DECAPx6_ASAP7_75t_R FILLER_97_844 ();
 DECAPx1_ASAP7_75t_R FILLER_97_858 ();
 DECAPx2_ASAP7_75t_R FILLER_97_868 ();
 DECAPx10_ASAP7_75t_R FILLER_97_893 ();
 DECAPx10_ASAP7_75t_R FILLER_97_915 ();
 FILLER_ASAP7_75t_R FILLER_97_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_939 ();
 DECAPx10_ASAP7_75t_R FILLER_97_978 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1112 ();
 FILLER_ASAP7_75t_R FILLER_97_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1134 ();
 FILLER_ASAP7_75t_R FILLER_97_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1176 ();
 FILLER_ASAP7_75t_R FILLER_97_1186 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1208 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1233 ();
 FILLER_ASAP7_75t_R FILLER_97_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_98_512 ();
 FILLER_ASAP7_75t_R FILLER_98_553 ();
 DECAPx6_ASAP7_75t_R FILLER_98_561 ();
 DECAPx6_ASAP7_75t_R FILLER_98_605 ();
 FILLER_ASAP7_75t_R FILLER_98_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_621 ();
 DECAPx6_ASAP7_75t_R FILLER_98_642 ();
 FILLER_ASAP7_75t_R FILLER_98_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_658 ();
 FILLER_ASAP7_75t_R FILLER_98_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_670 ();
 DECAPx10_ASAP7_75t_R FILLER_98_681 ();
 FILLER_ASAP7_75t_R FILLER_98_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_705 ();
 DECAPx2_ASAP7_75t_R FILLER_98_720 ();
 DECAPx6_ASAP7_75t_R FILLER_98_729 ();
 FILLER_ASAP7_75t_R FILLER_98_743 ();
 DECAPx4_ASAP7_75t_R FILLER_98_764 ();
 FILLER_ASAP7_75t_R FILLER_98_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_776 ();
 FILLER_ASAP7_75t_R FILLER_98_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_785 ();
 DECAPx10_ASAP7_75t_R FILLER_98_792 ();
 DECAPx10_ASAP7_75t_R FILLER_98_814 ();
 DECAPx10_ASAP7_75t_R FILLER_98_836 ();
 DECAPx10_ASAP7_75t_R FILLER_98_858 ();
 DECAPx10_ASAP7_75t_R FILLER_98_880 ();
 DECAPx6_ASAP7_75t_R FILLER_98_902 ();
 FILLER_ASAP7_75t_R FILLER_98_916 ();
 DECAPx4_ASAP7_75t_R FILLER_98_932 ();
 DECAPx10_ASAP7_75t_R FILLER_98_950 ();
 DECAPx10_ASAP7_75t_R FILLER_98_974 ();
 DECAPx4_ASAP7_75t_R FILLER_98_996 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1083 ();
 FILLER_ASAP7_75t_R FILLER_98_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1170 ();
 FILLER_ASAP7_75t_R FILLER_98_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1227 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1284 ();
 FILLER_ASAP7_75t_R FILLER_98_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_99_512 ();
 DECAPx6_ASAP7_75t_R FILLER_99_534 ();
 DECAPx2_ASAP7_75t_R FILLER_99_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_554 ();
 DECAPx2_ASAP7_75t_R FILLER_99_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_582 ();
 DECAPx6_ASAP7_75t_R FILLER_99_613 ();
 DECAPx10_ASAP7_75t_R FILLER_99_641 ();
 DECAPx10_ASAP7_75t_R FILLER_99_663 ();
 DECAPx10_ASAP7_75t_R FILLER_99_685 ();
 DECAPx1_ASAP7_75t_R FILLER_99_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_711 ();
 DECAPx10_ASAP7_75t_R FILLER_99_745 ();
 DECAPx2_ASAP7_75t_R FILLER_99_767 ();
 FILLER_ASAP7_75t_R FILLER_99_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_775 ();
 DECAPx1_ASAP7_75t_R FILLER_99_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_786 ();
 DECAPx1_ASAP7_75t_R FILLER_99_793 ();
 DECAPx6_ASAP7_75t_R FILLER_99_807 ();
 DECAPx2_ASAP7_75t_R FILLER_99_821 ();
 DECAPx6_ASAP7_75t_R FILLER_99_849 ();
 FILLER_ASAP7_75t_R FILLER_99_863 ();
 DECAPx10_ASAP7_75t_R FILLER_99_883 ();
 DECAPx1_ASAP7_75t_R FILLER_99_925 ();
 DECAPx4_ASAP7_75t_R FILLER_99_945 ();
 DECAPx10_ASAP7_75t_R FILLER_99_973 ();
 FILLER_ASAP7_75t_R FILLER_99_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_997 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1012 ();
 FILLER_ASAP7_75t_R FILLER_99_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1203 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_100_512 ();
 FILLER_ASAP7_75t_R FILLER_100_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_545 ();
 DECAPx6_ASAP7_75t_R FILLER_100_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_586 ();
 DECAPx4_ASAP7_75t_R FILLER_100_596 ();
 FILLER_ASAP7_75t_R FILLER_100_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_623 ();
 DECAPx6_ASAP7_75t_R FILLER_100_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_648 ();
 DECAPx1_ASAP7_75t_R FILLER_100_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_660 ();
 DECAPx10_ASAP7_75t_R FILLER_100_667 ();
 DECAPx1_ASAP7_75t_R FILLER_100_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_693 ();
 DECAPx10_ASAP7_75t_R FILLER_100_714 ();
 DECAPx10_ASAP7_75t_R FILLER_100_736 ();
 DECAPx6_ASAP7_75t_R FILLER_100_758 ();
 DECAPx2_ASAP7_75t_R FILLER_100_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_778 ();
 DECAPx6_ASAP7_75t_R FILLER_100_797 ();
 DECAPx1_ASAP7_75t_R FILLER_100_811 ();
 DECAPx10_ASAP7_75t_R FILLER_100_831 ();
 DECAPx10_ASAP7_75t_R FILLER_100_853 ();
 DECAPx10_ASAP7_75t_R FILLER_100_875 ();
 DECAPx10_ASAP7_75t_R FILLER_100_897 ();
 DECAPx10_ASAP7_75t_R FILLER_100_919 ();
 DECAPx1_ASAP7_75t_R FILLER_100_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_945 ();
 DECAPx6_ASAP7_75t_R FILLER_100_974 ();
 DECAPx1_ASAP7_75t_R FILLER_100_988 ();
 DECAPx6_ASAP7_75t_R FILLER_100_998 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1157 ();
 FILLER_ASAP7_75t_R FILLER_100_1167 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1224 ();
 FILLER_ASAP7_75t_R FILLER_100_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_101_512 ();
 FILLER_ASAP7_75t_R FILLER_101_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_536 ();
 DECAPx10_ASAP7_75t_R FILLER_101_546 ();
 FILLER_ASAP7_75t_R FILLER_101_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_570 ();
 DECAPx1_ASAP7_75t_R FILLER_101_589 ();
 DECAPx10_ASAP7_75t_R FILLER_101_599 ();
 DECAPx6_ASAP7_75t_R FILLER_101_621 ();
 FILLER_ASAP7_75t_R FILLER_101_635 ();
 DECAPx10_ASAP7_75t_R FILLER_101_644 ();
 DECAPx10_ASAP7_75t_R FILLER_101_666 ();
 DECAPx1_ASAP7_75t_R FILLER_101_688 ();
 DECAPx4_ASAP7_75t_R FILLER_101_704 ();
 FILLER_ASAP7_75t_R FILLER_101_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_720 ();
 DECAPx10_ASAP7_75t_R FILLER_101_751 ();
 DECAPx10_ASAP7_75t_R FILLER_101_773 ();
 DECAPx10_ASAP7_75t_R FILLER_101_795 ();
 DECAPx10_ASAP7_75t_R FILLER_101_817 ();
 DECAPx6_ASAP7_75t_R FILLER_101_839 ();
 DECAPx2_ASAP7_75t_R FILLER_101_853 ();
 DECAPx10_ASAP7_75t_R FILLER_101_893 ();
 DECAPx6_ASAP7_75t_R FILLER_101_915 ();
 DECAPx1_ASAP7_75t_R FILLER_101_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_933 ();
 DECAPx6_ASAP7_75t_R FILLER_101_948 ();
 DECAPx2_ASAP7_75t_R FILLER_101_962 ();
 DECAPx6_ASAP7_75t_R FILLER_101_975 ();
 FILLER_ASAP7_75t_R FILLER_101_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1025 ();
 FILLER_ASAP7_75t_R FILLER_101_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1046 ();
 FILLER_ASAP7_75t_R FILLER_101_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1145 ();
 FILLER_ASAP7_75t_R FILLER_101_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1160 ();
 FILLER_ASAP7_75t_R FILLER_101_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1215 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1237 ();
 FILLER_ASAP7_75t_R FILLER_101_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_102_512 ();
 DECAPx2_ASAP7_75t_R FILLER_102_534 ();
 DECAPx10_ASAP7_75t_R FILLER_102_550 ();
 DECAPx2_ASAP7_75t_R FILLER_102_572 ();
 DECAPx10_ASAP7_75t_R FILLER_102_599 ();
 DECAPx10_ASAP7_75t_R FILLER_102_621 ();
 FILLER_ASAP7_75t_R FILLER_102_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_645 ();
 DECAPx10_ASAP7_75t_R FILLER_102_653 ();
 DECAPx10_ASAP7_75t_R FILLER_102_675 ();
 DECAPx1_ASAP7_75t_R FILLER_102_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_701 ();
 DECAPx10_ASAP7_75t_R FILLER_102_714 ();
 DECAPx2_ASAP7_75t_R FILLER_102_736 ();
 FILLER_ASAP7_75t_R FILLER_102_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_744 ();
 DECAPx10_ASAP7_75t_R FILLER_102_754 ();
 FILLER_ASAP7_75t_R FILLER_102_776 ();
 DECAPx6_ASAP7_75t_R FILLER_102_784 ();
 DECAPx2_ASAP7_75t_R FILLER_102_798 ();
 DECAPx10_ASAP7_75t_R FILLER_102_818 ();
 DECAPx1_ASAP7_75t_R FILLER_102_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_844 ();
 DECAPx10_ASAP7_75t_R FILLER_102_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_881 ();
 DECAPx6_ASAP7_75t_R FILLER_102_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_910 ();
 FILLER_ASAP7_75t_R FILLER_102_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_945 ();
 DECAPx6_ASAP7_75t_R FILLER_102_953 ();
 DECAPx1_ASAP7_75t_R FILLER_102_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_971 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1031 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1070 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1150 ();
 FILLER_ASAP7_75t_R FILLER_102_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1194 ();
 FILLER_ASAP7_75t_R FILLER_102_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_103_512 ();
 DECAPx6_ASAP7_75t_R FILLER_103_534 ();
 FILLER_ASAP7_75t_R FILLER_103_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_550 ();
 DECAPx10_ASAP7_75t_R FILLER_103_565 ();
 DECAPx10_ASAP7_75t_R FILLER_103_587 ();
 DECAPx10_ASAP7_75t_R FILLER_103_609 ();
 DECAPx10_ASAP7_75t_R FILLER_103_631 ();
 DECAPx6_ASAP7_75t_R FILLER_103_653 ();
 DECAPx1_ASAP7_75t_R FILLER_103_667 ();
 DECAPx10_ASAP7_75t_R FILLER_103_681 ();
 DECAPx4_ASAP7_75t_R FILLER_103_703 ();
 FILLER_ASAP7_75t_R FILLER_103_713 ();
 DECAPx10_ASAP7_75t_R FILLER_103_729 ();
 DECAPx10_ASAP7_75t_R FILLER_103_751 ();
 DECAPx2_ASAP7_75t_R FILLER_103_773 ();
 DECAPx6_ASAP7_75t_R FILLER_103_795 ();
 DECAPx10_ASAP7_75t_R FILLER_103_821 ();
 DECAPx6_ASAP7_75t_R FILLER_103_843 ();
 DECAPx10_ASAP7_75t_R FILLER_103_867 ();
 DECAPx2_ASAP7_75t_R FILLER_103_889 ();
 DECAPx10_ASAP7_75t_R FILLER_103_927 ();
 FILLER_ASAP7_75t_R FILLER_103_949 ();
 DECAPx10_ASAP7_75t_R FILLER_103_961 ();
 DECAPx4_ASAP7_75t_R FILLER_103_983 ();
 DECAPx4_ASAP7_75t_R FILLER_103_999 ();
 FILLER_ASAP7_75t_R FILLER_103_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1040 ();
 FILLER_ASAP7_75t_R FILLER_103_1062 ();
 FILLER_ASAP7_75t_R FILLER_103_1086 ();
 FILLER_ASAP7_75t_R FILLER_103_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1172 ();
 FILLER_ASAP7_75t_R FILLER_103_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1281 ();
 FILLER_ASAP7_75t_R FILLER_103_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_104_512 ();
 FILLER_ASAP7_75t_R FILLER_104_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_573 ();
 DECAPx10_ASAP7_75t_R FILLER_104_580 ();
 DECAPx10_ASAP7_75t_R FILLER_104_602 ();
 DECAPx10_ASAP7_75t_R FILLER_104_624 ();
 DECAPx10_ASAP7_75t_R FILLER_104_646 ();
 DECAPx10_ASAP7_75t_R FILLER_104_668 ();
 DECAPx10_ASAP7_75t_R FILLER_104_690 ();
 DECAPx10_ASAP7_75t_R FILLER_104_712 ();
 DECAPx6_ASAP7_75t_R FILLER_104_734 ();
 FILLER_ASAP7_75t_R FILLER_104_748 ();
 DECAPx10_ASAP7_75t_R FILLER_104_764 ();
 DECAPx10_ASAP7_75t_R FILLER_104_786 ();
 DECAPx4_ASAP7_75t_R FILLER_104_808 ();
 DECAPx10_ASAP7_75t_R FILLER_104_834 ();
 DECAPx2_ASAP7_75t_R FILLER_104_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_862 ();
 DECAPx10_ASAP7_75t_R FILLER_104_877 ();
 DECAPx4_ASAP7_75t_R FILLER_104_899 ();
 DECAPx10_ASAP7_75t_R FILLER_104_947 ();
 FILLER_ASAP7_75t_R FILLER_104_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_971 ();
 DECAPx10_ASAP7_75t_R FILLER_104_974 ();
 DECAPx10_ASAP7_75t_R FILLER_104_996 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1102 ();
 FILLER_ASAP7_75t_R FILLER_104_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1142 ();
 FILLER_ASAP7_75t_R FILLER_104_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_105_512 ();
 DECAPx6_ASAP7_75t_R FILLER_105_542 ();
 DECAPx2_ASAP7_75t_R FILLER_105_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_562 ();
 FILLER_ASAP7_75t_R FILLER_105_584 ();
 DECAPx10_ASAP7_75t_R FILLER_105_594 ();
 DECAPx6_ASAP7_75t_R FILLER_105_616 ();
 DECAPx1_ASAP7_75t_R FILLER_105_630 ();
 DECAPx2_ASAP7_75t_R FILLER_105_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_646 ();
 DECAPx1_ASAP7_75t_R FILLER_105_653 ();
 DECAPx10_ASAP7_75t_R FILLER_105_668 ();
 FILLER_ASAP7_75t_R FILLER_105_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_692 ();
 DECAPx1_ASAP7_75t_R FILLER_105_705 ();
 DECAPx10_ASAP7_75t_R FILLER_105_728 ();
 DECAPx10_ASAP7_75t_R FILLER_105_750 ();
 DECAPx10_ASAP7_75t_R FILLER_105_772 ();
 DECAPx4_ASAP7_75t_R FILLER_105_794 ();
 DECAPx6_ASAP7_75t_R FILLER_105_814 ();
 DECAPx6_ASAP7_75t_R FILLER_105_836 ();
 FILLER_ASAP7_75t_R FILLER_105_850 ();
 DECAPx4_ASAP7_75t_R FILLER_105_862 ();
 FILLER_ASAP7_75t_R FILLER_105_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_874 ();
 DECAPx2_ASAP7_75t_R FILLER_105_889 ();
 FILLER_ASAP7_75t_R FILLER_105_895 ();
 DECAPx4_ASAP7_75t_R FILLER_105_911 ();
 DECAPx10_ASAP7_75t_R FILLER_105_933 ();
 DECAPx2_ASAP7_75t_R FILLER_105_965 ();
 DECAPx10_ASAP7_75t_R FILLER_105_977 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_105_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1211 ();
 FILLER_ASAP7_75t_R FILLER_105_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1219 ();
 FILLER_ASAP7_75t_R FILLER_105_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1238 ();
 DECAPx6_ASAP7_75t_R FILLER_105_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_106_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_526 ();
 DECAPx4_ASAP7_75t_R FILLER_106_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_547 ();
 DECAPx4_ASAP7_75t_R FILLER_106_562 ();
 DECAPx10_ASAP7_75t_R FILLER_106_609 ();
 DECAPx10_ASAP7_75t_R FILLER_106_631 ();
 DECAPx6_ASAP7_75t_R FILLER_106_653 ();
 FILLER_ASAP7_75t_R FILLER_106_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_669 ();
 DECAPx4_ASAP7_75t_R FILLER_106_682 ();
 FILLER_ASAP7_75t_R FILLER_106_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_701 ();
 DECAPx4_ASAP7_75t_R FILLER_106_708 ();
 DECAPx6_ASAP7_75t_R FILLER_106_727 ();
 FILLER_ASAP7_75t_R FILLER_106_741 ();
 DECAPx10_ASAP7_75t_R FILLER_106_762 ();
 DECAPx10_ASAP7_75t_R FILLER_106_784 ();
 DECAPx10_ASAP7_75t_R FILLER_106_806 ();
 DECAPx10_ASAP7_75t_R FILLER_106_828 ();
 DECAPx10_ASAP7_75t_R FILLER_106_850 ();
 DECAPx10_ASAP7_75t_R FILLER_106_872 ();
 DECAPx4_ASAP7_75t_R FILLER_106_894 ();
 FILLER_ASAP7_75t_R FILLER_106_904 ();
 DECAPx6_ASAP7_75t_R FILLER_106_920 ();
 DECAPx1_ASAP7_75t_R FILLER_106_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_938 ();
 FILLER_ASAP7_75t_R FILLER_106_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_971 ();
 DECAPx6_ASAP7_75t_R FILLER_106_974 ();
 FILLER_ASAP7_75t_R FILLER_106_988 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1070 ();
 FILLER_ASAP7_75t_R FILLER_106_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1091 ();
 FILLER_ASAP7_75t_R FILLER_106_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1117 ();
 FILLER_ASAP7_75t_R FILLER_106_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1257 ();
 FILLER_ASAP7_75t_R FILLER_106_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_107_512 ();
 DECAPx2_ASAP7_75t_R FILLER_107_534 ();
 FILLER_ASAP7_75t_R FILLER_107_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_542 ();
 DECAPx10_ASAP7_75t_R FILLER_107_547 ();
 FILLER_ASAP7_75t_R FILLER_107_569 ();
 DECAPx10_ASAP7_75t_R FILLER_107_581 ();
 DECAPx10_ASAP7_75t_R FILLER_107_603 ();
 DECAPx10_ASAP7_75t_R FILLER_107_625 ();
 DECAPx10_ASAP7_75t_R FILLER_107_647 ();
 DECAPx10_ASAP7_75t_R FILLER_107_669 ();
 DECAPx2_ASAP7_75t_R FILLER_107_691 ();
 FILLER_ASAP7_75t_R FILLER_107_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_699 ();
 DECAPx2_ASAP7_75t_R FILLER_107_712 ();
 DECAPx10_ASAP7_75t_R FILLER_107_727 ();
 DECAPx1_ASAP7_75t_R FILLER_107_749 ();
 DECAPx2_ASAP7_75t_R FILLER_107_759 ();
 DECAPx10_ASAP7_75t_R FILLER_107_771 ();
 DECAPx6_ASAP7_75t_R FILLER_107_793 ();
 DECAPx1_ASAP7_75t_R FILLER_107_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_811 ();
 DECAPx10_ASAP7_75t_R FILLER_107_820 ();
 DECAPx10_ASAP7_75t_R FILLER_107_842 ();
 DECAPx4_ASAP7_75t_R FILLER_107_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_874 ();
 DECAPx1_ASAP7_75t_R FILLER_107_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_897 ();
 DECAPx10_ASAP7_75t_R FILLER_107_926 ();
 DECAPx10_ASAP7_75t_R FILLER_107_948 ();
 DECAPx2_ASAP7_75t_R FILLER_107_970 ();
 FILLER_ASAP7_75t_R FILLER_107_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_978 ();
 DECAPx4_ASAP7_75t_R FILLER_107_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_999 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1028 ();
 FILLER_ASAP7_75t_R FILLER_107_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1071 ();
 FILLER_ASAP7_75t_R FILLER_107_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1123 ();
 DECAPx4_ASAP7_75t_R FILLER_107_1145 ();
 FILLER_ASAP7_75t_R FILLER_107_1155 ();
 FILLER_ASAP7_75t_R FILLER_107_1178 ();
 FILLER_ASAP7_75t_R FILLER_107_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1207 ();
 FILLER_ASAP7_75t_R FILLER_107_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_107_1280 ();
 FILLER_ASAP7_75t_R FILLER_107_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_108_512 ();
 DECAPx6_ASAP7_75t_R FILLER_108_534 ();
 FILLER_ASAP7_75t_R FILLER_108_548 ();
 DECAPx10_ASAP7_75t_R FILLER_108_583 ();
 DECAPx10_ASAP7_75t_R FILLER_108_605 ();
 DECAPx10_ASAP7_75t_R FILLER_108_627 ();
 DECAPx10_ASAP7_75t_R FILLER_108_649 ();
 DECAPx10_ASAP7_75t_R FILLER_108_671 ();
 DECAPx2_ASAP7_75t_R FILLER_108_693 ();
 FILLER_ASAP7_75t_R FILLER_108_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_701 ();
 DECAPx2_ASAP7_75t_R FILLER_108_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_716 ();
 DECAPx1_ASAP7_75t_R FILLER_108_726 ();
 DECAPx10_ASAP7_75t_R FILLER_108_733 ();
 DECAPx10_ASAP7_75t_R FILLER_108_755 ();
 DECAPx2_ASAP7_75t_R FILLER_108_777 ();
 FILLER_ASAP7_75t_R FILLER_108_783 ();
 DECAPx2_ASAP7_75t_R FILLER_108_805 ();
 FILLER_ASAP7_75t_R FILLER_108_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_813 ();
 DECAPx4_ASAP7_75t_R FILLER_108_826 ();
 DECAPx10_ASAP7_75t_R FILLER_108_858 ();
 DECAPx6_ASAP7_75t_R FILLER_108_880 ();
 DECAPx2_ASAP7_75t_R FILLER_108_894 ();
 DECAPx6_ASAP7_75t_R FILLER_108_914 ();
 FILLER_ASAP7_75t_R FILLER_108_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_930 ();
 DECAPx1_ASAP7_75t_R FILLER_108_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_949 ();
 DECAPx4_ASAP7_75t_R FILLER_108_960 ();
 FILLER_ASAP7_75t_R FILLER_108_970 ();
 DECAPx2_ASAP7_75t_R FILLER_108_974 ();
 DECAPx6_ASAP7_75t_R FILLER_108_986 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1008 ();
 FILLER_ASAP7_75t_R FILLER_108_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1093 ();
 FILLER_ASAP7_75t_R FILLER_108_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_109_512 ();
 DECAPx4_ASAP7_75t_R FILLER_109_562 ();
 DECAPx10_ASAP7_75t_R FILLER_109_582 ();
 DECAPx10_ASAP7_75t_R FILLER_109_604 ();
 DECAPx2_ASAP7_75t_R FILLER_109_626 ();
 FILLER_ASAP7_75t_R FILLER_109_632 ();
 DECAPx10_ASAP7_75t_R FILLER_109_643 ();
 DECAPx10_ASAP7_75t_R FILLER_109_665 ();
 DECAPx4_ASAP7_75t_R FILLER_109_687 ();
 FILLER_ASAP7_75t_R FILLER_109_697 ();
 FILLER_ASAP7_75t_R FILLER_109_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_726 ();
 FILLER_ASAP7_75t_R FILLER_109_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_750 ();
 DECAPx10_ASAP7_75t_R FILLER_109_769 ();
 DECAPx10_ASAP7_75t_R FILLER_109_791 ();
 DECAPx6_ASAP7_75t_R FILLER_109_813 ();
 FILLER_ASAP7_75t_R FILLER_109_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_850 ();
 DECAPx1_ASAP7_75t_R FILLER_109_859 ();
 DECAPx10_ASAP7_75t_R FILLER_109_869 ();
 DECAPx10_ASAP7_75t_R FILLER_109_891 ();
 DECAPx6_ASAP7_75t_R FILLER_109_913 ();
 FILLER_ASAP7_75t_R FILLER_109_927 ();
 DECAPx1_ASAP7_75t_R FILLER_109_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_947 ();
 DECAPx1_ASAP7_75t_R FILLER_109_956 ();
 DECAPx4_ASAP7_75t_R FILLER_109_978 ();
 FILLER_ASAP7_75t_R FILLER_109_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1116 ();
 FILLER_ASAP7_75t_R FILLER_109_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1215 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_110_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_526 ();
 DECAPx6_ASAP7_75t_R FILLER_110_535 ();
 DECAPx10_ASAP7_75t_R FILLER_110_570 ();
 DECAPx2_ASAP7_75t_R FILLER_110_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_598 ();
 DECAPx10_ASAP7_75t_R FILLER_110_613 ();
 DECAPx6_ASAP7_75t_R FILLER_110_635 ();
 DECAPx2_ASAP7_75t_R FILLER_110_655 ();
 DECAPx10_ASAP7_75t_R FILLER_110_675 ();
 DECAPx10_ASAP7_75t_R FILLER_110_697 ();
 DECAPx10_ASAP7_75t_R FILLER_110_719 ();
 DECAPx10_ASAP7_75t_R FILLER_110_741 ();
 DECAPx10_ASAP7_75t_R FILLER_110_763 ();
 FILLER_ASAP7_75t_R FILLER_110_785 ();
 DECAPx10_ASAP7_75t_R FILLER_110_801 ();
 DECAPx10_ASAP7_75t_R FILLER_110_823 ();
 DECAPx1_ASAP7_75t_R FILLER_110_845 ();
 DECAPx2_ASAP7_75t_R FILLER_110_855 ();
 DECAPx2_ASAP7_75t_R FILLER_110_877 ();
 DECAPx6_ASAP7_75t_R FILLER_110_893 ();
 DECAPx6_ASAP7_75t_R FILLER_110_921 ();
 DECAPx2_ASAP7_75t_R FILLER_110_935 ();
 DECAPx10_ASAP7_75t_R FILLER_110_974 ();
 DECAPx6_ASAP7_75t_R FILLER_110_996 ();
 FILLER_ASAP7_75t_R FILLER_110_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1092 ();
 FILLER_ASAP7_75t_R FILLER_110_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1197 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1285 ();
 FILLER_ASAP7_75t_R FILLER_110_1291 ();
 DECAPx4_ASAP7_75t_R FILLER_111_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_522 ();
 DECAPx6_ASAP7_75t_R FILLER_111_532 ();
 DECAPx1_ASAP7_75t_R FILLER_111_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_562 ();
 DECAPx10_ASAP7_75t_R FILLER_111_596 ();
 DECAPx10_ASAP7_75t_R FILLER_111_618 ();
 DECAPx10_ASAP7_75t_R FILLER_111_640 ();
 DECAPx6_ASAP7_75t_R FILLER_111_662 ();
 DECAPx10_ASAP7_75t_R FILLER_111_688 ();
 FILLER_ASAP7_75t_R FILLER_111_710 ();
 DECAPx10_ASAP7_75t_R FILLER_111_728 ();
 DECAPx4_ASAP7_75t_R FILLER_111_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_760 ();
 DECAPx10_ASAP7_75t_R FILLER_111_771 ();
 DECAPx1_ASAP7_75t_R FILLER_111_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_797 ();
 DECAPx10_ASAP7_75t_R FILLER_111_804 ();
 DECAPx6_ASAP7_75t_R FILLER_111_826 ();
 DECAPx10_ASAP7_75t_R FILLER_111_850 ();
 DECAPx10_ASAP7_75t_R FILLER_111_872 ();
 DECAPx2_ASAP7_75t_R FILLER_111_894 ();
 DECAPx10_ASAP7_75t_R FILLER_111_944 ();
 DECAPx1_ASAP7_75t_R FILLER_111_966 ();
 DECAPx1_ASAP7_75t_R FILLER_111_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_980 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_111_1200 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_112_512 ();
 FILLER_ASAP7_75t_R FILLER_112_518 ();
 DECAPx6_ASAP7_75t_R FILLER_112_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_556 ();
 FILLER_ASAP7_75t_R FILLER_112_565 ();
 DECAPx10_ASAP7_75t_R FILLER_112_581 ();
 DECAPx10_ASAP7_75t_R FILLER_112_603 ();
 DECAPx10_ASAP7_75t_R FILLER_112_625 ();
 DECAPx2_ASAP7_75t_R FILLER_112_647 ();
 FILLER_ASAP7_75t_R FILLER_112_653 ();
 DECAPx6_ASAP7_75t_R FILLER_112_673 ();
 DECAPx1_ASAP7_75t_R FILLER_112_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_691 ();
 DECAPx10_ASAP7_75t_R FILLER_112_700 ();
 DECAPx10_ASAP7_75t_R FILLER_112_722 ();
 DECAPx10_ASAP7_75t_R FILLER_112_744 ();
 FILLER_ASAP7_75t_R FILLER_112_766 ();
 DECAPx6_ASAP7_75t_R FILLER_112_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_800 ();
 DECAPx2_ASAP7_75t_R FILLER_112_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_815 ();
 DECAPx1_ASAP7_75t_R FILLER_112_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_834 ();
 DECAPx10_ASAP7_75t_R FILLER_112_845 ();
 DECAPx2_ASAP7_75t_R FILLER_112_867 ();
 FILLER_ASAP7_75t_R FILLER_112_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_875 ();
 DECAPx4_ASAP7_75t_R FILLER_112_920 ();
 FILLER_ASAP7_75t_R FILLER_112_930 ();
 DECAPx10_ASAP7_75t_R FILLER_112_940 ();
 DECAPx4_ASAP7_75t_R FILLER_112_962 ();
 DECAPx2_ASAP7_75t_R FILLER_112_974 ();
 FILLER_ASAP7_75t_R FILLER_112_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_982 ();
 DECAPx6_ASAP7_75t_R FILLER_112_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1095 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1147 ();
 FILLER_ASAP7_75t_R FILLER_112_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1223 ();
 FILLER_ASAP7_75t_R FILLER_112_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1231 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1238 ();
 FILLER_ASAP7_75t_R FILLER_112_1252 ();
 DECAPx4_ASAP7_75t_R FILLER_112_1281 ();
 FILLER_ASAP7_75t_R FILLER_112_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_113_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_526 ();
 DECAPx10_ASAP7_75t_R FILLER_113_571 ();
 DECAPx4_ASAP7_75t_R FILLER_113_593 ();
 FILLER_ASAP7_75t_R FILLER_113_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_605 ();
 DECAPx10_ASAP7_75t_R FILLER_113_619 ();
 DECAPx2_ASAP7_75t_R FILLER_113_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_647 ();
 DECAPx6_ASAP7_75t_R FILLER_113_669 ();
 DECAPx1_ASAP7_75t_R FILLER_113_683 ();
 DECAPx10_ASAP7_75t_R FILLER_113_695 ();
 DECAPx2_ASAP7_75t_R FILLER_113_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_723 ();
 DECAPx1_ASAP7_75t_R FILLER_113_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_754 ();
 DECAPx4_ASAP7_75t_R FILLER_113_779 ();
 FILLER_ASAP7_75t_R FILLER_113_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_791 ();
 FILLER_ASAP7_75t_R FILLER_113_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_824 ();
 DECAPx1_ASAP7_75t_R FILLER_113_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_839 ();
 DECAPx2_ASAP7_75t_R FILLER_113_852 ();
 FILLER_ASAP7_75t_R FILLER_113_858 ();
 FILLER_ASAP7_75t_R FILLER_113_874 ();
 DECAPx2_ASAP7_75t_R FILLER_113_898 ();
 DECAPx4_ASAP7_75t_R FILLER_113_918 ();
 DECAPx10_ASAP7_75t_R FILLER_113_949 ();
 FILLER_ASAP7_75t_R FILLER_113_971 ();
 DECAPx6_ASAP7_75t_R FILLER_113_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_993 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1078 ();
 FILLER_ASAP7_75t_R FILLER_113_1088 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1096 ();
 FILLER_ASAP7_75t_R FILLER_113_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1141 ();
 FILLER_ASAP7_75t_R FILLER_113_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1160 ();
 FILLER_ASAP7_75t_R FILLER_113_1166 ();
 FILLER_ASAP7_75t_R FILLER_113_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1232 ();
 FILLER_ASAP7_75t_R FILLER_113_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1248 ();
 FILLER_ASAP7_75t_R FILLER_113_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_114_512 ();
 DECAPx1_ASAP7_75t_R FILLER_114_526 ();
 DECAPx1_ASAP7_75t_R FILLER_114_540 ();
 DECAPx2_ASAP7_75t_R FILLER_114_554 ();
 FILLER_ASAP7_75t_R FILLER_114_560 ();
 DECAPx10_ASAP7_75t_R FILLER_114_570 ();
 DECAPx6_ASAP7_75t_R FILLER_114_606 ();
 DECAPx1_ASAP7_75t_R FILLER_114_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_624 ();
 DECAPx4_ASAP7_75t_R FILLER_114_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_655 ();
 DECAPx1_ASAP7_75t_R FILLER_114_663 ();
 FILLER_ASAP7_75t_R FILLER_114_689 ();
 DECAPx2_ASAP7_75t_R FILLER_114_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_703 ();
 DECAPx10_ASAP7_75t_R FILLER_114_714 ();
 DECAPx1_ASAP7_75t_R FILLER_114_736 ();
 DECAPx6_ASAP7_75t_R FILLER_114_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_766 ();
 DECAPx10_ASAP7_75t_R FILLER_114_770 ();
 DECAPx10_ASAP7_75t_R FILLER_114_792 ();
 DECAPx2_ASAP7_75t_R FILLER_114_814 ();
 FILLER_ASAP7_75t_R FILLER_114_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_822 ();
 DECAPx4_ASAP7_75t_R FILLER_114_839 ();
 DECAPx10_ASAP7_75t_R FILLER_114_859 ();
 DECAPx4_ASAP7_75t_R FILLER_114_903 ();
 FILLER_ASAP7_75t_R FILLER_114_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_915 ();
 FILLER_ASAP7_75t_R FILLER_114_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_936 ();
 DECAPx10_ASAP7_75t_R FILLER_114_943 ();
 DECAPx2_ASAP7_75t_R FILLER_114_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_971 ();
 DECAPx2_ASAP7_75t_R FILLER_114_983 ();
 FILLER_ASAP7_75t_R FILLER_114_989 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1146 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1182 ();
 FILLER_ASAP7_75t_R FILLER_114_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1277 ();
 FILLER_ASAP7_75t_R FILLER_114_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_115_512 ();
 FILLER_ASAP7_75t_R FILLER_115_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_536 ();
 DECAPx10_ASAP7_75t_R FILLER_115_547 ();
 FILLER_ASAP7_75t_R FILLER_115_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_584 ();
 DECAPx10_ASAP7_75t_R FILLER_115_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_631 ();
 DECAPx1_ASAP7_75t_R FILLER_115_650 ();
 FILLER_ASAP7_75t_R FILLER_115_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_670 ();
 FILLER_ASAP7_75t_R FILLER_115_674 ();
 DECAPx2_ASAP7_75t_R FILLER_115_682 ();
 FILLER_ASAP7_75t_R FILLER_115_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_690 ();
 FILLER_ASAP7_75t_R FILLER_115_697 ();
 FILLER_ASAP7_75t_R FILLER_115_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_707 ();
 DECAPx1_ASAP7_75t_R FILLER_115_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_722 ();
 DECAPx2_ASAP7_75t_R FILLER_115_737 ();
 FILLER_ASAP7_75t_R FILLER_115_743 ();
 FILLER_ASAP7_75t_R FILLER_115_772 ();
 DECAPx10_ASAP7_75t_R FILLER_115_780 ();
 DECAPx10_ASAP7_75t_R FILLER_115_802 ();
 DECAPx2_ASAP7_75t_R FILLER_115_824 ();
 FILLER_ASAP7_75t_R FILLER_115_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_832 ();
 DECAPx10_ASAP7_75t_R FILLER_115_843 ();
 DECAPx10_ASAP7_75t_R FILLER_115_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_917 ();
 DECAPx10_ASAP7_75t_R FILLER_115_928 ();
 DECAPx4_ASAP7_75t_R FILLER_115_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_960 ();
 DECAPx10_ASAP7_75t_R FILLER_115_967 ();
 DECAPx10_ASAP7_75t_R FILLER_115_989 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1055 ();
 FILLER_ASAP7_75t_R FILLER_115_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1075 ();
 FILLER_ASAP7_75t_R FILLER_115_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1087 ();
 FILLER_ASAP7_75t_R FILLER_115_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1210 ();
 FILLER_ASAP7_75t_R FILLER_115_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1233 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1255 ();
 FILLER_ASAP7_75t_R FILLER_115_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1271 ();
 DECAPx1_ASAP7_75t_R FILLER_116_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_516 ();
 DECAPx10_ASAP7_75t_R FILLER_116_523 ();
 DECAPx6_ASAP7_75t_R FILLER_116_570 ();
 DECAPx2_ASAP7_75t_R FILLER_116_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_590 ();
 DECAPx6_ASAP7_75t_R FILLER_116_599 ();
 DECAPx2_ASAP7_75t_R FILLER_116_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_619 ();
 DECAPx10_ASAP7_75t_R FILLER_116_649 ();
 DECAPx6_ASAP7_75t_R FILLER_116_671 ();
 DECAPx1_ASAP7_75t_R FILLER_116_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_696 ();
 DECAPx10_ASAP7_75t_R FILLER_116_705 ();
 DECAPx10_ASAP7_75t_R FILLER_116_727 ();
 DECAPx10_ASAP7_75t_R FILLER_116_749 ();
 DECAPx1_ASAP7_75t_R FILLER_116_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_775 ();
 DECAPx10_ASAP7_75t_R FILLER_116_786 ();
 DECAPx6_ASAP7_75t_R FILLER_116_808 ();
 DECAPx2_ASAP7_75t_R FILLER_116_822 ();
 DECAPx10_ASAP7_75t_R FILLER_116_840 ();
 DECAPx10_ASAP7_75t_R FILLER_116_862 ();
 FILLER_ASAP7_75t_R FILLER_116_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_886 ();
 DECAPx10_ASAP7_75t_R FILLER_116_909 ();
 DECAPx10_ASAP7_75t_R FILLER_116_931 ();
 DECAPx6_ASAP7_75t_R FILLER_116_953 ();
 DECAPx1_ASAP7_75t_R FILLER_116_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_971 ();
 DECAPx10_ASAP7_75t_R FILLER_116_974 ();
 DECAPx10_ASAP7_75t_R FILLER_116_996 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1040 ();
 FILLER_ASAP7_75t_R FILLER_116_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1055 ();
 FILLER_ASAP7_75t_R FILLER_116_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1104 ();
 FILLER_ASAP7_75t_R FILLER_116_1114 ();
 FILLER_ASAP7_75t_R FILLER_116_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_116_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1280 ();
 FILLER_ASAP7_75t_R FILLER_116_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_117_2 ();
 DECAPx10_ASAP7_75t_R FILLER_117_24 ();
 DECAPx10_ASAP7_75t_R FILLER_117_46 ();
 DECAPx10_ASAP7_75t_R FILLER_117_68 ();
 DECAPx10_ASAP7_75t_R FILLER_117_90 ();
 DECAPx10_ASAP7_75t_R FILLER_117_112 ();
 DECAPx10_ASAP7_75t_R FILLER_117_134 ();
 DECAPx10_ASAP7_75t_R FILLER_117_156 ();
 DECAPx10_ASAP7_75t_R FILLER_117_178 ();
 DECAPx10_ASAP7_75t_R FILLER_117_200 ();
 DECAPx10_ASAP7_75t_R FILLER_117_222 ();
 DECAPx10_ASAP7_75t_R FILLER_117_244 ();
 DECAPx10_ASAP7_75t_R FILLER_117_266 ();
 DECAPx10_ASAP7_75t_R FILLER_117_288 ();
 DECAPx10_ASAP7_75t_R FILLER_117_310 ();
 DECAPx10_ASAP7_75t_R FILLER_117_332 ();
 DECAPx10_ASAP7_75t_R FILLER_117_354 ();
 DECAPx10_ASAP7_75t_R FILLER_117_376 ();
 DECAPx10_ASAP7_75t_R FILLER_117_398 ();
 DECAPx10_ASAP7_75t_R FILLER_117_420 ();
 DECAPx6_ASAP7_75t_R FILLER_117_442 ();
 DECAPx2_ASAP7_75t_R FILLER_117_456 ();
 DECAPx10_ASAP7_75t_R FILLER_117_464 ();
 DECAPx10_ASAP7_75t_R FILLER_117_486 ();
 DECAPx4_ASAP7_75t_R FILLER_117_508 ();
 DECAPx6_ASAP7_75t_R FILLER_117_528 ();
 DECAPx2_ASAP7_75t_R FILLER_117_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_548 ();
 DECAPx10_ASAP7_75t_R FILLER_117_570 ();
 DECAPx10_ASAP7_75t_R FILLER_117_592 ();
 DECAPx6_ASAP7_75t_R FILLER_117_614 ();
 FILLER_ASAP7_75t_R FILLER_117_628 ();
 DECAPx10_ASAP7_75t_R FILLER_117_640 ();
 DECAPx10_ASAP7_75t_R FILLER_117_662 ();
 DECAPx10_ASAP7_75t_R FILLER_117_684 ();
 DECAPx6_ASAP7_75t_R FILLER_117_706 ();
 DECAPx1_ASAP7_75t_R FILLER_117_720 ();
 DECAPx10_ASAP7_75t_R FILLER_117_738 ();
 DECAPx10_ASAP7_75t_R FILLER_117_760 ();
 DECAPx10_ASAP7_75t_R FILLER_117_782 ();
 DECAPx4_ASAP7_75t_R FILLER_117_804 ();
 FILLER_ASAP7_75t_R FILLER_117_814 ();
 DECAPx4_ASAP7_75t_R FILLER_117_832 ();
 FILLER_ASAP7_75t_R FILLER_117_842 ();
 DECAPx4_ASAP7_75t_R FILLER_117_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_864 ();
 DECAPx10_ASAP7_75t_R FILLER_117_881 ();
 DECAPx6_ASAP7_75t_R FILLER_117_903 ();
 DECAPx2_ASAP7_75t_R FILLER_117_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_923 ();
 FILLER_ASAP7_75t_R FILLER_117_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_928 ();
 DECAPx4_ASAP7_75t_R FILLER_117_937 ();
 FILLER_ASAP7_75t_R FILLER_117_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_955 ();
 DECAPx6_ASAP7_75t_R FILLER_117_962 ();
 DECAPx1_ASAP7_75t_R FILLER_117_976 ();
 FILLER_ASAP7_75t_R FILLER_117_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_989 ();
 DECAPx10_ASAP7_75t_R FILLER_117_996 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1040 ();
 FILLER_ASAP7_75t_R FILLER_117_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1103 ();
 FILLER_ASAP7_75t_R FILLER_117_1113 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1121 ();
 FILLER_ASAP7_75t_R FILLER_117_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1162 ();
 FILLER_ASAP7_75t_R FILLER_117_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1174 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_118_2 ();
 DECAPx10_ASAP7_75t_R FILLER_118_24 ();
 DECAPx10_ASAP7_75t_R FILLER_118_46 ();
 DECAPx10_ASAP7_75t_R FILLER_118_68 ();
 DECAPx10_ASAP7_75t_R FILLER_118_90 ();
 DECAPx10_ASAP7_75t_R FILLER_118_112 ();
 DECAPx10_ASAP7_75t_R FILLER_118_134 ();
 DECAPx10_ASAP7_75t_R FILLER_118_156 ();
 DECAPx10_ASAP7_75t_R FILLER_118_178 ();
 DECAPx10_ASAP7_75t_R FILLER_118_200 ();
 DECAPx10_ASAP7_75t_R FILLER_118_222 ();
 DECAPx10_ASAP7_75t_R FILLER_118_244 ();
 DECAPx10_ASAP7_75t_R FILLER_118_266 ();
 DECAPx10_ASAP7_75t_R FILLER_118_288 ();
 DECAPx10_ASAP7_75t_R FILLER_118_310 ();
 DECAPx10_ASAP7_75t_R FILLER_118_332 ();
 DECAPx10_ASAP7_75t_R FILLER_118_354 ();
 DECAPx10_ASAP7_75t_R FILLER_118_376 ();
 DECAPx10_ASAP7_75t_R FILLER_118_398 ();
 DECAPx10_ASAP7_75t_R FILLER_118_420 ();
 DECAPx6_ASAP7_75t_R FILLER_118_442 ();
 DECAPx2_ASAP7_75t_R FILLER_118_456 ();
 DECAPx10_ASAP7_75t_R FILLER_118_464 ();
 DECAPx6_ASAP7_75t_R FILLER_118_486 ();
 DECAPx1_ASAP7_75t_R FILLER_118_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_530 ();
 DECAPx10_ASAP7_75t_R FILLER_118_541 ();
 DECAPx2_ASAP7_75t_R FILLER_118_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_569 ();
 DECAPx1_ASAP7_75t_R FILLER_118_584 ();
 DECAPx4_ASAP7_75t_R FILLER_118_594 ();
 FILLER_ASAP7_75t_R FILLER_118_604 ();
 DECAPx10_ASAP7_75t_R FILLER_118_612 ();
 DECAPx2_ASAP7_75t_R FILLER_118_634 ();
 FILLER_ASAP7_75t_R FILLER_118_640 ();
 DECAPx10_ASAP7_75t_R FILLER_118_660 ();
 DECAPx10_ASAP7_75t_R FILLER_118_682 ();
 DECAPx10_ASAP7_75t_R FILLER_118_704 ();
 DECAPx6_ASAP7_75t_R FILLER_118_726 ();
 DECAPx1_ASAP7_75t_R FILLER_118_740 ();
 DECAPx10_ASAP7_75t_R FILLER_118_753 ();
 DECAPx10_ASAP7_75t_R FILLER_118_775 ();
 DECAPx10_ASAP7_75t_R FILLER_118_797 ();
 DECAPx2_ASAP7_75t_R FILLER_118_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_825 ();
 DECAPx10_ASAP7_75t_R FILLER_118_836 ();
 DECAPx10_ASAP7_75t_R FILLER_118_858 ();
 DECAPx10_ASAP7_75t_R FILLER_118_880 ();
 DECAPx10_ASAP7_75t_R FILLER_118_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_924 ();
 DECAPx10_ASAP7_75t_R FILLER_118_952 ();
 DECAPx10_ASAP7_75t_R FILLER_118_974 ();
 DECAPx4_ASAP7_75t_R FILLER_118_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1006 ();
 FILLER_ASAP7_75t_R FILLER_118_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1280 ();
 FILLER_ASAP7_75t_R FILLER_118_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_119_2 ();
 DECAPx10_ASAP7_75t_R FILLER_119_24 ();
 DECAPx10_ASAP7_75t_R FILLER_119_46 ();
 DECAPx10_ASAP7_75t_R FILLER_119_68 ();
 DECAPx10_ASAP7_75t_R FILLER_119_90 ();
 DECAPx6_ASAP7_75t_R FILLER_119_112 ();
 DECAPx1_ASAP7_75t_R FILLER_119_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_130 ();
 DECAPx10_ASAP7_75t_R FILLER_119_171 ();
 DECAPx10_ASAP7_75t_R FILLER_119_193 ();
 DECAPx10_ASAP7_75t_R FILLER_119_215 ();
 DECAPx10_ASAP7_75t_R FILLER_119_237 ();
 DECAPx10_ASAP7_75t_R FILLER_119_259 ();
 DECAPx2_ASAP7_75t_R FILLER_119_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_300 ();
 DECAPx10_ASAP7_75t_R FILLER_119_307 ();
 DECAPx10_ASAP7_75t_R FILLER_119_329 ();
 DECAPx10_ASAP7_75t_R FILLER_119_351 ();
 DECAPx10_ASAP7_75t_R FILLER_119_373 ();
 DECAPx10_ASAP7_75t_R FILLER_119_395 ();
 DECAPx2_ASAP7_75t_R FILLER_119_417 ();
 DECAPx1_ASAP7_75t_R FILLER_119_434 ();
 DECAPx1_ASAP7_75t_R FILLER_119_444 ();
 DECAPx10_ASAP7_75t_R FILLER_119_464 ();
 DECAPx10_ASAP7_75t_R FILLER_119_486 ();
 DECAPx2_ASAP7_75t_R FILLER_119_508 ();
 FILLER_ASAP7_75t_R FILLER_119_514 ();
 DECAPx6_ASAP7_75t_R FILLER_119_526 ();
 DECAPx2_ASAP7_75t_R FILLER_119_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_554 ();
 DECAPx6_ASAP7_75t_R FILLER_119_561 ();
 DECAPx2_ASAP7_75t_R FILLER_119_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_581 ();
 DECAPx1_ASAP7_75t_R FILLER_119_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_597 ();
 DECAPx4_ASAP7_75t_R FILLER_119_604 ();
 FILLER_ASAP7_75t_R FILLER_119_614 ();
 DECAPx2_ASAP7_75t_R FILLER_119_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_661 ();
 DECAPx1_ASAP7_75t_R FILLER_119_665 ();
 DECAPx6_ASAP7_75t_R FILLER_119_675 ();
 DECAPx1_ASAP7_75t_R FILLER_119_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_693 ();
 FILLER_ASAP7_75t_R FILLER_119_704 ();
 DECAPx10_ASAP7_75t_R FILLER_119_716 ();
 FILLER_ASAP7_75t_R FILLER_119_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_740 ();
 DECAPx10_ASAP7_75t_R FILLER_119_750 ();
 DECAPx1_ASAP7_75t_R FILLER_119_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_776 ();
 DECAPx10_ASAP7_75t_R FILLER_119_786 ();
 DECAPx10_ASAP7_75t_R FILLER_119_808 ();
 DECAPx10_ASAP7_75t_R FILLER_119_830 ();
 DECAPx4_ASAP7_75t_R FILLER_119_858 ();
 FILLER_ASAP7_75t_R FILLER_119_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_870 ();
 FILLER_ASAP7_75t_R FILLER_119_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_889 ();
 DECAPx6_ASAP7_75t_R FILLER_119_899 ();
 FILLER_ASAP7_75t_R FILLER_119_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_923 ();
 DECAPx2_ASAP7_75t_R FILLER_119_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_932 ();
 DECAPx10_ASAP7_75t_R FILLER_119_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_961 ();
 DECAPx10_ASAP7_75t_R FILLER_119_970 ();
 DECAPx4_ASAP7_75t_R FILLER_119_992 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1074 ();
 FILLER_ASAP7_75t_R FILLER_119_1084 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1200 ();
 FILLER_ASAP7_75t_R FILLER_119_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1248 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_120_2 ();
 DECAPx10_ASAP7_75t_R FILLER_120_24 ();
 DECAPx10_ASAP7_75t_R FILLER_120_46 ();
 DECAPx10_ASAP7_75t_R FILLER_120_68 ();
 DECAPx10_ASAP7_75t_R FILLER_120_90 ();
 DECAPx1_ASAP7_75t_R FILLER_120_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_116 ();
 FILLER_ASAP7_75t_R FILLER_120_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_127 ();
 DECAPx1_ASAP7_75t_R FILLER_120_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_140 ();
 DECAPx6_ASAP7_75t_R FILLER_120_149 ();
 FILLER_ASAP7_75t_R FILLER_120_163 ();
 DECAPx1_ASAP7_75t_R FILLER_120_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_177 ();
 DECAPx10_ASAP7_75t_R FILLER_120_186 ();
 DECAPx10_ASAP7_75t_R FILLER_120_208 ();
 DECAPx10_ASAP7_75t_R FILLER_120_230 ();
 DECAPx6_ASAP7_75t_R FILLER_120_252 ();
 DECAPx10_ASAP7_75t_R FILLER_120_272 ();
 DECAPx6_ASAP7_75t_R FILLER_120_312 ();
 DECAPx2_ASAP7_75t_R FILLER_120_326 ();
 DECAPx10_ASAP7_75t_R FILLER_120_338 ();
 DECAPx10_ASAP7_75t_R FILLER_120_360 ();
 DECAPx10_ASAP7_75t_R FILLER_120_382 ();
 DECAPx1_ASAP7_75t_R FILLER_120_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_408 ();
 FILLER_ASAP7_75t_R FILLER_120_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_453 ();
 DECAPx10_ASAP7_75t_R FILLER_120_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_486 ();
 FILLER_ASAP7_75t_R FILLER_120_511 ();
 DECAPx2_ASAP7_75t_R FILLER_120_522 ();
 FILLER_ASAP7_75t_R FILLER_120_528 ();
 DECAPx4_ASAP7_75t_R FILLER_120_538 ();
 FILLER_ASAP7_75t_R FILLER_120_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_550 ();
 DECAPx4_ASAP7_75t_R FILLER_120_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_575 ();
 DECAPx10_ASAP7_75t_R FILLER_120_597 ();
 DECAPx1_ASAP7_75t_R FILLER_120_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_623 ();
 DECAPx2_ASAP7_75t_R FILLER_120_631 ();
 DECAPx10_ASAP7_75t_R FILLER_120_643 ();
 FILLER_ASAP7_75t_R FILLER_120_665 ();
 DECAPx2_ASAP7_75t_R FILLER_120_676 ();
 FILLER_ASAP7_75t_R FILLER_120_682 ();
 DECAPx10_ASAP7_75t_R FILLER_120_690 ();
 DECAPx6_ASAP7_75t_R FILLER_120_712 ();
 FILLER_ASAP7_75t_R FILLER_120_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_728 ();
 DECAPx10_ASAP7_75t_R FILLER_120_739 ();
 DECAPx6_ASAP7_75t_R FILLER_120_761 ();
 DECAPx1_ASAP7_75t_R FILLER_120_775 ();
 DECAPx10_ASAP7_75t_R FILLER_120_793 ();
 DECAPx10_ASAP7_75t_R FILLER_120_815 ();
 DECAPx10_ASAP7_75t_R FILLER_120_837 ();
 DECAPx10_ASAP7_75t_R FILLER_120_859 ();
 DECAPx6_ASAP7_75t_R FILLER_120_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_895 ();
 DECAPx10_ASAP7_75t_R FILLER_120_906 ();
 DECAPx10_ASAP7_75t_R FILLER_120_928 ();
 DECAPx4_ASAP7_75t_R FILLER_120_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_960 ();
 DECAPx2_ASAP7_75t_R FILLER_120_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_988 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1093 ();
 FILLER_ASAP7_75t_R FILLER_120_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1119 ();
 FILLER_ASAP7_75t_R FILLER_120_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1127 ();
 FILLER_ASAP7_75t_R FILLER_120_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_121_2 ();
 DECAPx10_ASAP7_75t_R FILLER_121_24 ();
 DECAPx10_ASAP7_75t_R FILLER_121_46 ();
 DECAPx10_ASAP7_75t_R FILLER_121_68 ();
 DECAPx10_ASAP7_75t_R FILLER_121_90 ();
 DECAPx6_ASAP7_75t_R FILLER_121_112 ();
 FILLER_ASAP7_75t_R FILLER_121_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_144 ();
 DECAPx10_ASAP7_75t_R FILLER_121_153 ();
 DECAPx10_ASAP7_75t_R FILLER_121_175 ();
 DECAPx6_ASAP7_75t_R FILLER_121_197 ();
 DECAPx2_ASAP7_75t_R FILLER_121_211 ();
 DECAPx6_ASAP7_75t_R FILLER_121_223 ();
 FILLER_ASAP7_75t_R FILLER_121_237 ();
 DECAPx6_ASAP7_75t_R FILLER_121_245 ();
 FILLER_ASAP7_75t_R FILLER_121_259 ();
 DECAPx10_ASAP7_75t_R FILLER_121_267 ();
 DECAPx2_ASAP7_75t_R FILLER_121_289 ();
 FILLER_ASAP7_75t_R FILLER_121_295 ();
 DECAPx10_ASAP7_75t_R FILLER_121_309 ();
 DECAPx2_ASAP7_75t_R FILLER_121_331 ();
 DECAPx4_ASAP7_75t_R FILLER_121_347 ();
 FILLER_ASAP7_75t_R FILLER_121_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_376 ();
 DECAPx2_ASAP7_75t_R FILLER_121_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_449 ();
 DECAPx6_ASAP7_75t_R FILLER_121_468 ();
 DECAPx1_ASAP7_75t_R FILLER_121_482 ();
 FILLER_ASAP7_75t_R FILLER_121_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_491 ();
 FILLER_ASAP7_75t_R FILLER_121_514 ();
 DECAPx2_ASAP7_75t_R FILLER_121_523 ();
 FILLER_ASAP7_75t_R FILLER_121_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_531 ();
 DECAPx6_ASAP7_75t_R FILLER_121_539 ();
 DECAPx4_ASAP7_75t_R FILLER_121_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_569 ();
 DECAPx6_ASAP7_75t_R FILLER_121_580 ();
 FILLER_ASAP7_75t_R FILLER_121_594 ();
 DECAPx6_ASAP7_75t_R FILLER_121_602 ();
 FILLER_ASAP7_75t_R FILLER_121_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_628 ();
 DECAPx10_ASAP7_75t_R FILLER_121_641 ();
 DECAPx6_ASAP7_75t_R FILLER_121_663 ();
 DECAPx1_ASAP7_75t_R FILLER_121_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_681 ();
 DECAPx10_ASAP7_75t_R FILLER_121_694 ();
 DECAPx10_ASAP7_75t_R FILLER_121_716 ();
 DECAPx10_ASAP7_75t_R FILLER_121_738 ();
 DECAPx10_ASAP7_75t_R FILLER_121_760 ();
 DECAPx10_ASAP7_75t_R FILLER_121_782 ();
 DECAPx6_ASAP7_75t_R FILLER_121_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_818 ();
 DECAPx10_ASAP7_75t_R FILLER_121_831 ();
 DECAPx10_ASAP7_75t_R FILLER_121_853 ();
 DECAPx10_ASAP7_75t_R FILLER_121_875 ();
 DECAPx10_ASAP7_75t_R FILLER_121_897 ();
 DECAPx1_ASAP7_75t_R FILLER_121_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_923 ();
 DECAPx10_ASAP7_75t_R FILLER_121_926 ();
 DECAPx6_ASAP7_75t_R FILLER_121_948 ();
 DECAPx10_ASAP7_75t_R FILLER_121_968 ();
 DECAPx10_ASAP7_75t_R FILLER_121_996 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1018 ();
 FILLER_ASAP7_75t_R FILLER_121_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1084 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1217 ();
 DECAPx6_ASAP7_75t_R FILLER_121_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_122_2 ();
 DECAPx10_ASAP7_75t_R FILLER_122_24 ();
 DECAPx10_ASAP7_75t_R FILLER_122_46 ();
 DECAPx10_ASAP7_75t_R FILLER_122_68 ();
 DECAPx10_ASAP7_75t_R FILLER_122_90 ();
 DECAPx10_ASAP7_75t_R FILLER_122_112 ();
 DECAPx10_ASAP7_75t_R FILLER_122_134 ();
 DECAPx10_ASAP7_75t_R FILLER_122_156 ();
 DECAPx10_ASAP7_75t_R FILLER_122_178 ();
 DECAPx10_ASAP7_75t_R FILLER_122_200 ();
 DECAPx10_ASAP7_75t_R FILLER_122_222 ();
 DECAPx10_ASAP7_75t_R FILLER_122_244 ();
 DECAPx10_ASAP7_75t_R FILLER_122_266 ();
 DECAPx6_ASAP7_75t_R FILLER_122_288 ();
 DECAPx2_ASAP7_75t_R FILLER_122_302 ();
 DECAPx10_ASAP7_75t_R FILLER_122_318 ();
 DECAPx10_ASAP7_75t_R FILLER_122_340 ();
 DECAPx10_ASAP7_75t_R FILLER_122_362 ();
 DECAPx10_ASAP7_75t_R FILLER_122_384 ();
 DECAPx2_ASAP7_75t_R FILLER_122_406 ();
 FILLER_ASAP7_75t_R FILLER_122_412 ();
 DECAPx1_ASAP7_75t_R FILLER_122_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_427 ();
 DECAPx1_ASAP7_75t_R FILLER_122_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_445 ();
 DECAPx4_ASAP7_75t_R FILLER_122_449 ();
 FILLER_ASAP7_75t_R FILLER_122_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_461 ();
 DECAPx6_ASAP7_75t_R FILLER_122_464 ();
 DECAPx2_ASAP7_75t_R FILLER_122_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_491 ();
 DECAPx2_ASAP7_75t_R FILLER_122_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_521 ();
 FILLER_ASAP7_75t_R FILLER_122_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_534 ();
 DECAPx6_ASAP7_75t_R FILLER_122_557 ();
 DECAPx1_ASAP7_75t_R FILLER_122_571 ();
 DECAPx10_ASAP7_75t_R FILLER_122_581 ();
 DECAPx10_ASAP7_75t_R FILLER_122_603 ();
 DECAPx10_ASAP7_75t_R FILLER_122_625 ();
 DECAPx10_ASAP7_75t_R FILLER_122_647 ();
 DECAPx10_ASAP7_75t_R FILLER_122_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_698 ();
 DECAPx1_ASAP7_75t_R FILLER_122_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_727 ();
 DECAPx10_ASAP7_75t_R FILLER_122_736 ();
 DECAPx10_ASAP7_75t_R FILLER_122_758 ();
 DECAPx10_ASAP7_75t_R FILLER_122_780 ();
 DECAPx6_ASAP7_75t_R FILLER_122_802 ();
 DECAPx2_ASAP7_75t_R FILLER_122_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_822 ();
 DECAPx6_ASAP7_75t_R FILLER_122_841 ();
 DECAPx1_ASAP7_75t_R FILLER_122_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_859 ();
 DECAPx6_ASAP7_75t_R FILLER_122_874 ();
 FILLER_ASAP7_75t_R FILLER_122_888 ();
 DECAPx4_ASAP7_75t_R FILLER_122_896 ();
 FILLER_ASAP7_75t_R FILLER_122_906 ();
 DECAPx4_ASAP7_75t_R FILLER_122_922 ();
 FILLER_ASAP7_75t_R FILLER_122_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_934 ();
 DECAPx1_ASAP7_75t_R FILLER_122_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_953 ();
 DECAPx10_ASAP7_75t_R FILLER_122_960 ();
 DECAPx10_ASAP7_75t_R FILLER_122_982 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1004 ();
 FILLER_ASAP7_75t_R FILLER_122_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_122_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1241 ();
 FILLER_ASAP7_75t_R FILLER_122_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1277 ();
 FILLER_ASAP7_75t_R FILLER_122_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_123_24 ();
 DECAPx10_ASAP7_75t_R FILLER_123_46 ();
 DECAPx10_ASAP7_75t_R FILLER_123_68 ();
 DECAPx10_ASAP7_75t_R FILLER_123_90 ();
 DECAPx6_ASAP7_75t_R FILLER_123_112 ();
 DECAPx1_ASAP7_75t_R FILLER_123_126 ();
 DECAPx6_ASAP7_75t_R FILLER_123_154 ();
 DECAPx1_ASAP7_75t_R FILLER_123_168 ();
 DECAPx10_ASAP7_75t_R FILLER_123_180 ();
 DECAPx10_ASAP7_75t_R FILLER_123_202 ();
 DECAPx10_ASAP7_75t_R FILLER_123_224 ();
 DECAPx2_ASAP7_75t_R FILLER_123_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_252 ();
 DECAPx6_ASAP7_75t_R FILLER_123_259 ();
 DECAPx2_ASAP7_75t_R FILLER_123_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_279 ();
 DECAPx2_ASAP7_75t_R FILLER_123_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_307 ();
 DECAPx10_ASAP7_75t_R FILLER_123_318 ();
 DECAPx10_ASAP7_75t_R FILLER_123_340 ();
 DECAPx10_ASAP7_75t_R FILLER_123_362 ();
 DECAPx10_ASAP7_75t_R FILLER_123_384 ();
 DECAPx4_ASAP7_75t_R FILLER_123_406 ();
 FILLER_ASAP7_75t_R FILLER_123_416 ();
 DECAPx2_ASAP7_75t_R FILLER_123_426 ();
 FILLER_ASAP7_75t_R FILLER_123_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_434 ();
 FILLER_ASAP7_75t_R FILLER_123_442 ();
 DECAPx10_ASAP7_75t_R FILLER_123_455 ();
 DECAPx10_ASAP7_75t_R FILLER_123_487 ();
 DECAPx2_ASAP7_75t_R FILLER_123_509 ();
 DECAPx2_ASAP7_75t_R FILLER_123_522 ();
 FILLER_ASAP7_75t_R FILLER_123_528 ();
 DECAPx6_ASAP7_75t_R FILLER_123_536 ();
 FILLER_ASAP7_75t_R FILLER_123_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_552 ();
 DECAPx4_ASAP7_75t_R FILLER_123_559 ();
 FILLER_ASAP7_75t_R FILLER_123_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_571 ();
 DECAPx6_ASAP7_75t_R FILLER_123_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_603 ();
 DECAPx10_ASAP7_75t_R FILLER_123_610 ();
 DECAPx6_ASAP7_75t_R FILLER_123_632 ();
 DECAPx10_ASAP7_75t_R FILLER_123_653 ();
 DECAPx10_ASAP7_75t_R FILLER_123_675 ();
 DECAPx10_ASAP7_75t_R FILLER_123_697 ();
 DECAPx4_ASAP7_75t_R FILLER_123_719 ();
 FILLER_ASAP7_75t_R FILLER_123_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_731 ();
 FILLER_ASAP7_75t_R FILLER_123_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_747 ();
 DECAPx10_ASAP7_75t_R FILLER_123_754 ();
 DECAPx6_ASAP7_75t_R FILLER_123_776 ();
 DECAPx2_ASAP7_75t_R FILLER_123_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_796 ();
 FILLER_ASAP7_75t_R FILLER_123_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_813 ();
 DECAPx10_ASAP7_75t_R FILLER_123_834 ();
 DECAPx4_ASAP7_75t_R FILLER_123_856 ();
 DECAPx10_ASAP7_75t_R FILLER_123_872 ();
 DECAPx10_ASAP7_75t_R FILLER_123_894 ();
 DECAPx2_ASAP7_75t_R FILLER_123_916 ();
 FILLER_ASAP7_75t_R FILLER_123_922 ();
 DECAPx10_ASAP7_75t_R FILLER_123_926 ();
 DECAPx6_ASAP7_75t_R FILLER_123_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_962 ();
 DECAPx1_ASAP7_75t_R FILLER_123_969 ();
 DECAPx10_ASAP7_75t_R FILLER_123_983 ();
 FILLER_ASAP7_75t_R FILLER_123_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1041 ();
 FILLER_ASAP7_75t_R FILLER_123_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1097 ();
 FILLER_ASAP7_75t_R FILLER_123_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1213 ();
 FILLER_ASAP7_75t_R FILLER_123_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1247 ();
 FILLER_ASAP7_75t_R FILLER_123_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_124_2 ();
 DECAPx10_ASAP7_75t_R FILLER_124_24 ();
 DECAPx10_ASAP7_75t_R FILLER_124_46 ();
 DECAPx10_ASAP7_75t_R FILLER_124_68 ();
 DECAPx10_ASAP7_75t_R FILLER_124_90 ();
 FILLER_ASAP7_75t_R FILLER_124_112 ();
 DECAPx6_ASAP7_75t_R FILLER_124_120 ();
 DECAPx2_ASAP7_75t_R FILLER_124_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_140 ();
 DECAPx10_ASAP7_75t_R FILLER_124_149 ();
 DECAPx4_ASAP7_75t_R FILLER_124_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_181 ();
 DECAPx10_ASAP7_75t_R FILLER_124_190 ();
 FILLER_ASAP7_75t_R FILLER_124_212 ();
 DECAPx4_ASAP7_75t_R FILLER_124_220 ();
 DECAPx10_ASAP7_75t_R FILLER_124_236 ();
 DECAPx10_ASAP7_75t_R FILLER_124_258 ();
 DECAPx2_ASAP7_75t_R FILLER_124_280 ();
 DECAPx2_ASAP7_75t_R FILLER_124_292 ();
 DECAPx6_ASAP7_75t_R FILLER_124_308 ();
 DECAPx2_ASAP7_75t_R FILLER_124_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_328 ();
 DECAPx10_ASAP7_75t_R FILLER_124_335 ();
 FILLER_ASAP7_75t_R FILLER_124_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_359 ();
 DECAPx10_ASAP7_75t_R FILLER_124_376 ();
 DECAPx6_ASAP7_75t_R FILLER_124_398 ();
 DECAPx2_ASAP7_75t_R FILLER_124_412 ();
 DECAPx2_ASAP7_75t_R FILLER_124_426 ();
 FILLER_ASAP7_75t_R FILLER_124_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_441 ();
 DECAPx1_ASAP7_75t_R FILLER_124_458 ();
 DECAPx2_ASAP7_75t_R FILLER_124_464 ();
 FILLER_ASAP7_75t_R FILLER_124_470 ();
 DECAPx4_ASAP7_75t_R FILLER_124_496 ();
 FILLER_ASAP7_75t_R FILLER_124_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_508 ();
 FILLER_ASAP7_75t_R FILLER_124_516 ();
 DECAPx2_ASAP7_75t_R FILLER_124_553 ();
 FILLER_ASAP7_75t_R FILLER_124_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_561 ();
 DECAPx10_ASAP7_75t_R FILLER_124_583 ();
 FILLER_ASAP7_75t_R FILLER_124_605 ();
 DECAPx6_ASAP7_75t_R FILLER_124_615 ();
 DECAPx6_ASAP7_75t_R FILLER_124_638 ();
 FILLER_ASAP7_75t_R FILLER_124_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_654 ();
 DECAPx2_ASAP7_75t_R FILLER_124_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_679 ();
 DECAPx10_ASAP7_75t_R FILLER_124_686 ();
 DECAPx10_ASAP7_75t_R FILLER_124_708 ();
 DECAPx2_ASAP7_75t_R FILLER_124_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_736 ();
 FILLER_ASAP7_75t_R FILLER_124_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_751 ();
 DECAPx10_ASAP7_75t_R FILLER_124_758 ();
 DECAPx1_ASAP7_75t_R FILLER_124_780 ();
 DECAPx4_ASAP7_75t_R FILLER_124_787 ();
 FILLER_ASAP7_75t_R FILLER_124_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_815 ();
 DECAPx10_ASAP7_75t_R FILLER_124_822 ();
 DECAPx10_ASAP7_75t_R FILLER_124_844 ();
 DECAPx10_ASAP7_75t_R FILLER_124_866 ();
 DECAPx10_ASAP7_75t_R FILLER_124_894 ();
 DECAPx10_ASAP7_75t_R FILLER_124_916 ();
 DECAPx10_ASAP7_75t_R FILLER_124_938 ();
 DECAPx10_ASAP7_75t_R FILLER_124_960 ();
 DECAPx2_ASAP7_75t_R FILLER_124_982 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1061 ();
 FILLER_ASAP7_75t_R FILLER_124_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1096 ();
 FILLER_ASAP7_75t_R FILLER_124_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1231 ();
 FILLER_ASAP7_75t_R FILLER_124_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1258 ();
 FILLER_ASAP7_75t_R FILLER_124_1264 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1280 ();
 FILLER_ASAP7_75t_R FILLER_124_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_125_2 ();
 DECAPx10_ASAP7_75t_R FILLER_125_24 ();
 DECAPx10_ASAP7_75t_R FILLER_125_46 ();
 DECAPx10_ASAP7_75t_R FILLER_125_68 ();
 DECAPx10_ASAP7_75t_R FILLER_125_90 ();
 DECAPx6_ASAP7_75t_R FILLER_125_112 ();
 DECAPx2_ASAP7_75t_R FILLER_125_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_132 ();
 DECAPx10_ASAP7_75t_R FILLER_125_147 ();
 DECAPx10_ASAP7_75t_R FILLER_125_169 ();
 DECAPx10_ASAP7_75t_R FILLER_125_191 ();
 DECAPx10_ASAP7_75t_R FILLER_125_213 ();
 DECAPx2_ASAP7_75t_R FILLER_125_235 ();
 FILLER_ASAP7_75t_R FILLER_125_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_243 ();
 DECAPx10_ASAP7_75t_R FILLER_125_250 ();
 DECAPx2_ASAP7_75t_R FILLER_125_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_278 ();
 DECAPx2_ASAP7_75t_R FILLER_125_289 ();
 DECAPx10_ASAP7_75t_R FILLER_125_315 ();
 DECAPx10_ASAP7_75t_R FILLER_125_337 ();
 DECAPx1_ASAP7_75t_R FILLER_125_359 ();
 DECAPx10_ASAP7_75t_R FILLER_125_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_417 ();
 DECAPx1_ASAP7_75t_R FILLER_125_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_451 ();
 FILLER_ASAP7_75t_R FILLER_125_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_462 ();
 FILLER_ASAP7_75t_R FILLER_125_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_471 ();
 FILLER_ASAP7_75t_R FILLER_125_480 ();
 DECAPx2_ASAP7_75t_R FILLER_125_488 ();
 DECAPx10_ASAP7_75t_R FILLER_125_501 ();
 DECAPx10_ASAP7_75t_R FILLER_125_523 ();
 DECAPx1_ASAP7_75t_R FILLER_125_545 ();
 DECAPx10_ASAP7_75t_R FILLER_125_552 ();
 DECAPx2_ASAP7_75t_R FILLER_125_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_580 ();
 FILLER_ASAP7_75t_R FILLER_125_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_604 ();
 FILLER_ASAP7_75t_R FILLER_125_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_628 ();
 DECAPx10_ASAP7_75t_R FILLER_125_635 ();
 DECAPx10_ASAP7_75t_R FILLER_125_657 ();
 DECAPx10_ASAP7_75t_R FILLER_125_679 ();
 DECAPx10_ASAP7_75t_R FILLER_125_701 ();
 DECAPx10_ASAP7_75t_R FILLER_125_723 ();
 DECAPx10_ASAP7_75t_R FILLER_125_745 ();
 DECAPx10_ASAP7_75t_R FILLER_125_767 ();
 DECAPx10_ASAP7_75t_R FILLER_125_789 ();
 DECAPx2_ASAP7_75t_R FILLER_125_811 ();
 FILLER_ASAP7_75t_R FILLER_125_817 ();
 DECAPx10_ASAP7_75t_R FILLER_125_829 ();
 FILLER_ASAP7_75t_R FILLER_125_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_853 ();
 DECAPx1_ASAP7_75t_R FILLER_125_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_864 ();
 DECAPx10_ASAP7_75t_R FILLER_125_886 ();
 FILLER_ASAP7_75t_R FILLER_125_908 ();
 DECAPx6_ASAP7_75t_R FILLER_125_926 ();
 FILLER_ASAP7_75t_R FILLER_125_940 ();
 DECAPx2_ASAP7_75t_R FILLER_125_948 ();
 FILLER_ASAP7_75t_R FILLER_125_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_956 ();
 DECAPx10_ASAP7_75t_R FILLER_125_965 ();
 FILLER_ASAP7_75t_R FILLER_125_987 ();
 DECAPx10_ASAP7_75t_R FILLER_125_995 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_126_2 ();
 DECAPx10_ASAP7_75t_R FILLER_126_24 ();
 DECAPx10_ASAP7_75t_R FILLER_126_46 ();
 DECAPx10_ASAP7_75t_R FILLER_126_68 ();
 DECAPx10_ASAP7_75t_R FILLER_126_90 ();
 DECAPx6_ASAP7_75t_R FILLER_126_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_126 ();
 DECAPx6_ASAP7_75t_R FILLER_126_137 ();
 DECAPx10_ASAP7_75t_R FILLER_126_167 ();
 DECAPx10_ASAP7_75t_R FILLER_126_189 ();
 DECAPx10_ASAP7_75t_R FILLER_126_211 ();
 DECAPx10_ASAP7_75t_R FILLER_126_233 ();
 DECAPx6_ASAP7_75t_R FILLER_126_255 ();
 DECAPx2_ASAP7_75t_R FILLER_126_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_275 ();
 DECAPx2_ASAP7_75t_R FILLER_126_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_288 ();
 DECAPx1_ASAP7_75t_R FILLER_126_299 ();
 DECAPx10_ASAP7_75t_R FILLER_126_313 ();
 DECAPx2_ASAP7_75t_R FILLER_126_335 ();
 FILLER_ASAP7_75t_R FILLER_126_341 ();
 DECAPx10_ASAP7_75t_R FILLER_126_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_415 ();
 DECAPx2_ASAP7_75t_R FILLER_126_432 ();
 FILLER_ASAP7_75t_R FILLER_126_438 ();
 DECAPx2_ASAP7_75t_R FILLER_126_454 ();
 FILLER_ASAP7_75t_R FILLER_126_460 ();
 DECAPx6_ASAP7_75t_R FILLER_126_464 ();
 DECAPx2_ASAP7_75t_R FILLER_126_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_484 ();
 DECAPx6_ASAP7_75t_R FILLER_126_494 ();
 DECAPx2_ASAP7_75t_R FILLER_126_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_547 ();
 DECAPx2_ASAP7_75t_R FILLER_126_572 ();
 FILLER_ASAP7_75t_R FILLER_126_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_595 ();
 DECAPx10_ASAP7_75t_R FILLER_126_599 ();
 DECAPx6_ASAP7_75t_R FILLER_126_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_635 ();
 DECAPx4_ASAP7_75t_R FILLER_126_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_655 ();
 DECAPx10_ASAP7_75t_R FILLER_126_662 ();
 DECAPx2_ASAP7_75t_R FILLER_126_684 ();
 DECAPx1_ASAP7_75t_R FILLER_126_697 ();
 FILLER_ASAP7_75t_R FILLER_126_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_719 ();
 DECAPx1_ASAP7_75t_R FILLER_126_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_730 ();
 DECAPx4_ASAP7_75t_R FILLER_126_748 ();
 FILLER_ASAP7_75t_R FILLER_126_758 ();
 DECAPx10_ASAP7_75t_R FILLER_126_763 ();
 DECAPx10_ASAP7_75t_R FILLER_126_785 ();
 DECAPx10_ASAP7_75t_R FILLER_126_807 ();
 DECAPx10_ASAP7_75t_R FILLER_126_829 ();
 DECAPx10_ASAP7_75t_R FILLER_126_851 ();
 DECAPx10_ASAP7_75t_R FILLER_126_873 ();
 DECAPx6_ASAP7_75t_R FILLER_126_895 ();
 DECAPx2_ASAP7_75t_R FILLER_126_952 ();
 FILLER_ASAP7_75t_R FILLER_126_964 ();
 DECAPx10_ASAP7_75t_R FILLER_126_972 ();
 DECAPx4_ASAP7_75t_R FILLER_126_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1095 ();
 FILLER_ASAP7_75t_R FILLER_126_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1134 ();
 FILLER_ASAP7_75t_R FILLER_126_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1158 ();
 FILLER_ASAP7_75t_R FILLER_126_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1189 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1280 ();
 FILLER_ASAP7_75t_R FILLER_126_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_127_2 ();
 DECAPx10_ASAP7_75t_R FILLER_127_24 ();
 DECAPx10_ASAP7_75t_R FILLER_127_46 ();
 DECAPx10_ASAP7_75t_R FILLER_127_68 ();
 DECAPx10_ASAP7_75t_R FILLER_127_90 ();
 DECAPx6_ASAP7_75t_R FILLER_127_112 ();
 FILLER_ASAP7_75t_R FILLER_127_126 ();
 DECAPx2_ASAP7_75t_R FILLER_127_142 ();
 FILLER_ASAP7_75t_R FILLER_127_148 ();
 DECAPx10_ASAP7_75t_R FILLER_127_176 ();
 DECAPx10_ASAP7_75t_R FILLER_127_198 ();
 DECAPx10_ASAP7_75t_R FILLER_127_220 ();
 DECAPx4_ASAP7_75t_R FILLER_127_242 ();
 DECAPx4_ASAP7_75t_R FILLER_127_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_272 ();
 DECAPx10_ASAP7_75t_R FILLER_127_283 ();
 DECAPx10_ASAP7_75t_R FILLER_127_305 ();
 DECAPx10_ASAP7_75t_R FILLER_127_327 ();
 FILLER_ASAP7_75t_R FILLER_127_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_351 ();
 DECAPx10_ASAP7_75t_R FILLER_127_368 ();
 DECAPx10_ASAP7_75t_R FILLER_127_390 ();
 DECAPx4_ASAP7_75t_R FILLER_127_412 ();
 DECAPx10_ASAP7_75t_R FILLER_127_428 ();
 DECAPx10_ASAP7_75t_R FILLER_127_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_472 ();
 DECAPx6_ASAP7_75t_R FILLER_127_480 ();
 FILLER_ASAP7_75t_R FILLER_127_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_496 ();
 DECAPx10_ASAP7_75t_R FILLER_127_505 ();
 DECAPx10_ASAP7_75t_R FILLER_127_527 ();
 FILLER_ASAP7_75t_R FILLER_127_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_560 ();
 DECAPx10_ASAP7_75t_R FILLER_127_591 ();
 DECAPx10_ASAP7_75t_R FILLER_127_613 ();
 DECAPx10_ASAP7_75t_R FILLER_127_635 ();
 DECAPx6_ASAP7_75t_R FILLER_127_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_671 ();
 FILLER_ASAP7_75t_R FILLER_127_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_680 ();
 DECAPx1_ASAP7_75t_R FILLER_127_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_699 ();
 DECAPx2_ASAP7_75t_R FILLER_127_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_726 ();
 DECAPx6_ASAP7_75t_R FILLER_127_734 ();
 DECAPx2_ASAP7_75t_R FILLER_127_748 ();
 DECAPx10_ASAP7_75t_R FILLER_127_775 ();
 FILLER_ASAP7_75t_R FILLER_127_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_799 ();
 DECAPx2_ASAP7_75t_R FILLER_127_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_827 ();
 DECAPx2_ASAP7_75t_R FILLER_127_837 ();
 DECAPx10_ASAP7_75t_R FILLER_127_849 ();
 FILLER_ASAP7_75t_R FILLER_127_871 ();
 DECAPx10_ASAP7_75t_R FILLER_127_876 ();
 DECAPx10_ASAP7_75t_R FILLER_127_898 ();
 DECAPx1_ASAP7_75t_R FILLER_127_920 ();
 DECAPx10_ASAP7_75t_R FILLER_127_950 ();
 DECAPx10_ASAP7_75t_R FILLER_127_972 ();
 DECAPx4_ASAP7_75t_R FILLER_127_994 ();
 FILLER_ASAP7_75t_R FILLER_127_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1012 ();
 FILLER_ASAP7_75t_R FILLER_127_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1052 ();
 FILLER_ASAP7_75t_R FILLER_127_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1092 ();
 FILLER_ASAP7_75t_R FILLER_127_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1172 ();
 FILLER_ASAP7_75t_R FILLER_127_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_128_2 ();
 DECAPx10_ASAP7_75t_R FILLER_128_24 ();
 DECAPx10_ASAP7_75t_R FILLER_128_46 ();
 DECAPx10_ASAP7_75t_R FILLER_128_68 ();
 DECAPx10_ASAP7_75t_R FILLER_128_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_112 ();
 DECAPx10_ASAP7_75t_R FILLER_128_121 ();
 DECAPx10_ASAP7_75t_R FILLER_128_143 ();
 DECAPx2_ASAP7_75t_R FILLER_128_171 ();
 FILLER_ASAP7_75t_R FILLER_128_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_179 ();
 DECAPx1_ASAP7_75t_R FILLER_128_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_197 ();
 DECAPx4_ASAP7_75t_R FILLER_128_208 ();
 FILLER_ASAP7_75t_R FILLER_128_218 ();
 FILLER_ASAP7_75t_R FILLER_128_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_232 ();
 DECAPx1_ASAP7_75t_R FILLER_128_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_253 ();
 FILLER_ASAP7_75t_R FILLER_128_264 ();
 FILLER_ASAP7_75t_R FILLER_128_288 ();
 DECAPx10_ASAP7_75t_R FILLER_128_303 ();
 DECAPx6_ASAP7_75t_R FILLER_128_325 ();
 DECAPx1_ASAP7_75t_R FILLER_128_339 ();
 DECAPx1_ASAP7_75t_R FILLER_128_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_373 ();
 DECAPx6_ASAP7_75t_R FILLER_128_390 ();
 DECAPx2_ASAP7_75t_R FILLER_128_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_410 ();
 FILLER_ASAP7_75t_R FILLER_128_425 ();
 DECAPx1_ASAP7_75t_R FILLER_128_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_439 ();
 DECAPx4_ASAP7_75t_R FILLER_128_452 ();
 DECAPx10_ASAP7_75t_R FILLER_128_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_516 ();
 DECAPx4_ASAP7_75t_R FILLER_128_548 ();
 FILLER_ASAP7_75t_R FILLER_128_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_560 ();
 FILLER_ASAP7_75t_R FILLER_128_577 ();
 DECAPx2_ASAP7_75t_R FILLER_128_586 ();
 FILLER_ASAP7_75t_R FILLER_128_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_594 ();
 DECAPx1_ASAP7_75t_R FILLER_128_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_628 ();
 FILLER_ASAP7_75t_R FILLER_128_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_634 ();
 DECAPx10_ASAP7_75t_R FILLER_128_684 ();
 DECAPx10_ASAP7_75t_R FILLER_128_706 ();
 DECAPx10_ASAP7_75t_R FILLER_128_728 ();
 DECAPx6_ASAP7_75t_R FILLER_128_750 ();
 DECAPx10_ASAP7_75t_R FILLER_128_773 ();
 DECAPx2_ASAP7_75t_R FILLER_128_795 ();
 FILLER_ASAP7_75t_R FILLER_128_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_813 ();
 FILLER_ASAP7_75t_R FILLER_128_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_819 ();
 DECAPx6_ASAP7_75t_R FILLER_128_826 ();
 DECAPx2_ASAP7_75t_R FILLER_128_840 ();
 DECAPx1_ASAP7_75t_R FILLER_128_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_867 ();
 DECAPx2_ASAP7_75t_R FILLER_128_876 ();
 FILLER_ASAP7_75t_R FILLER_128_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_884 ();
 DECAPx10_ASAP7_75t_R FILLER_128_893 ();
 DECAPx10_ASAP7_75t_R FILLER_128_915 ();
 DECAPx10_ASAP7_75t_R FILLER_128_937 ();
 DECAPx4_ASAP7_75t_R FILLER_128_959 ();
 DECAPx10_ASAP7_75t_R FILLER_128_977 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1005 ();
 FILLER_ASAP7_75t_R FILLER_128_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1263 ();
 FILLER_ASAP7_75t_R FILLER_128_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_129_2 ();
 DECAPx10_ASAP7_75t_R FILLER_129_24 ();
 DECAPx10_ASAP7_75t_R FILLER_129_46 ();
 DECAPx10_ASAP7_75t_R FILLER_129_68 ();
 DECAPx10_ASAP7_75t_R FILLER_129_90 ();
 DECAPx6_ASAP7_75t_R FILLER_129_112 ();
 DECAPx10_ASAP7_75t_R FILLER_129_140 ();
 DECAPx10_ASAP7_75t_R FILLER_129_162 ();
 DECAPx10_ASAP7_75t_R FILLER_129_184 ();
 DECAPx2_ASAP7_75t_R FILLER_129_206 ();
 DECAPx1_ASAP7_75t_R FILLER_129_226 ();
 DECAPx6_ASAP7_75t_R FILLER_129_236 ();
 DECAPx2_ASAP7_75t_R FILLER_129_250 ();
 DECAPx6_ASAP7_75t_R FILLER_129_273 ();
 DECAPx10_ASAP7_75t_R FILLER_129_309 ();
 DECAPx10_ASAP7_75t_R FILLER_129_331 ();
 DECAPx10_ASAP7_75t_R FILLER_129_369 ();
 DECAPx10_ASAP7_75t_R FILLER_129_391 ();
 DECAPx6_ASAP7_75t_R FILLER_129_413 ();
 DECAPx1_ASAP7_75t_R FILLER_129_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_431 ();
 DECAPx2_ASAP7_75t_R FILLER_129_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_478 ();
 DECAPx2_ASAP7_75t_R FILLER_129_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_505 ();
 DECAPx6_ASAP7_75t_R FILLER_129_531 ();
 DECAPx2_ASAP7_75t_R FILLER_129_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_551 ();
 DECAPx1_ASAP7_75t_R FILLER_129_555 ();
 FILLER_ASAP7_75t_R FILLER_129_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_606 ();
 FILLER_ASAP7_75t_R FILLER_129_629 ();
 DECAPx10_ASAP7_75t_R FILLER_129_645 ();
 DECAPx10_ASAP7_75t_R FILLER_129_667 ();
 DECAPx6_ASAP7_75t_R FILLER_129_689 ();
 FILLER_ASAP7_75t_R FILLER_129_703 ();
 DECAPx10_ASAP7_75t_R FILLER_129_711 ();
 DECAPx10_ASAP7_75t_R FILLER_129_733 ();
 DECAPx6_ASAP7_75t_R FILLER_129_755 ();
 DECAPx2_ASAP7_75t_R FILLER_129_778 ();
 DECAPx10_ASAP7_75t_R FILLER_129_813 ();
 DECAPx10_ASAP7_75t_R FILLER_129_835 ();
 DECAPx10_ASAP7_75t_R FILLER_129_857 ();
 DECAPx1_ASAP7_75t_R FILLER_129_879 ();
 DECAPx2_ASAP7_75t_R FILLER_129_893 ();
 FILLER_ASAP7_75t_R FILLER_129_899 ();
 DECAPx6_ASAP7_75t_R FILLER_129_910 ();
 DECAPx6_ASAP7_75t_R FILLER_129_926 ();
 DECAPx2_ASAP7_75t_R FILLER_129_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_946 ();
 DECAPx6_ASAP7_75t_R FILLER_129_961 ();
 DECAPx1_ASAP7_75t_R FILLER_129_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_985 ();
 DECAPx10_ASAP7_75t_R FILLER_129_994 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1016 ();
 FILLER_ASAP7_75t_R FILLER_129_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1040 ();
 FILLER_ASAP7_75t_R FILLER_129_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1056 ();
 FILLER_ASAP7_75t_R FILLER_129_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_129_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_129_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_129_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1179 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1206 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1241 ();
 FILLER_ASAP7_75t_R FILLER_129_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_130_2 ();
 DECAPx10_ASAP7_75t_R FILLER_130_24 ();
 DECAPx10_ASAP7_75t_R FILLER_130_46 ();
 DECAPx10_ASAP7_75t_R FILLER_130_68 ();
 DECAPx10_ASAP7_75t_R FILLER_130_90 ();
 DECAPx4_ASAP7_75t_R FILLER_130_112 ();
 DECAPx10_ASAP7_75t_R FILLER_130_128 ();
 DECAPx10_ASAP7_75t_R FILLER_130_150 ();
 DECAPx10_ASAP7_75t_R FILLER_130_172 ();
 DECAPx10_ASAP7_75t_R FILLER_130_194 ();
 DECAPx10_ASAP7_75t_R FILLER_130_216 ();
 DECAPx1_ASAP7_75t_R FILLER_130_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_242 ();
 DECAPx2_ASAP7_75t_R FILLER_130_257 ();
 FILLER_ASAP7_75t_R FILLER_130_263 ();
 FILLER_ASAP7_75t_R FILLER_130_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_285 ();
 DECAPx10_ASAP7_75t_R FILLER_130_307 ();
 DECAPx10_ASAP7_75t_R FILLER_130_329 ();
 DECAPx1_ASAP7_75t_R FILLER_130_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_401 ();
 DECAPx2_ASAP7_75t_R FILLER_130_410 ();
 DECAPx10_ASAP7_75t_R FILLER_130_431 ();
 FILLER_ASAP7_75t_R FILLER_130_453 ();
 FILLER_ASAP7_75t_R FILLER_130_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_466 ();
 DECAPx4_ASAP7_75t_R FILLER_130_473 ();
 FILLER_ASAP7_75t_R FILLER_130_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_485 ();
 DECAPx10_ASAP7_75t_R FILLER_130_499 ();
 DECAPx1_ASAP7_75t_R FILLER_130_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_525 ();
 FILLER_ASAP7_75t_R FILLER_130_557 ();
 FILLER_ASAP7_75t_R FILLER_130_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_569 ();
 DECAPx1_ASAP7_75t_R FILLER_130_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_577 ();
 DECAPx10_ASAP7_75t_R FILLER_130_593 ();
 DECAPx2_ASAP7_75t_R FILLER_130_615 ();
 DECAPx1_ASAP7_75t_R FILLER_130_629 ();
 DECAPx10_ASAP7_75t_R FILLER_130_641 ();
 DECAPx6_ASAP7_75t_R FILLER_130_663 ();
 DECAPx2_ASAP7_75t_R FILLER_130_677 ();
 DECAPx2_ASAP7_75t_R FILLER_130_695 ();
 FILLER_ASAP7_75t_R FILLER_130_701 ();
 DECAPx6_ASAP7_75t_R FILLER_130_715 ();
 DECAPx1_ASAP7_75t_R FILLER_130_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_733 ();
 DECAPx10_ASAP7_75t_R FILLER_130_756 ();
 DECAPx10_ASAP7_75t_R FILLER_130_778 ();
 DECAPx10_ASAP7_75t_R FILLER_130_800 ();
 DECAPx10_ASAP7_75t_R FILLER_130_822 ();
 DECAPx10_ASAP7_75t_R FILLER_130_844 ();
 DECAPx10_ASAP7_75t_R FILLER_130_866 ();
 DECAPx10_ASAP7_75t_R FILLER_130_888 ();
 DECAPx10_ASAP7_75t_R FILLER_130_910 ();
 DECAPx6_ASAP7_75t_R FILLER_130_932 ();
 DECAPx1_ASAP7_75t_R FILLER_130_946 ();
 DECAPx4_ASAP7_75t_R FILLER_130_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_974 ();
 DECAPx10_ASAP7_75t_R FILLER_130_981 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1003 ();
 FILLER_ASAP7_75t_R FILLER_130_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1022 ();
 FILLER_ASAP7_75t_R FILLER_130_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_131_2 ();
 DECAPx10_ASAP7_75t_R FILLER_131_24 ();
 DECAPx10_ASAP7_75t_R FILLER_131_46 ();
 DECAPx10_ASAP7_75t_R FILLER_131_68 ();
 DECAPx10_ASAP7_75t_R FILLER_131_90 ();
 DECAPx10_ASAP7_75t_R FILLER_131_112 ();
 DECAPx4_ASAP7_75t_R FILLER_131_134 ();
 FILLER_ASAP7_75t_R FILLER_131_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_146 ();
 DECAPx1_ASAP7_75t_R FILLER_131_153 ();
 DECAPx10_ASAP7_75t_R FILLER_131_171 ();
 DECAPx10_ASAP7_75t_R FILLER_131_193 ();
 DECAPx10_ASAP7_75t_R FILLER_131_223 ();
 DECAPx10_ASAP7_75t_R FILLER_131_245 ();
 DECAPx10_ASAP7_75t_R FILLER_131_267 ();
 DECAPx2_ASAP7_75t_R FILLER_131_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_312 ();
 DECAPx10_ASAP7_75t_R FILLER_131_321 ();
 DECAPx2_ASAP7_75t_R FILLER_131_343 ();
 FILLER_ASAP7_75t_R FILLER_131_349 ();
 DECAPx10_ASAP7_75t_R FILLER_131_367 ();
 DECAPx6_ASAP7_75t_R FILLER_131_389 ();
 DECAPx1_ASAP7_75t_R FILLER_131_403 ();
 DECAPx2_ASAP7_75t_R FILLER_131_410 ();
 DECAPx10_ASAP7_75t_R FILLER_131_425 ();
 DECAPx1_ASAP7_75t_R FILLER_131_447 ();
 DECAPx10_ASAP7_75t_R FILLER_131_459 ();
 DECAPx10_ASAP7_75t_R FILLER_131_481 ();
 DECAPx4_ASAP7_75t_R FILLER_131_503 ();
 DECAPx1_ASAP7_75t_R FILLER_131_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_541 ();
 DECAPx1_ASAP7_75t_R FILLER_131_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_554 ();
 DECAPx10_ASAP7_75t_R FILLER_131_561 ();
 DECAPx4_ASAP7_75t_R FILLER_131_583 ();
 FILLER_ASAP7_75t_R FILLER_131_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_595 ();
 DECAPx10_ASAP7_75t_R FILLER_131_602 ();
 DECAPx2_ASAP7_75t_R FILLER_131_624 ();
 FILLER_ASAP7_75t_R FILLER_131_630 ();
 DECAPx10_ASAP7_75t_R FILLER_131_652 ();
 FILLER_ASAP7_75t_R FILLER_131_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_676 ();
 FILLER_ASAP7_75t_R FILLER_131_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_691 ();
 DECAPx2_ASAP7_75t_R FILLER_131_698 ();
 DECAPx10_ASAP7_75t_R FILLER_131_728 ();
 DECAPx1_ASAP7_75t_R FILLER_131_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_754 ();
 DECAPx10_ASAP7_75t_R FILLER_131_761 ();
 DECAPx10_ASAP7_75t_R FILLER_131_783 ();
 DECAPx10_ASAP7_75t_R FILLER_131_805 ();
 DECAPx10_ASAP7_75t_R FILLER_131_827 ();
 DECAPx10_ASAP7_75t_R FILLER_131_849 ();
 DECAPx10_ASAP7_75t_R FILLER_131_871 ();
 FILLER_ASAP7_75t_R FILLER_131_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_895 ();
 DECAPx6_ASAP7_75t_R FILLER_131_910 ();
 DECAPx10_ASAP7_75t_R FILLER_131_926 ();
 DECAPx2_ASAP7_75t_R FILLER_131_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_954 ();
 DECAPx10_ASAP7_75t_R FILLER_131_979 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1087 ();
 FILLER_ASAP7_75t_R FILLER_131_1109 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1121 ();
 FILLER_ASAP7_75t_R FILLER_131_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1208 ();
 FILLER_ASAP7_75t_R FILLER_131_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_132_2 ();
 DECAPx10_ASAP7_75t_R FILLER_132_24 ();
 DECAPx10_ASAP7_75t_R FILLER_132_46 ();
 DECAPx10_ASAP7_75t_R FILLER_132_68 ();
 DECAPx10_ASAP7_75t_R FILLER_132_90 ();
 DECAPx2_ASAP7_75t_R FILLER_132_112 ();
 FILLER_ASAP7_75t_R FILLER_132_118 ();
 DECAPx10_ASAP7_75t_R FILLER_132_126 ();
 DECAPx10_ASAP7_75t_R FILLER_132_148 ();
 DECAPx10_ASAP7_75t_R FILLER_132_170 ();
 DECAPx10_ASAP7_75t_R FILLER_132_192 ();
 DECAPx10_ASAP7_75t_R FILLER_132_214 ();
 DECAPx10_ASAP7_75t_R FILLER_132_236 ();
 DECAPx2_ASAP7_75t_R FILLER_132_268 ();
 FILLER_ASAP7_75t_R FILLER_132_274 ();
 DECAPx4_ASAP7_75t_R FILLER_132_283 ();
 FILLER_ASAP7_75t_R FILLER_132_300 ();
 FILLER_ASAP7_75t_R FILLER_132_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_310 ();
 DECAPx2_ASAP7_75t_R FILLER_132_336 ();
 FILLER_ASAP7_75t_R FILLER_132_342 ();
 DECAPx10_ASAP7_75t_R FILLER_132_360 ();
 DECAPx10_ASAP7_75t_R FILLER_132_382 ();
 DECAPx6_ASAP7_75t_R FILLER_132_404 ();
 FILLER_ASAP7_75t_R FILLER_132_418 ();
 DECAPx6_ASAP7_75t_R FILLER_132_429 ();
 FILLER_ASAP7_75t_R FILLER_132_443 ();
 FILLER_ASAP7_75t_R FILLER_132_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_461 ();
 DECAPx10_ASAP7_75t_R FILLER_132_464 ();
 DECAPx10_ASAP7_75t_R FILLER_132_486 ();
 DECAPx1_ASAP7_75t_R FILLER_132_508 ();
 DECAPx4_ASAP7_75t_R FILLER_132_527 ();
 FILLER_ASAP7_75t_R FILLER_132_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_539 ();
 DECAPx10_ASAP7_75t_R FILLER_132_546 ();
 DECAPx10_ASAP7_75t_R FILLER_132_568 ();
 DECAPx1_ASAP7_75t_R FILLER_132_590 ();
 DECAPx4_ASAP7_75t_R FILLER_132_618 ();
 FILLER_ASAP7_75t_R FILLER_132_628 ();
 DECAPx4_ASAP7_75t_R FILLER_132_638 ();
 DECAPx10_ASAP7_75t_R FILLER_132_664 ();
 DECAPx10_ASAP7_75t_R FILLER_132_686 ();
 DECAPx4_ASAP7_75t_R FILLER_132_708 ();
 FILLER_ASAP7_75t_R FILLER_132_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_720 ();
 DECAPx4_ASAP7_75t_R FILLER_132_732 ();
 FILLER_ASAP7_75t_R FILLER_132_742 ();
 DECAPx10_ASAP7_75t_R FILLER_132_750 ();
 DECAPx6_ASAP7_75t_R FILLER_132_772 ();
 DECAPx1_ASAP7_75t_R FILLER_132_786 ();
 DECAPx10_ASAP7_75t_R FILLER_132_812 ();
 DECAPx10_ASAP7_75t_R FILLER_132_834 ();
 FILLER_ASAP7_75t_R FILLER_132_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_858 ();
 DECAPx10_ASAP7_75t_R FILLER_132_865 ();
 DECAPx10_ASAP7_75t_R FILLER_132_887 ();
 DECAPx6_ASAP7_75t_R FILLER_132_909 ();
 DECAPx2_ASAP7_75t_R FILLER_132_923 ();
 DECAPx2_ASAP7_75t_R FILLER_132_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_945 ();
 DECAPx10_ASAP7_75t_R FILLER_132_978 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1066 ();
 FILLER_ASAP7_75t_R FILLER_132_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1141 ();
 FILLER_ASAP7_75t_R FILLER_132_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1181 ();
 FILLER_ASAP7_75t_R FILLER_132_1195 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1206 ();
 FILLER_ASAP7_75t_R FILLER_132_1220 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_133_2 ();
 DECAPx10_ASAP7_75t_R FILLER_133_24 ();
 DECAPx10_ASAP7_75t_R FILLER_133_46 ();
 DECAPx10_ASAP7_75t_R FILLER_133_68 ();
 DECAPx10_ASAP7_75t_R FILLER_133_90 ();
 DECAPx1_ASAP7_75t_R FILLER_133_130 ();
 DECAPx10_ASAP7_75t_R FILLER_133_142 ();
 FILLER_ASAP7_75t_R FILLER_133_164 ();
 FILLER_ASAP7_75t_R FILLER_133_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_182 ();
 DECAPx6_ASAP7_75t_R FILLER_133_202 ();
 DECAPx2_ASAP7_75t_R FILLER_133_216 ();
 DECAPx2_ASAP7_75t_R FILLER_133_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_254 ();
 DECAPx10_ASAP7_75t_R FILLER_133_263 ();
 FILLER_ASAP7_75t_R FILLER_133_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_287 ();
 DECAPx10_ASAP7_75t_R FILLER_133_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_336 ();
 DECAPx1_ASAP7_75t_R FILLER_133_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_351 ();
 DECAPx10_ASAP7_75t_R FILLER_133_368 ();
 DECAPx2_ASAP7_75t_R FILLER_133_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_396 ();
 DECAPx2_ASAP7_75t_R FILLER_133_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_418 ();
 DECAPx2_ASAP7_75t_R FILLER_133_425 ();
 FILLER_ASAP7_75t_R FILLER_133_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_433 ();
 FILLER_ASAP7_75t_R FILLER_133_450 ();
 DECAPx6_ASAP7_75t_R FILLER_133_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_498 ();
 DECAPx10_ASAP7_75t_R FILLER_133_520 ();
 FILLER_ASAP7_75t_R FILLER_133_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_552 ();
 DECAPx1_ASAP7_75t_R FILLER_133_556 ();
 DECAPx6_ASAP7_75t_R FILLER_133_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_598 ();
 DECAPx10_ASAP7_75t_R FILLER_133_607 ();
 DECAPx6_ASAP7_75t_R FILLER_133_629 ();
 DECAPx10_ASAP7_75t_R FILLER_133_683 ();
 DECAPx10_ASAP7_75t_R FILLER_133_705 ();
 DECAPx10_ASAP7_75t_R FILLER_133_727 ();
 DECAPx10_ASAP7_75t_R FILLER_133_749 ();
 DECAPx10_ASAP7_75t_R FILLER_133_771 ();
 DECAPx10_ASAP7_75t_R FILLER_133_793 ();
 DECAPx1_ASAP7_75t_R FILLER_133_815 ();
 DECAPx4_ASAP7_75t_R FILLER_133_831 ();
 FILLER_ASAP7_75t_R FILLER_133_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_843 ();
 DECAPx10_ASAP7_75t_R FILLER_133_858 ();
 DECAPx10_ASAP7_75t_R FILLER_133_880 ();
 DECAPx10_ASAP7_75t_R FILLER_133_902 ();
 DECAPx2_ASAP7_75t_R FILLER_133_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_932 ();
 DECAPx10_ASAP7_75t_R FILLER_133_951 ();
 DECAPx10_ASAP7_75t_R FILLER_133_973 ();
 DECAPx2_ASAP7_75t_R FILLER_133_995 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1092 ();
 FILLER_ASAP7_75t_R FILLER_133_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1186 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_134_2 ();
 DECAPx10_ASAP7_75t_R FILLER_134_24 ();
 DECAPx10_ASAP7_75t_R FILLER_134_46 ();
 DECAPx10_ASAP7_75t_R FILLER_134_68 ();
 DECAPx10_ASAP7_75t_R FILLER_134_90 ();
 DECAPx10_ASAP7_75t_R FILLER_134_112 ();
 DECAPx1_ASAP7_75t_R FILLER_134_134 ();
 DECAPx6_ASAP7_75t_R FILLER_134_144 ();
 FILLER_ASAP7_75t_R FILLER_134_158 ();
 DECAPx10_ASAP7_75t_R FILLER_134_166 ();
 DECAPx2_ASAP7_75t_R FILLER_134_188 ();
 FILLER_ASAP7_75t_R FILLER_134_194 ();
 FILLER_ASAP7_75t_R FILLER_134_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_205 ();
 DECAPx2_ASAP7_75t_R FILLER_134_216 ();
 DECAPx4_ASAP7_75t_R FILLER_134_230 ();
 FILLER_ASAP7_75t_R FILLER_134_240 ();
 DECAPx6_ASAP7_75t_R FILLER_134_252 ();
 DECAPx2_ASAP7_75t_R FILLER_134_266 ();
 DECAPx6_ASAP7_75t_R FILLER_134_282 ();
 FILLER_ASAP7_75t_R FILLER_134_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_298 ();
 DECAPx6_ASAP7_75t_R FILLER_134_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_319 ();
 DECAPx10_ASAP7_75t_R FILLER_134_329 ();
 DECAPx6_ASAP7_75t_R FILLER_134_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_365 ();
 DECAPx6_ASAP7_75t_R FILLER_134_374 ();
 FILLER_ASAP7_75t_R FILLER_134_388 ();
 FILLER_ASAP7_75t_R FILLER_134_403 ();
 DECAPx2_ASAP7_75t_R FILLER_134_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_425 ();
 DECAPx1_ASAP7_75t_R FILLER_134_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_436 ();
 FILLER_ASAP7_75t_R FILLER_134_447 ();
 DECAPx1_ASAP7_75t_R FILLER_134_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_461 ();
 DECAPx4_ASAP7_75t_R FILLER_134_472 ();
 FILLER_ASAP7_75t_R FILLER_134_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_484 ();
 DECAPx10_ASAP7_75t_R FILLER_134_494 ();
 DECAPx2_ASAP7_75t_R FILLER_134_516 ();
 FILLER_ASAP7_75t_R FILLER_134_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_524 ();
 FILLER_ASAP7_75t_R FILLER_134_533 ();
 FILLER_ASAP7_75t_R FILLER_134_556 ();
 DECAPx2_ASAP7_75t_R FILLER_134_573 ();
 DECAPx6_ASAP7_75t_R FILLER_134_600 ();
 DECAPx6_ASAP7_75t_R FILLER_134_620 ();
 FILLER_ASAP7_75t_R FILLER_134_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_636 ();
 DECAPx4_ASAP7_75t_R FILLER_134_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_653 ();
 DECAPx10_ASAP7_75t_R FILLER_134_662 ();
 DECAPx6_ASAP7_75t_R FILLER_134_684 ();
 DECAPx10_ASAP7_75t_R FILLER_134_710 ();
 DECAPx10_ASAP7_75t_R FILLER_134_732 ();
 DECAPx4_ASAP7_75t_R FILLER_134_754 ();
 FILLER_ASAP7_75t_R FILLER_134_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_766 ();
 DECAPx4_ASAP7_75t_R FILLER_134_779 ();
 DECAPx10_ASAP7_75t_R FILLER_134_797 ();
 DECAPx10_ASAP7_75t_R FILLER_134_819 ();
 DECAPx10_ASAP7_75t_R FILLER_134_841 ();
 DECAPx10_ASAP7_75t_R FILLER_134_863 ();
 FILLER_ASAP7_75t_R FILLER_134_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_887 ();
 DECAPx6_ASAP7_75t_R FILLER_134_904 ();
 DECAPx1_ASAP7_75t_R FILLER_134_918 ();
 DECAPx6_ASAP7_75t_R FILLER_134_936 ();
 DECAPx2_ASAP7_75t_R FILLER_134_950 ();
 DECAPx10_ASAP7_75t_R FILLER_134_966 ();
 DECAPx10_ASAP7_75t_R FILLER_134_988 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1054 ();
 FILLER_ASAP7_75t_R FILLER_134_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1127 ();
 FILLER_ASAP7_75t_R FILLER_134_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1157 ();
 FILLER_ASAP7_75t_R FILLER_134_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1208 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1230 ();
 FILLER_ASAP7_75t_R FILLER_134_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1269 ();
 FILLER_ASAP7_75t_R FILLER_134_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_135_2 ();
 DECAPx10_ASAP7_75t_R FILLER_135_24 ();
 DECAPx10_ASAP7_75t_R FILLER_135_46 ();
 DECAPx10_ASAP7_75t_R FILLER_135_68 ();
 DECAPx10_ASAP7_75t_R FILLER_135_90 ();
 DECAPx10_ASAP7_75t_R FILLER_135_112 ();
 FILLER_ASAP7_75t_R FILLER_135_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_136 ();
 DECAPx6_ASAP7_75t_R FILLER_135_159 ();
 DECAPx1_ASAP7_75t_R FILLER_135_173 ();
 DECAPx10_ASAP7_75t_R FILLER_135_183 ();
 DECAPx6_ASAP7_75t_R FILLER_135_205 ();
 DECAPx1_ASAP7_75t_R FILLER_135_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_223 ();
 DECAPx2_ASAP7_75t_R FILLER_135_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_236 ();
 DECAPx10_ASAP7_75t_R FILLER_135_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_288 ();
 DECAPx2_ASAP7_75t_R FILLER_135_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_302 ();
 DECAPx4_ASAP7_75t_R FILLER_135_311 ();
 DECAPx2_ASAP7_75t_R FILLER_135_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_333 ();
 DECAPx10_ASAP7_75t_R FILLER_135_344 ();
 DECAPx4_ASAP7_75t_R FILLER_135_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_376 ();
 FILLER_ASAP7_75t_R FILLER_135_383 ();
 DECAPx4_ASAP7_75t_R FILLER_135_421 ();
 DECAPx4_ASAP7_75t_R FILLER_135_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_449 ();
 FILLER_ASAP7_75t_R FILLER_135_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_461 ();
 FILLER_ASAP7_75t_R FILLER_135_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_472 ();
 DECAPx10_ASAP7_75t_R FILLER_135_483 ();
 DECAPx2_ASAP7_75t_R FILLER_135_505 ();
 FILLER_ASAP7_75t_R FILLER_135_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_513 ();
 FILLER_ASAP7_75t_R FILLER_135_538 ();
 DECAPx10_ASAP7_75t_R FILLER_135_546 ();
 DECAPx10_ASAP7_75t_R FILLER_135_568 ();
 DECAPx1_ASAP7_75t_R FILLER_135_590 ();
 DECAPx10_ASAP7_75t_R FILLER_135_597 ();
 DECAPx10_ASAP7_75t_R FILLER_135_619 ();
 DECAPx6_ASAP7_75t_R FILLER_135_641 ();
 DECAPx1_ASAP7_75t_R FILLER_135_655 ();
 DECAPx10_ASAP7_75t_R FILLER_135_665 ();
 DECAPx4_ASAP7_75t_R FILLER_135_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_704 ();
 DECAPx6_ASAP7_75t_R FILLER_135_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_725 ();
 DECAPx10_ASAP7_75t_R FILLER_135_738 ();
 DECAPx10_ASAP7_75t_R FILLER_135_760 ();
 DECAPx6_ASAP7_75t_R FILLER_135_782 ();
 FILLER_ASAP7_75t_R FILLER_135_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_798 ();
 DECAPx10_ASAP7_75t_R FILLER_135_817 ();
 DECAPx10_ASAP7_75t_R FILLER_135_839 ();
 DECAPx10_ASAP7_75t_R FILLER_135_861 ();
 DECAPx10_ASAP7_75t_R FILLER_135_883 ();
 DECAPx6_ASAP7_75t_R FILLER_135_905 ();
 DECAPx1_ASAP7_75t_R FILLER_135_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_923 ();
 DECAPx10_ASAP7_75t_R FILLER_135_926 ();
 DECAPx2_ASAP7_75t_R FILLER_135_948 ();
 FILLER_ASAP7_75t_R FILLER_135_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_956 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1001 ();
 FILLER_ASAP7_75t_R FILLER_135_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1067 ();
 FILLER_ASAP7_75t_R FILLER_135_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1123 ();
 FILLER_ASAP7_75t_R FILLER_135_1133 ();
 FILLER_ASAP7_75t_R FILLER_135_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1152 ();
 FILLER_ASAP7_75t_R FILLER_135_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1241 ();
 FILLER_ASAP7_75t_R FILLER_135_1247 ();
 FILLER_ASAP7_75t_R FILLER_135_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1259 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_136_2 ();
 DECAPx10_ASAP7_75t_R FILLER_136_24 ();
 DECAPx10_ASAP7_75t_R FILLER_136_46 ();
 DECAPx10_ASAP7_75t_R FILLER_136_68 ();
 DECAPx10_ASAP7_75t_R FILLER_136_90 ();
 DECAPx10_ASAP7_75t_R FILLER_136_112 ();
 DECAPx6_ASAP7_75t_R FILLER_136_134 ();
 FILLER_ASAP7_75t_R FILLER_136_148 ();
 DECAPx10_ASAP7_75t_R FILLER_136_156 ();
 DECAPx10_ASAP7_75t_R FILLER_136_178 ();
 DECAPx6_ASAP7_75t_R FILLER_136_200 ();
 DECAPx2_ASAP7_75t_R FILLER_136_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_220 ();
 DECAPx10_ASAP7_75t_R FILLER_136_227 ();
 DECAPx2_ASAP7_75t_R FILLER_136_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_255 ();
 DECAPx2_ASAP7_75t_R FILLER_136_266 ();
 FILLER_ASAP7_75t_R FILLER_136_272 ();
 DECAPx10_ASAP7_75t_R FILLER_136_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_302 ();
 DECAPx2_ASAP7_75t_R FILLER_136_310 ();
 FILLER_ASAP7_75t_R FILLER_136_316 ();
 DECAPx2_ASAP7_75t_R FILLER_136_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_336 ();
 DECAPx6_ASAP7_75t_R FILLER_136_347 ();
 DECAPx2_ASAP7_75t_R FILLER_136_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_367 ();
 FILLER_ASAP7_75t_R FILLER_136_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_394 ();
 DECAPx10_ASAP7_75t_R FILLER_136_415 ();
 DECAPx6_ASAP7_75t_R FILLER_136_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_451 ();
 FILLER_ASAP7_75t_R FILLER_136_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_466 ();
 DECAPx1_ASAP7_75t_R FILLER_136_475 ();
 DECAPx6_ASAP7_75t_R FILLER_136_495 ();
 DECAPx2_ASAP7_75t_R FILLER_136_509 ();
 FILLER_ASAP7_75t_R FILLER_136_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_531 ();
 DECAPx10_ASAP7_75t_R FILLER_136_536 ();
 DECAPx10_ASAP7_75t_R FILLER_136_558 ();
 FILLER_ASAP7_75t_R FILLER_136_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_582 ();
 FILLER_ASAP7_75t_R FILLER_136_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_599 ();
 DECAPx2_ASAP7_75t_R FILLER_136_614 ();
 DECAPx6_ASAP7_75t_R FILLER_136_623 ();
 DECAPx1_ASAP7_75t_R FILLER_136_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_641 ();
 DECAPx2_ASAP7_75t_R FILLER_136_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_670 ();
 DECAPx4_ASAP7_75t_R FILLER_136_678 ();
 DECAPx10_ASAP7_75t_R FILLER_136_698 ();
 DECAPx10_ASAP7_75t_R FILLER_136_720 ();
 FILLER_ASAP7_75t_R FILLER_136_742 ();
 DECAPx10_ASAP7_75t_R FILLER_136_754 ();
 DECAPx10_ASAP7_75t_R FILLER_136_776 ();
 DECAPx10_ASAP7_75t_R FILLER_136_798 ();
 DECAPx10_ASAP7_75t_R FILLER_136_820 ();
 DECAPx10_ASAP7_75t_R FILLER_136_842 ();
 DECAPx10_ASAP7_75t_R FILLER_136_864 ();
 DECAPx10_ASAP7_75t_R FILLER_136_886 ();
 DECAPx10_ASAP7_75t_R FILLER_136_908 ();
 DECAPx10_ASAP7_75t_R FILLER_136_950 ();
 DECAPx6_ASAP7_75t_R FILLER_136_972 ();
 FILLER_ASAP7_75t_R FILLER_136_986 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1012 ();
 FILLER_ASAP7_75t_R FILLER_136_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1034 ();
 FILLER_ASAP7_75t_R FILLER_136_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1071 ();
 FILLER_ASAP7_75t_R FILLER_136_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1102 ();
 FILLER_ASAP7_75t_R FILLER_136_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1231 ();
 FILLER_ASAP7_75t_R FILLER_136_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_137_2 ();
 DECAPx10_ASAP7_75t_R FILLER_137_24 ();
 DECAPx10_ASAP7_75t_R FILLER_137_46 ();
 DECAPx10_ASAP7_75t_R FILLER_137_68 ();
 DECAPx4_ASAP7_75t_R FILLER_137_90 ();
 FILLER_ASAP7_75t_R FILLER_137_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_102 ();
 DECAPx2_ASAP7_75t_R FILLER_137_127 ();
 FILLER_ASAP7_75t_R FILLER_137_133 ();
 DECAPx10_ASAP7_75t_R FILLER_137_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_165 ();
 DECAPx10_ASAP7_75t_R FILLER_137_178 ();
 DECAPx2_ASAP7_75t_R FILLER_137_200 ();
 DECAPx10_ASAP7_75t_R FILLER_137_216 ();
 DECAPx1_ASAP7_75t_R FILLER_137_238 ();
 DECAPx10_ASAP7_75t_R FILLER_137_247 ();
 DECAPx6_ASAP7_75t_R FILLER_137_269 ();
 DECAPx1_ASAP7_75t_R FILLER_137_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_287 ();
 DECAPx10_ASAP7_75t_R FILLER_137_294 ();
 DECAPx6_ASAP7_75t_R FILLER_137_328 ();
 DECAPx10_ASAP7_75t_R FILLER_137_348 ();
 DECAPx10_ASAP7_75t_R FILLER_137_377 ();
 DECAPx4_ASAP7_75t_R FILLER_137_399 ();
 FILLER_ASAP7_75t_R FILLER_137_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_451 ();
 DECAPx10_ASAP7_75t_R FILLER_137_462 ();
 DECAPx4_ASAP7_75t_R FILLER_137_484 ();
 FILLER_ASAP7_75t_R FILLER_137_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_496 ();
 DECAPx2_ASAP7_75t_R FILLER_137_505 ();
 FILLER_ASAP7_75t_R FILLER_137_511 ();
 DECAPx10_ASAP7_75t_R FILLER_137_519 ();
 FILLER_ASAP7_75t_R FILLER_137_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_552 ();
 DECAPx2_ASAP7_75t_R FILLER_137_556 ();
 FILLER_ASAP7_75t_R FILLER_137_562 ();
 FILLER_ASAP7_75t_R FILLER_137_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_574 ();
 DECAPx2_ASAP7_75t_R FILLER_137_578 ();
 FILLER_ASAP7_75t_R FILLER_137_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_586 ();
 DECAPx2_ASAP7_75t_R FILLER_137_595 ();
 FILLER_ASAP7_75t_R FILLER_137_601 ();
 DECAPx10_ASAP7_75t_R FILLER_137_624 ();
 DECAPx1_ASAP7_75t_R FILLER_137_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_650 ();
 DECAPx4_ASAP7_75t_R FILLER_137_661 ();
 FILLER_ASAP7_75t_R FILLER_137_671 ();
 FILLER_ASAP7_75t_R FILLER_137_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_685 ();
 DECAPx1_ASAP7_75t_R FILLER_137_698 ();
 DECAPx6_ASAP7_75t_R FILLER_137_708 ();
 FILLER_ASAP7_75t_R FILLER_137_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_724 ();
 FILLER_ASAP7_75t_R FILLER_137_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_733 ();
 FILLER_ASAP7_75t_R FILLER_137_740 ();
 DECAPx10_ASAP7_75t_R FILLER_137_750 ();
 DECAPx10_ASAP7_75t_R FILLER_137_772 ();
 DECAPx10_ASAP7_75t_R FILLER_137_794 ();
 DECAPx10_ASAP7_75t_R FILLER_137_816 ();
 DECAPx10_ASAP7_75t_R FILLER_137_838 ();
 DECAPx2_ASAP7_75t_R FILLER_137_860 ();
 FILLER_ASAP7_75t_R FILLER_137_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_868 ();
 DECAPx10_ASAP7_75t_R FILLER_137_875 ();
 DECAPx10_ASAP7_75t_R FILLER_137_897 ();
 DECAPx1_ASAP7_75t_R FILLER_137_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_923 ();
 DECAPx4_ASAP7_75t_R FILLER_137_942 ();
 FILLER_ASAP7_75t_R FILLER_137_952 ();
 DECAPx10_ASAP7_75t_R FILLER_137_978 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1050 ();
 FILLER_ASAP7_75t_R FILLER_137_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1073 ();
 FILLER_ASAP7_75t_R FILLER_137_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1195 ();
 FILLER_ASAP7_75t_R FILLER_137_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1280 ();
 FILLER_ASAP7_75t_R FILLER_137_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_138_2 ();
 DECAPx10_ASAP7_75t_R FILLER_138_24 ();
 DECAPx10_ASAP7_75t_R FILLER_138_46 ();
 DECAPx10_ASAP7_75t_R FILLER_138_68 ();
 DECAPx10_ASAP7_75t_R FILLER_138_90 ();
 DECAPx6_ASAP7_75t_R FILLER_138_112 ();
 FILLER_ASAP7_75t_R FILLER_138_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_148 ();
 DECAPx10_ASAP7_75t_R FILLER_138_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_196 ();
 DECAPx10_ASAP7_75t_R FILLER_138_219 ();
 DECAPx1_ASAP7_75t_R FILLER_138_241 ();
 DECAPx2_ASAP7_75t_R FILLER_138_254 ();
 DECAPx1_ASAP7_75t_R FILLER_138_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_280 ();
 DECAPx2_ASAP7_75t_R FILLER_138_291 ();
 FILLER_ASAP7_75t_R FILLER_138_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_299 ();
 DECAPx1_ASAP7_75t_R FILLER_138_316 ();
 DECAPx1_ASAP7_75t_R FILLER_138_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_338 ();
 DECAPx10_ASAP7_75t_R FILLER_138_347 ();
 DECAPx10_ASAP7_75t_R FILLER_138_369 ();
 DECAPx2_ASAP7_75t_R FILLER_138_391 ();
 DECAPx2_ASAP7_75t_R FILLER_138_401 ();
 FILLER_ASAP7_75t_R FILLER_138_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_409 ();
 DECAPx2_ASAP7_75t_R FILLER_138_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_422 ();
 DECAPx4_ASAP7_75t_R FILLER_138_433 ();
 FILLER_ASAP7_75t_R FILLER_138_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_445 ();
 DECAPx2_ASAP7_75t_R FILLER_138_453 ();
 FILLER_ASAP7_75t_R FILLER_138_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_461 ();
 DECAPx2_ASAP7_75t_R FILLER_138_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_470 ();
 DECAPx4_ASAP7_75t_R FILLER_138_527 ();
 DECAPx1_ASAP7_75t_R FILLER_138_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_583 ();
 DECAPx1_ASAP7_75t_R FILLER_138_590 ();
 DECAPx10_ASAP7_75t_R FILLER_138_597 ();
 DECAPx10_ASAP7_75t_R FILLER_138_619 ();
 FILLER_ASAP7_75t_R FILLER_138_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_643 ();
 DECAPx10_ASAP7_75t_R FILLER_138_652 ();
 DECAPx10_ASAP7_75t_R FILLER_138_674 ();
 FILLER_ASAP7_75t_R FILLER_138_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_707 ();
 DECAPx10_ASAP7_75t_R FILLER_138_720 ();
 DECAPx10_ASAP7_75t_R FILLER_138_742 ();
 DECAPx10_ASAP7_75t_R FILLER_138_764 ();
 DECAPx10_ASAP7_75t_R FILLER_138_786 ();
 DECAPx6_ASAP7_75t_R FILLER_138_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_822 ();
 DECAPx10_ASAP7_75t_R FILLER_138_829 ();
 DECAPx4_ASAP7_75t_R FILLER_138_851 ();
 DECAPx10_ASAP7_75t_R FILLER_138_869 ();
 DECAPx6_ASAP7_75t_R FILLER_138_891 ();
 FILLER_ASAP7_75t_R FILLER_138_905 ();
 DECAPx10_ASAP7_75t_R FILLER_138_935 ();
 DECAPx10_ASAP7_75t_R FILLER_138_957 ();
 DECAPx10_ASAP7_75t_R FILLER_138_979 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1146 ();
 FILLER_ASAP7_75t_R FILLER_138_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1161 ();
 FILLER_ASAP7_75t_R FILLER_138_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_139_2 ();
 DECAPx10_ASAP7_75t_R FILLER_139_24 ();
 DECAPx10_ASAP7_75t_R FILLER_139_46 ();
 DECAPx10_ASAP7_75t_R FILLER_139_68 ();
 DECAPx10_ASAP7_75t_R FILLER_139_90 ();
 FILLER_ASAP7_75t_R FILLER_139_112 ();
 DECAPx10_ASAP7_75t_R FILLER_139_122 ();
 DECAPx10_ASAP7_75t_R FILLER_139_144 ();
 FILLER_ASAP7_75t_R FILLER_139_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_168 ();
 DECAPx1_ASAP7_75t_R FILLER_139_179 ();
 DECAPx2_ASAP7_75t_R FILLER_139_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_200 ();
 DECAPx2_ASAP7_75t_R FILLER_139_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_217 ();
 DECAPx6_ASAP7_75t_R FILLER_139_221 ();
 FILLER_ASAP7_75t_R FILLER_139_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_237 ();
 DECAPx1_ASAP7_75t_R FILLER_139_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_251 ();
 DECAPx4_ASAP7_75t_R FILLER_139_264 ();
 FILLER_ASAP7_75t_R FILLER_139_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_276 ();
 DECAPx6_ASAP7_75t_R FILLER_139_285 ();
 DECAPx2_ASAP7_75t_R FILLER_139_299 ();
 DECAPx4_ASAP7_75t_R FILLER_139_345 ();
 FILLER_ASAP7_75t_R FILLER_139_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_357 ();
 FILLER_ASAP7_75t_R FILLER_139_377 ();
 DECAPx2_ASAP7_75t_R FILLER_139_385 ();
 FILLER_ASAP7_75t_R FILLER_139_391 ();
 DECAPx2_ASAP7_75t_R FILLER_139_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_406 ();
 DECAPx6_ASAP7_75t_R FILLER_139_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_429 ();
 DECAPx10_ASAP7_75t_R FILLER_139_440 ();
 FILLER_ASAP7_75t_R FILLER_139_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_464 ();
 DECAPx10_ASAP7_75t_R FILLER_139_491 ();
 DECAPx4_ASAP7_75t_R FILLER_139_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_523 ();
 FILLER_ASAP7_75t_R FILLER_139_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_534 ();
 FILLER_ASAP7_75t_R FILLER_139_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_540 ();
 DECAPx4_ASAP7_75t_R FILLER_139_547 ();
 FILLER_ASAP7_75t_R FILLER_139_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_559 ();
 DECAPx6_ASAP7_75t_R FILLER_139_566 ();
 FILLER_ASAP7_75t_R FILLER_139_580 ();
 DECAPx10_ASAP7_75t_R FILLER_139_603 ();
 FILLER_ASAP7_75t_R FILLER_139_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_627 ();
 DECAPx4_ASAP7_75t_R FILLER_139_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_666 ();
 DECAPx4_ASAP7_75t_R FILLER_139_681 ();
 FILLER_ASAP7_75t_R FILLER_139_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_715 ();
 DECAPx10_ASAP7_75t_R FILLER_139_722 ();
 DECAPx10_ASAP7_75t_R FILLER_139_744 ();
 DECAPx2_ASAP7_75t_R FILLER_139_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_772 ();
 DECAPx6_ASAP7_75t_R FILLER_139_781 ();
 DECAPx1_ASAP7_75t_R FILLER_139_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_799 ();
 DECAPx10_ASAP7_75t_R FILLER_139_806 ();
 DECAPx10_ASAP7_75t_R FILLER_139_828 ();
 DECAPx10_ASAP7_75t_R FILLER_139_850 ();
 DECAPx10_ASAP7_75t_R FILLER_139_872 ();
 DECAPx10_ASAP7_75t_R FILLER_139_894 ();
 DECAPx2_ASAP7_75t_R FILLER_139_916 ();
 FILLER_ASAP7_75t_R FILLER_139_922 ();
 DECAPx4_ASAP7_75t_R FILLER_139_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_936 ();
 DECAPx10_ASAP7_75t_R FILLER_139_973 ();
 FILLER_ASAP7_75t_R FILLER_139_995 ();
 FILLER_ASAP7_75t_R FILLER_139_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1017 ();
 FILLER_ASAP7_75t_R FILLER_139_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1125 ();
 FILLER_ASAP7_75t_R FILLER_139_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1244 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1251 ();
 FILLER_ASAP7_75t_R FILLER_139_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_140_2 ();
 DECAPx10_ASAP7_75t_R FILLER_140_24 ();
 DECAPx10_ASAP7_75t_R FILLER_140_46 ();
 DECAPx10_ASAP7_75t_R FILLER_140_68 ();
 DECAPx10_ASAP7_75t_R FILLER_140_90 ();
 DECAPx10_ASAP7_75t_R FILLER_140_112 ();
 DECAPx10_ASAP7_75t_R FILLER_140_134 ();
 DECAPx6_ASAP7_75t_R FILLER_140_156 ();
 DECAPx2_ASAP7_75t_R FILLER_140_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_176 ();
 DECAPx10_ASAP7_75t_R FILLER_140_203 ();
 DECAPx2_ASAP7_75t_R FILLER_140_225 ();
 DECAPx1_ASAP7_75t_R FILLER_140_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_247 ();
 DECAPx2_ASAP7_75t_R FILLER_140_258 ();
 FILLER_ASAP7_75t_R FILLER_140_264 ();
 DECAPx2_ASAP7_75t_R FILLER_140_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_278 ();
 DECAPx2_ASAP7_75t_R FILLER_140_282 ();
 FILLER_ASAP7_75t_R FILLER_140_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_296 ();
 DECAPx6_ASAP7_75t_R FILLER_140_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_328 ();
 DECAPx4_ASAP7_75t_R FILLER_140_343 ();
 DECAPx6_ASAP7_75t_R FILLER_140_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_377 ();
 DECAPx2_ASAP7_75t_R FILLER_140_412 ();
 FILLER_ASAP7_75t_R FILLER_140_418 ();
 DECAPx10_ASAP7_75t_R FILLER_140_430 ();
 DECAPx4_ASAP7_75t_R FILLER_140_452 ();
 DECAPx6_ASAP7_75t_R FILLER_140_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_478 ();
 DECAPx10_ASAP7_75t_R FILLER_140_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_516 ();
 DECAPx10_ASAP7_75t_R FILLER_140_538 ();
 DECAPx10_ASAP7_75t_R FILLER_140_560 ();
 DECAPx6_ASAP7_75t_R FILLER_140_582 ();
 DECAPx2_ASAP7_75t_R FILLER_140_596 ();
 DECAPx4_ASAP7_75t_R FILLER_140_623 ();
 DECAPx10_ASAP7_75t_R FILLER_140_636 ();
 DECAPx10_ASAP7_75t_R FILLER_140_658 ();
 DECAPx6_ASAP7_75t_R FILLER_140_680 ();
 FILLER_ASAP7_75t_R FILLER_140_694 ();
 DECAPx2_ASAP7_75t_R FILLER_140_702 ();
 DECAPx10_ASAP7_75t_R FILLER_140_714 ();
 DECAPx10_ASAP7_75t_R FILLER_140_736 ();
 DECAPx10_ASAP7_75t_R FILLER_140_758 ();
 DECAPx10_ASAP7_75t_R FILLER_140_780 ();
 DECAPx4_ASAP7_75t_R FILLER_140_802 ();
 DECAPx10_ASAP7_75t_R FILLER_140_818 ();
 DECAPx10_ASAP7_75t_R FILLER_140_840 ();
 DECAPx10_ASAP7_75t_R FILLER_140_862 ();
 DECAPx10_ASAP7_75t_R FILLER_140_884 ();
 DECAPx10_ASAP7_75t_R FILLER_140_906 ();
 DECAPx10_ASAP7_75t_R FILLER_140_928 ();
 DECAPx10_ASAP7_75t_R FILLER_140_950 ();
 DECAPx10_ASAP7_75t_R FILLER_140_982 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1102 ();
 FILLER_ASAP7_75t_R FILLER_140_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1145 ();
 FILLER_ASAP7_75t_R FILLER_140_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1159 ();
 FILLER_ASAP7_75t_R FILLER_140_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1226 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_141_2 ();
 DECAPx10_ASAP7_75t_R FILLER_141_24 ();
 DECAPx10_ASAP7_75t_R FILLER_141_46 ();
 DECAPx10_ASAP7_75t_R FILLER_141_68 ();
 DECAPx10_ASAP7_75t_R FILLER_141_90 ();
 DECAPx10_ASAP7_75t_R FILLER_141_112 ();
 DECAPx10_ASAP7_75t_R FILLER_141_134 ();
 DECAPx6_ASAP7_75t_R FILLER_141_156 ();
 DECAPx10_ASAP7_75t_R FILLER_141_173 ();
 DECAPx4_ASAP7_75t_R FILLER_141_195 ();
 FILLER_ASAP7_75t_R FILLER_141_205 ();
 DECAPx10_ASAP7_75t_R FILLER_141_233 ();
 DECAPx4_ASAP7_75t_R FILLER_141_255 ();
 FILLER_ASAP7_75t_R FILLER_141_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_303 ();
 DECAPx10_ASAP7_75t_R FILLER_141_320 ();
 DECAPx10_ASAP7_75t_R FILLER_141_342 ();
 DECAPx2_ASAP7_75t_R FILLER_141_364 ();
 DECAPx4_ASAP7_75t_R FILLER_141_384 ();
 DECAPx1_ASAP7_75t_R FILLER_141_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_416 ();
 DECAPx1_ASAP7_75t_R FILLER_141_425 ();
 FILLER_ASAP7_75t_R FILLER_141_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_441 ();
 DECAPx10_ASAP7_75t_R FILLER_141_448 ();
 DECAPx1_ASAP7_75t_R FILLER_141_470 ();
 DECAPx10_ASAP7_75t_R FILLER_141_484 ();
 DECAPx6_ASAP7_75t_R FILLER_141_506 ();
 FILLER_ASAP7_75t_R FILLER_141_520 ();
 DECAPx1_ASAP7_75t_R FILLER_141_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_532 ();
 DECAPx6_ASAP7_75t_R FILLER_141_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_568 ();
 DECAPx4_ASAP7_75t_R FILLER_141_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_599 ();
 DECAPx10_ASAP7_75t_R FILLER_141_614 ();
 DECAPx4_ASAP7_75t_R FILLER_141_636 ();
 FILLER_ASAP7_75t_R FILLER_141_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_648 ();
 DECAPx1_ASAP7_75t_R FILLER_141_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_663 ();
 DECAPx1_ASAP7_75t_R FILLER_141_670 ();
 DECAPx4_ASAP7_75t_R FILLER_141_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_718 ();
 DECAPx2_ASAP7_75t_R FILLER_141_726 ();
 FILLER_ASAP7_75t_R FILLER_141_732 ();
 DECAPx10_ASAP7_75t_R FILLER_141_744 ();
 DECAPx10_ASAP7_75t_R FILLER_141_766 ();
 DECAPx10_ASAP7_75t_R FILLER_141_788 ();
 DECAPx10_ASAP7_75t_R FILLER_141_810 ();
 DECAPx4_ASAP7_75t_R FILLER_141_832 ();
 FILLER_ASAP7_75t_R FILLER_141_842 ();
 DECAPx6_ASAP7_75t_R FILLER_141_850 ();
 DECAPx1_ASAP7_75t_R FILLER_141_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_868 ();
 DECAPx10_ASAP7_75t_R FILLER_141_875 ();
 DECAPx10_ASAP7_75t_R FILLER_141_897 ();
 DECAPx1_ASAP7_75t_R FILLER_141_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_923 ();
 DECAPx10_ASAP7_75t_R FILLER_141_926 ();
 DECAPx1_ASAP7_75t_R FILLER_141_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_952 ();
 DECAPx6_ASAP7_75t_R FILLER_141_959 ();
 DECAPx2_ASAP7_75t_R FILLER_141_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_979 ();
 DECAPx10_ASAP7_75t_R FILLER_141_994 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1038 ();
 FILLER_ASAP7_75t_R FILLER_141_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1193 ();
 FILLER_ASAP7_75t_R FILLER_141_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1205 ();
 FILLER_ASAP7_75t_R FILLER_141_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1220 ();
 FILLER_ASAP7_75t_R FILLER_141_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1244 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1251 ();
 FILLER_ASAP7_75t_R FILLER_141_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_142_2 ();
 DECAPx10_ASAP7_75t_R FILLER_142_24 ();
 DECAPx10_ASAP7_75t_R FILLER_142_46 ();
 DECAPx10_ASAP7_75t_R FILLER_142_68 ();
 FILLER_ASAP7_75t_R FILLER_142_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_92 ();
 FILLER_ASAP7_75t_R FILLER_142_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_121 ();
 FILLER_ASAP7_75t_R FILLER_142_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_130 ();
 DECAPx6_ASAP7_75t_R FILLER_142_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_157 ();
 DECAPx4_ASAP7_75t_R FILLER_142_191 ();
 FILLER_ASAP7_75t_R FILLER_142_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_215 ();
 DECAPx10_ASAP7_75t_R FILLER_142_223 ();
 FILLER_ASAP7_75t_R FILLER_142_245 ();
 DECAPx6_ASAP7_75t_R FILLER_142_255 ();
 DECAPx1_ASAP7_75t_R FILLER_142_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_273 ();
 DECAPx4_ASAP7_75t_R FILLER_142_319 ();
 FILLER_ASAP7_75t_R FILLER_142_329 ();
 DECAPx10_ASAP7_75t_R FILLER_142_337 ();
 DECAPx4_ASAP7_75t_R FILLER_142_359 ();
 FILLER_ASAP7_75t_R FILLER_142_369 ();
 DECAPx6_ASAP7_75t_R FILLER_142_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_394 ();
 DECAPx6_ASAP7_75t_R FILLER_142_408 ();
 DECAPx2_ASAP7_75t_R FILLER_142_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_428 ();
 DECAPx2_ASAP7_75t_R FILLER_142_456 ();
 DECAPx10_ASAP7_75t_R FILLER_142_474 ();
 DECAPx6_ASAP7_75t_R FILLER_142_496 ();
 DECAPx10_ASAP7_75t_R FILLER_142_516 ();
 FILLER_ASAP7_75t_R FILLER_142_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_584 ();
 DECAPx4_ASAP7_75t_R FILLER_142_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_616 ();
 DECAPx4_ASAP7_75t_R FILLER_142_628 ();
 DECAPx6_ASAP7_75t_R FILLER_142_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_662 ();
 FILLER_ASAP7_75t_R FILLER_142_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_671 ();
 DECAPx10_ASAP7_75t_R FILLER_142_680 ();
 DECAPx10_ASAP7_75t_R FILLER_142_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_724 ();
 DECAPx10_ASAP7_75t_R FILLER_142_737 ();
 DECAPx10_ASAP7_75t_R FILLER_142_759 ();
 DECAPx10_ASAP7_75t_R FILLER_142_781 ();
 DECAPx4_ASAP7_75t_R FILLER_142_803 ();
 DECAPx1_ASAP7_75t_R FILLER_142_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_829 ();
 DECAPx10_ASAP7_75t_R FILLER_142_840 ();
 DECAPx10_ASAP7_75t_R FILLER_142_862 ();
 DECAPx6_ASAP7_75t_R FILLER_142_884 ();
 FILLER_ASAP7_75t_R FILLER_142_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_900 ();
 DECAPx6_ASAP7_75t_R FILLER_142_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_922 ();
 DECAPx10_ASAP7_75t_R FILLER_142_935 ();
 DECAPx1_ASAP7_75t_R FILLER_142_967 ();
 DECAPx2_ASAP7_75t_R FILLER_142_987 ();
 FILLER_ASAP7_75t_R FILLER_142_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_995 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1022 ();
 FILLER_ASAP7_75t_R FILLER_142_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1052 ();
 FILLER_ASAP7_75t_R FILLER_142_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1136 ();
 FILLER_ASAP7_75t_R FILLER_142_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1201 ();
 FILLER_ASAP7_75t_R FILLER_142_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1225 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1238 ();
 FILLER_ASAP7_75t_R FILLER_142_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_143_2 ();
 DECAPx10_ASAP7_75t_R FILLER_143_24 ();
 DECAPx10_ASAP7_75t_R FILLER_143_46 ();
 DECAPx4_ASAP7_75t_R FILLER_143_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_78 ();
 DECAPx4_ASAP7_75t_R FILLER_143_105 ();
 FILLER_ASAP7_75t_R FILLER_143_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_117 ();
 FILLER_ASAP7_75t_R FILLER_143_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_137 ();
 DECAPx1_ASAP7_75t_R FILLER_143_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_189 ();
 DECAPx2_ASAP7_75t_R FILLER_143_210 ();
 DECAPx2_ASAP7_75t_R FILLER_143_232 ();
 FILLER_ASAP7_75t_R FILLER_143_238 ();
 DECAPx10_ASAP7_75t_R FILLER_143_248 ();
 DECAPx6_ASAP7_75t_R FILLER_143_270 ();
 DECAPx2_ASAP7_75t_R FILLER_143_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_290 ();
 DECAPx10_ASAP7_75t_R FILLER_143_301 ();
 DECAPx6_ASAP7_75t_R FILLER_143_323 ();
 FILLER_ASAP7_75t_R FILLER_143_337 ();
 DECAPx2_ASAP7_75t_R FILLER_143_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_351 ();
 DECAPx10_ASAP7_75t_R FILLER_143_355 ();
 FILLER_ASAP7_75t_R FILLER_143_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_379 ();
 DECAPx10_ASAP7_75t_R FILLER_143_392 ();
 DECAPx4_ASAP7_75t_R FILLER_143_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_424 ();
 DECAPx6_ASAP7_75t_R FILLER_143_435 ();
 DECAPx2_ASAP7_75t_R FILLER_143_449 ();
 FILLER_ASAP7_75t_R FILLER_143_461 ();
 DECAPx2_ASAP7_75t_R FILLER_143_485 ();
 FILLER_ASAP7_75t_R FILLER_143_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_493 ();
 DECAPx4_ASAP7_75t_R FILLER_143_526 ();
 FILLER_ASAP7_75t_R FILLER_143_536 ();
 DECAPx2_ASAP7_75t_R FILLER_143_544 ();
 FILLER_ASAP7_75t_R FILLER_143_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_552 ();
 DECAPx4_ASAP7_75t_R FILLER_143_570 ();
 FILLER_ASAP7_75t_R FILLER_143_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_582 ();
 DECAPx2_ASAP7_75t_R FILLER_143_606 ();
 FILLER_ASAP7_75t_R FILLER_143_612 ();
 DECAPx4_ASAP7_75t_R FILLER_143_635 ();
 FILLER_ASAP7_75t_R FILLER_143_645 ();
 DECAPx2_ASAP7_75t_R FILLER_143_669 ();
 FILLER_ASAP7_75t_R FILLER_143_675 ();
 DECAPx4_ASAP7_75t_R FILLER_143_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_693 ();
 FILLER_ASAP7_75t_R FILLER_143_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_708 ();
 DECAPx10_ASAP7_75t_R FILLER_143_719 ();
 DECAPx4_ASAP7_75t_R FILLER_143_741 ();
 FILLER_ASAP7_75t_R FILLER_143_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_753 ();
 DECAPx10_ASAP7_75t_R FILLER_143_776 ();
 DECAPx10_ASAP7_75t_R FILLER_143_798 ();
 DECAPx10_ASAP7_75t_R FILLER_143_820 ();
 DECAPx10_ASAP7_75t_R FILLER_143_842 ();
 DECAPx10_ASAP7_75t_R FILLER_143_864 ();
 DECAPx10_ASAP7_75t_R FILLER_143_886 ();
 DECAPx6_ASAP7_75t_R FILLER_143_908 ();
 FILLER_ASAP7_75t_R FILLER_143_922 ();
 DECAPx4_ASAP7_75t_R FILLER_143_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_936 ();
 DECAPx6_ASAP7_75t_R FILLER_143_945 ();
 DECAPx6_ASAP7_75t_R FILLER_143_965 ();
 FILLER_ASAP7_75t_R FILLER_143_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_981 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1170 ();
 FILLER_ASAP7_75t_R FILLER_143_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1210 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_144_2 ();
 DECAPx10_ASAP7_75t_R FILLER_144_24 ();
 DECAPx10_ASAP7_75t_R FILLER_144_46 ();
 DECAPx10_ASAP7_75t_R FILLER_144_68 ();
 DECAPx1_ASAP7_75t_R FILLER_144_90 ();
 DECAPx2_ASAP7_75t_R FILLER_144_97 ();
 FILLER_ASAP7_75t_R FILLER_144_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_105 ();
 DECAPx2_ASAP7_75t_R FILLER_144_109 ();
 FILLER_ASAP7_75t_R FILLER_144_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_126 ();
 FILLER_ASAP7_75t_R FILLER_144_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_185 ();
 DECAPx2_ASAP7_75t_R FILLER_144_192 ();
 FILLER_ASAP7_75t_R FILLER_144_198 ();
 DECAPx2_ASAP7_75t_R FILLER_144_206 ();
 DECAPx4_ASAP7_75t_R FILLER_144_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_235 ();
 DECAPx1_ASAP7_75t_R FILLER_144_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_247 ();
 DECAPx6_ASAP7_75t_R FILLER_144_251 ();
 DECAPx10_ASAP7_75t_R FILLER_144_282 ();
 DECAPx6_ASAP7_75t_R FILLER_144_304 ();
 DECAPx1_ASAP7_75t_R FILLER_144_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_322 ();
 DECAPx6_ASAP7_75t_R FILLER_144_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_377 ();
 FILLER_ASAP7_75t_R FILLER_144_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_385 ();
 DECAPx4_ASAP7_75t_R FILLER_144_402 ();
 FILLER_ASAP7_75t_R FILLER_144_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_414 ();
 DECAPx4_ASAP7_75t_R FILLER_144_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_435 ();
 DECAPx2_ASAP7_75t_R FILLER_144_442 ();
 FILLER_ASAP7_75t_R FILLER_144_448 ();
 FILLER_ASAP7_75t_R FILLER_144_460 ();
 DECAPx1_ASAP7_75t_R FILLER_144_464 ();
 DECAPx4_ASAP7_75t_R FILLER_144_479 ();
 DECAPx4_ASAP7_75t_R FILLER_144_503 ();
 FILLER_ASAP7_75t_R FILLER_144_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_515 ();
 DECAPx1_ASAP7_75t_R FILLER_144_527 ();
 DECAPx10_ASAP7_75t_R FILLER_144_555 ();
 DECAPx10_ASAP7_75t_R FILLER_144_577 ();
 DECAPx10_ASAP7_75t_R FILLER_144_599 ();
 DECAPx10_ASAP7_75t_R FILLER_144_621 ();
 DECAPx10_ASAP7_75t_R FILLER_144_643 ();
 DECAPx1_ASAP7_75t_R FILLER_144_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_679 ();
 DECAPx10_ASAP7_75t_R FILLER_144_687 ();
 DECAPx2_ASAP7_75t_R FILLER_144_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_715 ();
 DECAPx10_ASAP7_75t_R FILLER_144_723 ();
 DECAPx10_ASAP7_75t_R FILLER_144_745 ();
 DECAPx2_ASAP7_75t_R FILLER_144_767 ();
 FILLER_ASAP7_75t_R FILLER_144_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_775 ();
 DECAPx10_ASAP7_75t_R FILLER_144_782 ();
 DECAPx10_ASAP7_75t_R FILLER_144_804 ();
 DECAPx10_ASAP7_75t_R FILLER_144_826 ();
 DECAPx10_ASAP7_75t_R FILLER_144_848 ();
 DECAPx10_ASAP7_75t_R FILLER_144_870 ();
 DECAPx10_ASAP7_75t_R FILLER_144_898 ();
 DECAPx10_ASAP7_75t_R FILLER_144_920 ();
 DECAPx6_ASAP7_75t_R FILLER_144_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_956 ();
 FILLER_ASAP7_75t_R FILLER_144_967 ();
 DECAPx10_ASAP7_75t_R FILLER_144_978 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1022 ();
 FILLER_ASAP7_75t_R FILLER_144_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1165 ();
 FILLER_ASAP7_75t_R FILLER_144_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1198 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1227 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1234 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_145_2 ();
 DECAPx10_ASAP7_75t_R FILLER_145_24 ();
 DECAPx10_ASAP7_75t_R FILLER_145_46 ();
 DECAPx10_ASAP7_75t_R FILLER_145_68 ();
 DECAPx6_ASAP7_75t_R FILLER_145_90 ();
 DECAPx1_ASAP7_75t_R FILLER_145_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_108 ();
 DECAPx6_ASAP7_75t_R FILLER_145_112 ();
 DECAPx2_ASAP7_75t_R FILLER_145_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_145 ();
 DECAPx2_ASAP7_75t_R FILLER_145_154 ();
 DECAPx10_ASAP7_75t_R FILLER_145_178 ();
 DECAPx6_ASAP7_75t_R FILLER_145_200 ();
 FILLER_ASAP7_75t_R FILLER_145_214 ();
 FILLER_ASAP7_75t_R FILLER_145_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_226 ();
 DECAPx10_ASAP7_75t_R FILLER_145_260 ();
 DECAPx2_ASAP7_75t_R FILLER_145_282 ();
 FILLER_ASAP7_75t_R FILLER_145_288 ();
 FILLER_ASAP7_75t_R FILLER_145_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_298 ();
 DECAPx10_ASAP7_75t_R FILLER_145_305 ();
 DECAPx6_ASAP7_75t_R FILLER_145_339 ();
 DECAPx2_ASAP7_75t_R FILLER_145_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_359 ();
 DECAPx10_ASAP7_75t_R FILLER_145_363 ();
 DECAPx2_ASAP7_75t_R FILLER_145_385 ();
 FILLER_ASAP7_75t_R FILLER_145_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_393 ();
 DECAPx6_ASAP7_75t_R FILLER_145_400 ();
 FILLER_ASAP7_75t_R FILLER_145_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_434 ();
 DECAPx6_ASAP7_75t_R FILLER_145_445 ();
 DECAPx1_ASAP7_75t_R FILLER_145_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_463 ();
 DECAPx4_ASAP7_75t_R FILLER_145_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_485 ();
 FILLER_ASAP7_75t_R FILLER_145_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_508 ();
 DECAPx4_ASAP7_75t_R FILLER_145_530 ();
 FILLER_ASAP7_75t_R FILLER_145_540 ();
 DECAPx2_ASAP7_75t_R FILLER_145_550 ();
 FILLER_ASAP7_75t_R FILLER_145_556 ();
 DECAPx1_ASAP7_75t_R FILLER_145_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_583 ();
 DECAPx10_ASAP7_75t_R FILLER_145_611 ();
 DECAPx6_ASAP7_75t_R FILLER_145_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_653 ();
 DECAPx6_ASAP7_75t_R FILLER_145_660 ();
 DECAPx1_ASAP7_75t_R FILLER_145_674 ();
 DECAPx1_ASAP7_75t_R FILLER_145_685 ();
 DECAPx4_ASAP7_75t_R FILLER_145_705 ();
 FILLER_ASAP7_75t_R FILLER_145_715 ();
 DECAPx10_ASAP7_75t_R FILLER_145_726 ();
 DECAPx10_ASAP7_75t_R FILLER_145_748 ();
 DECAPx10_ASAP7_75t_R FILLER_145_770 ();
 FILLER_ASAP7_75t_R FILLER_145_792 ();
 DECAPx6_ASAP7_75t_R FILLER_145_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_814 ();
 DECAPx10_ASAP7_75t_R FILLER_145_821 ();
 DECAPx10_ASAP7_75t_R FILLER_145_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_865 ();
 DECAPx10_ASAP7_75t_R FILLER_145_876 ();
 DECAPx10_ASAP7_75t_R FILLER_145_898 ();
 DECAPx1_ASAP7_75t_R FILLER_145_920 ();
 DECAPx1_ASAP7_75t_R FILLER_145_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_930 ();
 DECAPx10_ASAP7_75t_R FILLER_145_945 ();
 DECAPx1_ASAP7_75t_R FILLER_145_967 ();
 DECAPx10_ASAP7_75t_R FILLER_145_979 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1132 ();
 FILLER_ASAP7_75t_R FILLER_145_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1191 ();
 FILLER_ASAP7_75t_R FILLER_145_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1213 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1240 ();
 FILLER_ASAP7_75t_R FILLER_145_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1280 ();
 FILLER_ASAP7_75t_R FILLER_145_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_146_2 ();
 DECAPx10_ASAP7_75t_R FILLER_146_24 ();
 DECAPx10_ASAP7_75t_R FILLER_146_46 ();
 DECAPx10_ASAP7_75t_R FILLER_146_68 ();
 DECAPx2_ASAP7_75t_R FILLER_146_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_96 ();
 DECAPx2_ASAP7_75t_R FILLER_146_123 ();
 FILLER_ASAP7_75t_R FILLER_146_129 ();
 DECAPx1_ASAP7_75t_R FILLER_146_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_152 ();
 DECAPx2_ASAP7_75t_R FILLER_146_163 ();
 DECAPx10_ASAP7_75t_R FILLER_146_177 ();
 DECAPx6_ASAP7_75t_R FILLER_146_199 ();
 DECAPx2_ASAP7_75t_R FILLER_146_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_219 ();
 DECAPx2_ASAP7_75t_R FILLER_146_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_238 ();
 DECAPx6_ASAP7_75t_R FILLER_146_245 ();
 DECAPx1_ASAP7_75t_R FILLER_146_259 ();
 FILLER_ASAP7_75t_R FILLER_146_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_281 ();
 DECAPx2_ASAP7_75t_R FILLER_146_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_315 ();
 DECAPx1_ASAP7_75t_R FILLER_146_326 ();
 DECAPx2_ASAP7_75t_R FILLER_146_337 ();
 FILLER_ASAP7_75t_R FILLER_146_343 ();
 DECAPx1_ASAP7_75t_R FILLER_146_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_375 ();
 DECAPx4_ASAP7_75t_R FILLER_146_386 ();
 DECAPx6_ASAP7_75t_R FILLER_146_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_426 ();
 DECAPx6_ASAP7_75t_R FILLER_146_442 ();
 DECAPx2_ASAP7_75t_R FILLER_146_456 ();
 DECAPx2_ASAP7_75t_R FILLER_146_464 ();
 DECAPx6_ASAP7_75t_R FILLER_146_496 ();
 FILLER_ASAP7_75t_R FILLER_146_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_512 ();
 DECAPx6_ASAP7_75t_R FILLER_146_519 ();
 DECAPx1_ASAP7_75t_R FILLER_146_533 ();
 DECAPx4_ASAP7_75t_R FILLER_146_543 ();
 FILLER_ASAP7_75t_R FILLER_146_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_555 ();
 DECAPx4_ASAP7_75t_R FILLER_146_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_580 ();
 DECAPx2_ASAP7_75t_R FILLER_146_603 ();
 FILLER_ASAP7_75t_R FILLER_146_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_611 ();
 DECAPx10_ASAP7_75t_R FILLER_146_627 ();
 DECAPx10_ASAP7_75t_R FILLER_146_649 ();
 DECAPx10_ASAP7_75t_R FILLER_146_671 ();
 DECAPx2_ASAP7_75t_R FILLER_146_693 ();
 DECAPx10_ASAP7_75t_R FILLER_146_705 ();
 DECAPx1_ASAP7_75t_R FILLER_146_727 ();
 DECAPx10_ASAP7_75t_R FILLER_146_739 ();
 DECAPx1_ASAP7_75t_R FILLER_146_761 ();
 DECAPx10_ASAP7_75t_R FILLER_146_781 ();
 DECAPx10_ASAP7_75t_R FILLER_146_803 ();
 DECAPx6_ASAP7_75t_R FILLER_146_825 ();
 FILLER_ASAP7_75t_R FILLER_146_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_841 ();
 DECAPx6_ASAP7_75t_R FILLER_146_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_864 ();
 DECAPx10_ASAP7_75t_R FILLER_146_871 ();
 DECAPx10_ASAP7_75t_R FILLER_146_893 ();
 DECAPx10_ASAP7_75t_R FILLER_146_915 ();
 DECAPx10_ASAP7_75t_R FILLER_146_937 ();
 DECAPx10_ASAP7_75t_R FILLER_146_959 ();
 FILLER_ASAP7_75t_R FILLER_146_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_983 ();
 DECAPx10_ASAP7_75t_R FILLER_146_998 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1042 ();
 FILLER_ASAP7_75t_R FILLER_146_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1071 ();
 FILLER_ASAP7_75t_R FILLER_146_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_147_2 ();
 DECAPx10_ASAP7_75t_R FILLER_147_24 ();
 DECAPx10_ASAP7_75t_R FILLER_147_46 ();
 DECAPx10_ASAP7_75t_R FILLER_147_68 ();
 DECAPx10_ASAP7_75t_R FILLER_147_90 ();
 DECAPx6_ASAP7_75t_R FILLER_147_112 ();
 DECAPx2_ASAP7_75t_R FILLER_147_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_132 ();
 DECAPx10_ASAP7_75t_R FILLER_147_139 ();
 DECAPx4_ASAP7_75t_R FILLER_147_161 ();
 FILLER_ASAP7_75t_R FILLER_147_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_173 ();
 DECAPx10_ASAP7_75t_R FILLER_147_194 ();
 FILLER_ASAP7_75t_R FILLER_147_216 ();
 DECAPx2_ASAP7_75t_R FILLER_147_223 ();
 DECAPx4_ASAP7_75t_R FILLER_147_236 ();
 FILLER_ASAP7_75t_R FILLER_147_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_248 ();
 FILLER_ASAP7_75t_R FILLER_147_275 ();
 DECAPx10_ASAP7_75t_R FILLER_147_290 ();
 DECAPx6_ASAP7_75t_R FILLER_147_312 ();
 FILLER_ASAP7_75t_R FILLER_147_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_328 ();
 DECAPx10_ASAP7_75t_R FILLER_147_333 ();
 DECAPx10_ASAP7_75t_R FILLER_147_355 ();
 DECAPx4_ASAP7_75t_R FILLER_147_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_387 ();
 DECAPx10_ASAP7_75t_R FILLER_147_398 ();
 DECAPx2_ASAP7_75t_R FILLER_147_420 ();
 DECAPx10_ASAP7_75t_R FILLER_147_434 ();
 DECAPx2_ASAP7_75t_R FILLER_147_456 ();
 DECAPx4_ASAP7_75t_R FILLER_147_483 ();
 FILLER_ASAP7_75t_R FILLER_147_493 ();
 DECAPx10_ASAP7_75t_R FILLER_147_505 ();
 DECAPx10_ASAP7_75t_R FILLER_147_527 ();
 DECAPx10_ASAP7_75t_R FILLER_147_549 ();
 DECAPx10_ASAP7_75t_R FILLER_147_571 ();
 DECAPx10_ASAP7_75t_R FILLER_147_593 ();
 DECAPx1_ASAP7_75t_R FILLER_147_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_619 ();
 DECAPx2_ASAP7_75t_R FILLER_147_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_632 ();
 DECAPx10_ASAP7_75t_R FILLER_147_640 ();
 DECAPx10_ASAP7_75t_R FILLER_147_662 ();
 DECAPx10_ASAP7_75t_R FILLER_147_684 ();
 DECAPx10_ASAP7_75t_R FILLER_147_706 ();
 DECAPx10_ASAP7_75t_R FILLER_147_728 ();
 DECAPx10_ASAP7_75t_R FILLER_147_750 ();
 DECAPx10_ASAP7_75t_R FILLER_147_772 ();
 DECAPx1_ASAP7_75t_R FILLER_147_794 ();
 DECAPx10_ASAP7_75t_R FILLER_147_806 ();
 DECAPx10_ASAP7_75t_R FILLER_147_828 ();
 DECAPx10_ASAP7_75t_R FILLER_147_850 ();
 DECAPx4_ASAP7_75t_R FILLER_147_872 ();
 FILLER_ASAP7_75t_R FILLER_147_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_884 ();
 DECAPx2_ASAP7_75t_R FILLER_147_891 ();
 FILLER_ASAP7_75t_R FILLER_147_897 ();
 DECAPx6_ASAP7_75t_R FILLER_147_907 ();
 FILLER_ASAP7_75t_R FILLER_147_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_923 ();
 DECAPx10_ASAP7_75t_R FILLER_147_926 ();
 DECAPx10_ASAP7_75t_R FILLER_147_948 ();
 DECAPx10_ASAP7_75t_R FILLER_147_970 ();
 DECAPx10_ASAP7_75t_R FILLER_147_992 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1014 ();
 FILLER_ASAP7_75t_R FILLER_147_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1071 ();
 FILLER_ASAP7_75t_R FILLER_147_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1087 ();
 FILLER_ASAP7_75t_R FILLER_147_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1204 ();
 FILLER_ASAP7_75t_R FILLER_147_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_148_2 ();
 DECAPx10_ASAP7_75t_R FILLER_148_24 ();
 DECAPx10_ASAP7_75t_R FILLER_148_46 ();
 DECAPx6_ASAP7_75t_R FILLER_148_68 ();
 DECAPx2_ASAP7_75t_R FILLER_148_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_88 ();
 DECAPx6_ASAP7_75t_R FILLER_148_92 ();
 DECAPx2_ASAP7_75t_R FILLER_148_106 ();
 DECAPx4_ASAP7_75t_R FILLER_148_124 ();
 FILLER_ASAP7_75t_R FILLER_148_165 ();
 DECAPx10_ASAP7_75t_R FILLER_148_173 ();
 DECAPx10_ASAP7_75t_R FILLER_148_195 ();
 DECAPx2_ASAP7_75t_R FILLER_148_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_223 ();
 DECAPx2_ASAP7_75t_R FILLER_148_258 ();
 DECAPx4_ASAP7_75t_R FILLER_148_267 ();
 FILLER_ASAP7_75t_R FILLER_148_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_279 ();
 DECAPx10_ASAP7_75t_R FILLER_148_283 ();
 DECAPx1_ASAP7_75t_R FILLER_148_305 ();
 DECAPx6_ASAP7_75t_R FILLER_148_319 ();
 DECAPx2_ASAP7_75t_R FILLER_148_333 ();
 DECAPx6_ASAP7_75t_R FILLER_148_349 ();
 DECAPx1_ASAP7_75t_R FILLER_148_377 ();
 DECAPx10_ASAP7_75t_R FILLER_148_403 ();
 DECAPx4_ASAP7_75t_R FILLER_148_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_435 ();
 DECAPx6_ASAP7_75t_R FILLER_148_442 ();
 DECAPx2_ASAP7_75t_R FILLER_148_456 ();
 DECAPx10_ASAP7_75t_R FILLER_148_464 ();
 DECAPx10_ASAP7_75t_R FILLER_148_486 ();
 FILLER_ASAP7_75t_R FILLER_148_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_510 ();
 FILLER_ASAP7_75t_R FILLER_148_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_516 ();
 DECAPx6_ASAP7_75t_R FILLER_148_528 ();
 FILLER_ASAP7_75t_R FILLER_148_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_544 ();
 DECAPx2_ASAP7_75t_R FILLER_148_572 ();
 FILLER_ASAP7_75t_R FILLER_148_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_580 ();
 DECAPx10_ASAP7_75t_R FILLER_148_602 ();
 DECAPx6_ASAP7_75t_R FILLER_148_624 ();
 FILLER_ASAP7_75t_R FILLER_148_638 ();
 DECAPx2_ASAP7_75t_R FILLER_148_656 ();
 DECAPx10_ASAP7_75t_R FILLER_148_668 ();
 DECAPx10_ASAP7_75t_R FILLER_148_690 ();
 DECAPx10_ASAP7_75t_R FILLER_148_712 ();
 FILLER_ASAP7_75t_R FILLER_148_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_736 ();
 FILLER_ASAP7_75t_R FILLER_148_751 ();
 DECAPx10_ASAP7_75t_R FILLER_148_759 ();
 DECAPx10_ASAP7_75t_R FILLER_148_781 ();
 DECAPx10_ASAP7_75t_R FILLER_148_803 ();
 DECAPx10_ASAP7_75t_R FILLER_148_825 ();
 DECAPx10_ASAP7_75t_R FILLER_148_847 ();
 DECAPx6_ASAP7_75t_R FILLER_148_869 ();
 FILLER_ASAP7_75t_R FILLER_148_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_885 ();
 DECAPx10_ASAP7_75t_R FILLER_148_893 ();
 DECAPx10_ASAP7_75t_R FILLER_148_915 ();
 DECAPx1_ASAP7_75t_R FILLER_148_937 ();
 DECAPx10_ASAP7_75t_R FILLER_148_951 ();
 FILLER_ASAP7_75t_R FILLER_148_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_981 ();
 DECAPx1_ASAP7_75t_R FILLER_148_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_994 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1127 ();
 FILLER_ASAP7_75t_R FILLER_148_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1156 ();
 FILLER_ASAP7_75t_R FILLER_148_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_149_2 ();
 DECAPx10_ASAP7_75t_R FILLER_149_24 ();
 DECAPx10_ASAP7_75t_R FILLER_149_46 ();
 DECAPx2_ASAP7_75t_R FILLER_149_68 ();
 DECAPx4_ASAP7_75t_R FILLER_149_100 ();
 FILLER_ASAP7_75t_R FILLER_149_110 ();
 DECAPx2_ASAP7_75t_R FILLER_149_118 ();
 FILLER_ASAP7_75t_R FILLER_149_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_126 ();
 DECAPx2_ASAP7_75t_R FILLER_149_133 ();
 FILLER_ASAP7_75t_R FILLER_149_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_141 ();
 DECAPx4_ASAP7_75t_R FILLER_149_174 ();
 DECAPx6_ASAP7_75t_R FILLER_149_191 ();
 DECAPx1_ASAP7_75t_R FILLER_149_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_215 ();
 DECAPx1_ASAP7_75t_R FILLER_149_223 ();
 DECAPx4_ASAP7_75t_R FILLER_149_233 ();
 FILLER_ASAP7_75t_R FILLER_149_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_245 ();
 DECAPx10_ASAP7_75t_R FILLER_149_249 ();
 DECAPx10_ASAP7_75t_R FILLER_149_271 ();
 DECAPx4_ASAP7_75t_R FILLER_149_300 ();
 FILLER_ASAP7_75t_R FILLER_149_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_312 ();
 DECAPx1_ASAP7_75t_R FILLER_149_353 ();
 FILLER_ASAP7_75t_R FILLER_149_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_375 ();
 DECAPx6_ASAP7_75t_R FILLER_149_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_406 ();
 FILLER_ASAP7_75t_R FILLER_149_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_421 ();
 DECAPx2_ASAP7_75t_R FILLER_149_428 ();
 DECAPx10_ASAP7_75t_R FILLER_149_446 ();
 DECAPx6_ASAP7_75t_R FILLER_149_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_510 ();
 FILLER_ASAP7_75t_R FILLER_149_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_555 ();
 DECAPx6_ASAP7_75t_R FILLER_149_594 ();
 FILLER_ASAP7_75t_R FILLER_149_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_610 ();
 DECAPx6_ASAP7_75t_R FILLER_149_620 ();
 DECAPx1_ASAP7_75t_R FILLER_149_634 ();
 DECAPx6_ASAP7_75t_R FILLER_149_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_666 ();
 DECAPx10_ASAP7_75t_R FILLER_149_685 ();
 DECAPx10_ASAP7_75t_R FILLER_149_707 ();
 DECAPx10_ASAP7_75t_R FILLER_149_729 ();
 FILLER_ASAP7_75t_R FILLER_149_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_753 ();
 DECAPx10_ASAP7_75t_R FILLER_149_760 ();
 DECAPx1_ASAP7_75t_R FILLER_149_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_786 ();
 DECAPx4_ASAP7_75t_R FILLER_149_811 ();
 DECAPx10_ASAP7_75t_R FILLER_149_843 ();
 DECAPx10_ASAP7_75t_R FILLER_149_873 ();
 DECAPx10_ASAP7_75t_R FILLER_149_895 ();
 DECAPx2_ASAP7_75t_R FILLER_149_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_923 ();
 DECAPx10_ASAP7_75t_R FILLER_149_926 ();
 DECAPx10_ASAP7_75t_R FILLER_149_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_970 ();
 DECAPx10_ASAP7_75t_R FILLER_149_977 ();
 DECAPx4_ASAP7_75t_R FILLER_149_999 ();
 FILLER_ASAP7_75t_R FILLER_149_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1110 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1126 ();
 FILLER_ASAP7_75t_R FILLER_149_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1188 ();
 FILLER_ASAP7_75t_R FILLER_149_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1232 ();
 FILLER_ASAP7_75t_R FILLER_149_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1276 ();
 FILLER_ASAP7_75t_R FILLER_149_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_150_2 ();
 DECAPx10_ASAP7_75t_R FILLER_150_24 ();
 DECAPx10_ASAP7_75t_R FILLER_150_46 ();
 DECAPx10_ASAP7_75t_R FILLER_150_68 ();
 DECAPx6_ASAP7_75t_R FILLER_150_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_104 ();
 FILLER_ASAP7_75t_R FILLER_150_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_141 ();
 DECAPx10_ASAP7_75t_R FILLER_150_148 ();
 DECAPx10_ASAP7_75t_R FILLER_150_170 ();
 DECAPx2_ASAP7_75t_R FILLER_150_192 ();
 FILLER_ASAP7_75t_R FILLER_150_198 ();
 DECAPx10_ASAP7_75t_R FILLER_150_221 ();
 DECAPx6_ASAP7_75t_R FILLER_150_243 ();
 DECAPx6_ASAP7_75t_R FILLER_150_265 ();
 DECAPx6_ASAP7_75t_R FILLER_150_288 ();
 DECAPx1_ASAP7_75t_R FILLER_150_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_314 ();
 DECAPx2_ASAP7_75t_R FILLER_150_324 ();
 FILLER_ASAP7_75t_R FILLER_150_330 ();
 DECAPx2_ASAP7_75t_R FILLER_150_354 ();
 FILLER_ASAP7_75t_R FILLER_150_360 ();
 DECAPx4_ASAP7_75t_R FILLER_150_370 ();
 FILLER_ASAP7_75t_R FILLER_150_380 ();
 DECAPx10_ASAP7_75t_R FILLER_150_390 ();
 DECAPx2_ASAP7_75t_R FILLER_150_412 ();
 FILLER_ASAP7_75t_R FILLER_150_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_438 ();
 DECAPx2_ASAP7_75t_R FILLER_150_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_461 ();
 DECAPx1_ASAP7_75t_R FILLER_150_464 ();
 DECAPx10_ASAP7_75t_R FILLER_150_474 ();
 DECAPx4_ASAP7_75t_R FILLER_150_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_506 ();
 DECAPx1_ASAP7_75t_R FILLER_150_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_519 ();
 DECAPx2_ASAP7_75t_R FILLER_150_528 ();
 DECAPx6_ASAP7_75t_R FILLER_150_548 ();
 FILLER_ASAP7_75t_R FILLER_150_562 ();
 DECAPx6_ASAP7_75t_R FILLER_150_567 ();
 DECAPx10_ASAP7_75t_R FILLER_150_598 ();
 DECAPx10_ASAP7_75t_R FILLER_150_620 ();
 FILLER_ASAP7_75t_R FILLER_150_642 ();
 DECAPx2_ASAP7_75t_R FILLER_150_650 ();
 DECAPx6_ASAP7_75t_R FILLER_150_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_684 ();
 DECAPx2_ASAP7_75t_R FILLER_150_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_700 ();
 DECAPx10_ASAP7_75t_R FILLER_150_707 ();
 DECAPx10_ASAP7_75t_R FILLER_150_729 ();
 FILLER_ASAP7_75t_R FILLER_150_751 ();
 DECAPx10_ASAP7_75t_R FILLER_150_759 ();
 DECAPx10_ASAP7_75t_R FILLER_150_781 ();
 DECAPx1_ASAP7_75t_R FILLER_150_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_807 ();
 DECAPx10_ASAP7_75t_R FILLER_150_817 ();
 DECAPx10_ASAP7_75t_R FILLER_150_839 ();
 DECAPx10_ASAP7_75t_R FILLER_150_861 ();
 DECAPx10_ASAP7_75t_R FILLER_150_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_905 ();
 DECAPx10_ASAP7_75t_R FILLER_150_916 ();
 DECAPx6_ASAP7_75t_R FILLER_150_938 ();
 DECAPx2_ASAP7_75t_R FILLER_150_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_958 ();
 DECAPx10_ASAP7_75t_R FILLER_150_969 ();
 DECAPx6_ASAP7_75t_R FILLER_150_991 ();
 FILLER_ASAP7_75t_R FILLER_150_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1046 ();
 FILLER_ASAP7_75t_R FILLER_150_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1190 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1236 ();
 FILLER_ASAP7_75t_R FILLER_150_1242 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1277 ();
 FILLER_ASAP7_75t_R FILLER_150_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_151_2 ();
 DECAPx10_ASAP7_75t_R FILLER_151_24 ();
 DECAPx10_ASAP7_75t_R FILLER_151_46 ();
 DECAPx2_ASAP7_75t_R FILLER_151_68 ();
 DECAPx2_ASAP7_75t_R FILLER_151_100 ();
 FILLER_ASAP7_75t_R FILLER_151_106 ();
 DECAPx2_ASAP7_75t_R FILLER_151_111 ();
 DECAPx1_ASAP7_75t_R FILLER_151_153 ();
 FILLER_ASAP7_75t_R FILLER_151_163 ();
 FILLER_ASAP7_75t_R FILLER_151_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_179 ();
 FILLER_ASAP7_75t_R FILLER_151_205 ();
 FILLER_ASAP7_75t_R FILLER_151_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_216 ();
 DECAPx1_ASAP7_75t_R FILLER_151_229 ();
 DECAPx2_ASAP7_75t_R FILLER_151_239 ();
 FILLER_ASAP7_75t_R FILLER_151_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_294 ();
 DECAPx6_ASAP7_75t_R FILLER_151_298 ();
 DECAPx1_ASAP7_75t_R FILLER_151_312 ();
 DECAPx2_ASAP7_75t_R FILLER_151_324 ();
 FILLER_ASAP7_75t_R FILLER_151_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_332 ();
 DECAPx10_ASAP7_75t_R FILLER_151_355 ();
 DECAPx2_ASAP7_75t_R FILLER_151_377 ();
 DECAPx1_ASAP7_75t_R FILLER_151_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_393 ();
 DECAPx1_ASAP7_75t_R FILLER_151_414 ();
 DECAPx10_ASAP7_75t_R FILLER_151_426 ();
 DECAPx2_ASAP7_75t_R FILLER_151_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_461 ();
 FILLER_ASAP7_75t_R FILLER_151_468 ();
 DECAPx10_ASAP7_75t_R FILLER_151_476 ();
 DECAPx4_ASAP7_75t_R FILLER_151_498 ();
 FILLER_ASAP7_75t_R FILLER_151_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_516 ();
 DECAPx10_ASAP7_75t_R FILLER_151_523 ();
 DECAPx4_ASAP7_75t_R FILLER_151_545 ();
 DECAPx2_ASAP7_75t_R FILLER_151_561 ();
 DECAPx10_ASAP7_75t_R FILLER_151_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_597 ();
 FILLER_ASAP7_75t_R FILLER_151_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_614 ();
 DECAPx6_ASAP7_75t_R FILLER_151_618 ();
 DECAPx2_ASAP7_75t_R FILLER_151_632 ();
 DECAPx6_ASAP7_75t_R FILLER_151_648 ();
 DECAPx1_ASAP7_75t_R FILLER_151_662 ();
 FILLER_ASAP7_75t_R FILLER_151_678 ();
 DECAPx4_ASAP7_75t_R FILLER_151_686 ();
 FILLER_ASAP7_75t_R FILLER_151_696 ();
 DECAPx10_ASAP7_75t_R FILLER_151_704 ();
 DECAPx10_ASAP7_75t_R FILLER_151_726 ();
 DECAPx10_ASAP7_75t_R FILLER_151_748 ();
 DECAPx10_ASAP7_75t_R FILLER_151_770 ();
 DECAPx10_ASAP7_75t_R FILLER_151_792 ();
 DECAPx10_ASAP7_75t_R FILLER_151_814 ();
 DECAPx10_ASAP7_75t_R FILLER_151_836 ();
 DECAPx1_ASAP7_75t_R FILLER_151_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_862 ();
 DECAPx1_ASAP7_75t_R FILLER_151_879 ();
 FILLER_ASAP7_75t_R FILLER_151_889 ();
 DECAPx1_ASAP7_75t_R FILLER_151_897 ();
 DECAPx6_ASAP7_75t_R FILLER_151_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_923 ();
 DECAPx6_ASAP7_75t_R FILLER_151_926 ();
 DECAPx1_ASAP7_75t_R FILLER_151_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_944 ();
 FILLER_ASAP7_75t_R FILLER_151_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_953 ();
 DECAPx10_ASAP7_75t_R FILLER_151_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_996 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1081 ();
 FILLER_ASAP7_75t_R FILLER_151_1097 ();
 FILLER_ASAP7_75t_R FILLER_151_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1202 ();
 FILLER_ASAP7_75t_R FILLER_151_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1216 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_152_2 ();
 DECAPx10_ASAP7_75t_R FILLER_152_24 ();
 DECAPx10_ASAP7_75t_R FILLER_152_46 ();
 DECAPx6_ASAP7_75t_R FILLER_152_68 ();
 DECAPx2_ASAP7_75t_R FILLER_152_82 ();
 FILLER_ASAP7_75t_R FILLER_152_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_93 ();
 FILLER_ASAP7_75t_R FILLER_152_133 ();
 DECAPx6_ASAP7_75t_R FILLER_152_143 ();
 DECAPx2_ASAP7_75t_R FILLER_152_157 ();
 DECAPx2_ASAP7_75t_R FILLER_152_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_175 ();
 DECAPx2_ASAP7_75t_R FILLER_152_189 ();
 FILLER_ASAP7_75t_R FILLER_152_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_211 ();
 DECAPx2_ASAP7_75t_R FILLER_152_219 ();
 DECAPx2_ASAP7_75t_R FILLER_152_239 ();
 FILLER_ASAP7_75t_R FILLER_152_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_247 ();
 DECAPx10_ASAP7_75t_R FILLER_152_271 ();
 DECAPx1_ASAP7_75t_R FILLER_152_293 ();
 DECAPx4_ASAP7_75t_R FILLER_152_323 ();
 FILLER_ASAP7_75t_R FILLER_152_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_335 ();
 DECAPx2_ASAP7_75t_R FILLER_152_343 ();
 FILLER_ASAP7_75t_R FILLER_152_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_351 ();
 DECAPx10_ASAP7_75t_R FILLER_152_355 ();
 DECAPx2_ASAP7_75t_R FILLER_152_385 ();
 FILLER_ASAP7_75t_R FILLER_152_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_393 ();
 FILLER_ASAP7_75t_R FILLER_152_400 ();
 FILLER_ASAP7_75t_R FILLER_152_413 ();
 DECAPx10_ASAP7_75t_R FILLER_152_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_477 ();
 DECAPx6_ASAP7_75t_R FILLER_152_494 ();
 DECAPx2_ASAP7_75t_R FILLER_152_508 ();
 DECAPx4_ASAP7_75t_R FILLER_152_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_530 ();
 DECAPx2_ASAP7_75t_R FILLER_152_552 ();
 FILLER_ASAP7_75t_R FILLER_152_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_560 ();
 DECAPx6_ASAP7_75t_R FILLER_152_585 ();
 DECAPx6_ASAP7_75t_R FILLER_152_620 ();
 DECAPx1_ASAP7_75t_R FILLER_152_634 ();
 DECAPx2_ASAP7_75t_R FILLER_152_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_650 ();
 DECAPx10_ASAP7_75t_R FILLER_152_675 ();
 DECAPx10_ASAP7_75t_R FILLER_152_697 ();
 DECAPx2_ASAP7_75t_R FILLER_152_719 ();
 FILLER_ASAP7_75t_R FILLER_152_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_733 ();
 DECAPx2_ASAP7_75t_R FILLER_152_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_746 ();
 DECAPx10_ASAP7_75t_R FILLER_152_753 ();
 DECAPx10_ASAP7_75t_R FILLER_152_775 ();
 DECAPx4_ASAP7_75t_R FILLER_152_797 ();
 DECAPx10_ASAP7_75t_R FILLER_152_816 ();
 DECAPx10_ASAP7_75t_R FILLER_152_838 ();
 DECAPx10_ASAP7_75t_R FILLER_152_860 ();
 DECAPx10_ASAP7_75t_R FILLER_152_882 ();
 DECAPx6_ASAP7_75t_R FILLER_152_904 ();
 FILLER_ASAP7_75t_R FILLER_152_918 ();
 DECAPx10_ASAP7_75t_R FILLER_152_930 ();
 DECAPx10_ASAP7_75t_R FILLER_152_952 ();
 DECAPx6_ASAP7_75t_R FILLER_152_974 ();
 FILLER_ASAP7_75t_R FILLER_152_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_990 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1118 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1284 ();
 FILLER_ASAP7_75t_R FILLER_152_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_153_2 ();
 DECAPx10_ASAP7_75t_R FILLER_153_24 ();
 DECAPx10_ASAP7_75t_R FILLER_153_46 ();
 DECAPx10_ASAP7_75t_R FILLER_153_68 ();
 DECAPx6_ASAP7_75t_R FILLER_153_90 ();
 DECAPx4_ASAP7_75t_R FILLER_153_107 ();
 FILLER_ASAP7_75t_R FILLER_153_147 ();
 FILLER_ASAP7_75t_R FILLER_153_159 ();
 DECAPx10_ASAP7_75t_R FILLER_153_167 ();
 DECAPx6_ASAP7_75t_R FILLER_153_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_203 ();
 DECAPx2_ASAP7_75t_R FILLER_153_211 ();
 FILLER_ASAP7_75t_R FILLER_153_229 ();
 DECAPx10_ASAP7_75t_R FILLER_153_240 ();
 DECAPx10_ASAP7_75t_R FILLER_153_262 ();
 DECAPx2_ASAP7_75t_R FILLER_153_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_296 ();
 DECAPx2_ASAP7_75t_R FILLER_153_304 ();
 FILLER_ASAP7_75t_R FILLER_153_310 ();
 DECAPx6_ASAP7_75t_R FILLER_153_315 ();
 FILLER_ASAP7_75t_R FILLER_153_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_331 ();
 DECAPx6_ASAP7_75t_R FILLER_153_364 ();
 DECAPx1_ASAP7_75t_R FILLER_153_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_382 ();
 DECAPx6_ASAP7_75t_R FILLER_153_390 ();
 FILLER_ASAP7_75t_R FILLER_153_426 ();
 DECAPx4_ASAP7_75t_R FILLER_153_434 ();
 DECAPx2_ASAP7_75t_R FILLER_153_452 ();
 FILLER_ASAP7_75t_R FILLER_153_458 ();
 DECAPx10_ASAP7_75t_R FILLER_153_490 ();
 DECAPx1_ASAP7_75t_R FILLER_153_512 ();
 FILLER_ASAP7_75t_R FILLER_153_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_526 ();
 FILLER_ASAP7_75t_R FILLER_153_530 ();
 DECAPx10_ASAP7_75t_R FILLER_153_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_563 ();
 DECAPx10_ASAP7_75t_R FILLER_153_570 ();
 FILLER_ASAP7_75t_R FILLER_153_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_594 ();
 DECAPx10_ASAP7_75t_R FILLER_153_617 ();
 DECAPx10_ASAP7_75t_R FILLER_153_639 ();
 DECAPx6_ASAP7_75t_R FILLER_153_661 ();
 FILLER_ASAP7_75t_R FILLER_153_675 ();
 DECAPx10_ASAP7_75t_R FILLER_153_687 ();
 DECAPx6_ASAP7_75t_R FILLER_153_709 ();
 FILLER_ASAP7_75t_R FILLER_153_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_725 ();
 FILLER_ASAP7_75t_R FILLER_153_732 ();
 DECAPx10_ASAP7_75t_R FILLER_153_740 ();
 DECAPx10_ASAP7_75t_R FILLER_153_762 ();
 DECAPx10_ASAP7_75t_R FILLER_153_784 ();
 DECAPx10_ASAP7_75t_R FILLER_153_806 ();
 DECAPx10_ASAP7_75t_R FILLER_153_828 ();
 DECAPx10_ASAP7_75t_R FILLER_153_850 ();
 DECAPx10_ASAP7_75t_R FILLER_153_872 ();
 DECAPx10_ASAP7_75t_R FILLER_153_894 ();
 DECAPx2_ASAP7_75t_R FILLER_153_916 ();
 FILLER_ASAP7_75t_R FILLER_153_922 ();
 DECAPx10_ASAP7_75t_R FILLER_153_926 ();
 DECAPx1_ASAP7_75t_R FILLER_153_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_959 ();
 DECAPx10_ASAP7_75t_R FILLER_153_966 ();
 DECAPx4_ASAP7_75t_R FILLER_153_988 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1093 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1115 ();
 FILLER_ASAP7_75t_R FILLER_153_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1269 ();
 FILLER_ASAP7_75t_R FILLER_153_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_154_2 ();
 DECAPx10_ASAP7_75t_R FILLER_154_24 ();
 DECAPx10_ASAP7_75t_R FILLER_154_46 ();
 DECAPx10_ASAP7_75t_R FILLER_154_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_90 ();
 DECAPx6_ASAP7_75t_R FILLER_154_123 ();
 DECAPx2_ASAP7_75t_R FILLER_154_137 ();
 DECAPx1_ASAP7_75t_R FILLER_154_156 ();
 DECAPx10_ASAP7_75t_R FILLER_154_166 ();
 DECAPx10_ASAP7_75t_R FILLER_154_188 ();
 DECAPx10_ASAP7_75t_R FILLER_154_210 ();
 DECAPx2_ASAP7_75t_R FILLER_154_232 ();
 DECAPx10_ASAP7_75t_R FILLER_154_256 ();
 DECAPx1_ASAP7_75t_R FILLER_154_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_282 ();
 FILLER_ASAP7_75t_R FILLER_154_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_297 ();
 DECAPx6_ASAP7_75t_R FILLER_154_350 ();
 DECAPx6_ASAP7_75t_R FILLER_154_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_416 ();
 DECAPx1_ASAP7_75t_R FILLER_154_424 ();
 FILLER_ASAP7_75t_R FILLER_154_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_438 ();
 DECAPx4_ASAP7_75t_R FILLER_154_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_461 ();
 DECAPx4_ASAP7_75t_R FILLER_154_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_474 ();
 DECAPx6_ASAP7_75t_R FILLER_154_481 ();
 DECAPx1_ASAP7_75t_R FILLER_154_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_520 ();
 DECAPx1_ASAP7_75t_R FILLER_154_527 ();
 FILLER_ASAP7_75t_R FILLER_154_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_541 ();
 DECAPx4_ASAP7_75t_R FILLER_154_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_576 ();
 DECAPx6_ASAP7_75t_R FILLER_154_593 ();
 FILLER_ASAP7_75t_R FILLER_154_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_617 ();
 DECAPx10_ASAP7_75t_R FILLER_154_621 ();
 DECAPx10_ASAP7_75t_R FILLER_154_643 ();
 DECAPx4_ASAP7_75t_R FILLER_154_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_675 ();
 DECAPx4_ASAP7_75t_R FILLER_154_682 ();
 FILLER_ASAP7_75t_R FILLER_154_692 ();
 DECAPx10_ASAP7_75t_R FILLER_154_700 ();
 DECAPx10_ASAP7_75t_R FILLER_154_722 ();
 DECAPx6_ASAP7_75t_R FILLER_154_744 ();
 DECAPx1_ASAP7_75t_R FILLER_154_758 ();
 DECAPx1_ASAP7_75t_R FILLER_154_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_776 ();
 DECAPx10_ASAP7_75t_R FILLER_154_783 ();
 DECAPx6_ASAP7_75t_R FILLER_154_805 ();
 FILLER_ASAP7_75t_R FILLER_154_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_821 ();
 DECAPx10_ASAP7_75t_R FILLER_154_828 ();
 DECAPx4_ASAP7_75t_R FILLER_154_850 ();
 FILLER_ASAP7_75t_R FILLER_154_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_862 ();
 DECAPx10_ASAP7_75t_R FILLER_154_869 ();
 DECAPx10_ASAP7_75t_R FILLER_154_891 ();
 DECAPx10_ASAP7_75t_R FILLER_154_913 ();
 DECAPx6_ASAP7_75t_R FILLER_154_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_949 ();
 FILLER_ASAP7_75t_R FILLER_154_971 ();
 DECAPx10_ASAP7_75t_R FILLER_154_979 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1045 ();
 FILLER_ASAP7_75t_R FILLER_154_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1155 ();
 FILLER_ASAP7_75t_R FILLER_154_1215 ();
 FILLER_ASAP7_75t_R FILLER_154_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1233 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1248 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1276 ();
 FILLER_ASAP7_75t_R FILLER_154_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_155_2 ();
 DECAPx10_ASAP7_75t_R FILLER_155_24 ();
 DECAPx10_ASAP7_75t_R FILLER_155_46 ();
 DECAPx10_ASAP7_75t_R FILLER_155_68 ();
 DECAPx2_ASAP7_75t_R FILLER_155_90 ();
 FILLER_ASAP7_75t_R FILLER_155_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_98 ();
 DECAPx4_ASAP7_75t_R FILLER_155_107 ();
 FILLER_ASAP7_75t_R FILLER_155_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_119 ();
 DECAPx4_ASAP7_75t_R FILLER_155_128 ();
 FILLER_ASAP7_75t_R FILLER_155_138 ();
 FILLER_ASAP7_75t_R FILLER_155_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_154 ();
 FILLER_ASAP7_75t_R FILLER_155_164 ();
 DECAPx1_ASAP7_75t_R FILLER_155_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_184 ();
 DECAPx2_ASAP7_75t_R FILLER_155_194 ();
 DECAPx10_ASAP7_75t_R FILLER_155_215 ();
 FILLER_ASAP7_75t_R FILLER_155_237 ();
 DECAPx4_ASAP7_75t_R FILLER_155_249 ();
 FILLER_ASAP7_75t_R FILLER_155_259 ();
 DECAPx4_ASAP7_75t_R FILLER_155_317 ();
 FILLER_ASAP7_75t_R FILLER_155_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_329 ();
 FILLER_ASAP7_75t_R FILLER_155_333 ();
 DECAPx4_ASAP7_75t_R FILLER_155_341 ();
 FILLER_ASAP7_75t_R FILLER_155_351 ();
 DECAPx6_ASAP7_75t_R FILLER_155_365 ();
 DECAPx1_ASAP7_75t_R FILLER_155_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_383 ();
 DECAPx2_ASAP7_75t_R FILLER_155_391 ();
 FILLER_ASAP7_75t_R FILLER_155_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_399 ();
 DECAPx1_ASAP7_75t_R FILLER_155_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_418 ();
 DECAPx6_ASAP7_75t_R FILLER_155_427 ();
 DECAPx4_ASAP7_75t_R FILLER_155_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_467 ();
 DECAPx6_ASAP7_75t_R FILLER_155_485 ();
 DECAPx1_ASAP7_75t_R FILLER_155_499 ();
 DECAPx1_ASAP7_75t_R FILLER_155_511 ();
 FILLER_ASAP7_75t_R FILLER_155_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_527 ();
 DECAPx6_ASAP7_75t_R FILLER_155_531 ();
 FILLER_ASAP7_75t_R FILLER_155_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_547 ();
 DECAPx4_ASAP7_75t_R FILLER_155_556 ();
 FILLER_ASAP7_75t_R FILLER_155_566 ();
 FILLER_ASAP7_75t_R FILLER_155_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_578 ();
 DECAPx10_ASAP7_75t_R FILLER_155_582 ();
 DECAPx1_ASAP7_75t_R FILLER_155_604 ();
 DECAPx10_ASAP7_75t_R FILLER_155_629 ();
 DECAPx4_ASAP7_75t_R FILLER_155_651 ();
 FILLER_ASAP7_75t_R FILLER_155_661 ();
 DECAPx10_ASAP7_75t_R FILLER_155_669 ();
 DECAPx4_ASAP7_75t_R FILLER_155_691 ();
 FILLER_ASAP7_75t_R FILLER_155_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_703 ();
 DECAPx1_ASAP7_75t_R FILLER_155_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_723 ();
 DECAPx2_ASAP7_75t_R FILLER_155_730 ();
 FILLER_ASAP7_75t_R FILLER_155_736 ();
 DECAPx4_ASAP7_75t_R FILLER_155_748 ();
 FILLER_ASAP7_75t_R FILLER_155_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_760 ();
 DECAPx10_ASAP7_75t_R FILLER_155_775 ();
 DECAPx10_ASAP7_75t_R FILLER_155_797 ();
 DECAPx4_ASAP7_75t_R FILLER_155_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_829 ();
 DECAPx2_ASAP7_75t_R FILLER_155_840 ();
 FILLER_ASAP7_75t_R FILLER_155_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_848 ();
 DECAPx10_ASAP7_75t_R FILLER_155_863 ();
 DECAPx10_ASAP7_75t_R FILLER_155_885 ();
 DECAPx6_ASAP7_75t_R FILLER_155_907 ();
 FILLER_ASAP7_75t_R FILLER_155_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_923 ();
 DECAPx10_ASAP7_75t_R FILLER_155_926 ();
 DECAPx10_ASAP7_75t_R FILLER_155_948 ();
 DECAPx2_ASAP7_75t_R FILLER_155_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_976 ();
 DECAPx6_ASAP7_75t_R FILLER_155_984 ();
 DECAPx1_ASAP7_75t_R FILLER_155_998 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1012 ();
 FILLER_ASAP7_75t_R FILLER_155_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1065 ();
 FILLER_ASAP7_75t_R FILLER_155_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1150 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1166 ();
 FILLER_ASAP7_75t_R FILLER_155_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1269 ();
 FILLER_ASAP7_75t_R FILLER_155_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_156_2 ();
 DECAPx10_ASAP7_75t_R FILLER_156_24 ();
 DECAPx10_ASAP7_75t_R FILLER_156_46 ();
 DECAPx10_ASAP7_75t_R FILLER_156_68 ();
 DECAPx6_ASAP7_75t_R FILLER_156_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_104 ();
 DECAPx2_ASAP7_75t_R FILLER_156_114 ();
 FILLER_ASAP7_75t_R FILLER_156_120 ();
 DECAPx6_ASAP7_75t_R FILLER_156_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_149 ();
 DECAPx2_ASAP7_75t_R FILLER_156_162 ();
 DECAPx2_ASAP7_75t_R FILLER_156_175 ();
 FILLER_ASAP7_75t_R FILLER_156_181 ();
 DECAPx6_ASAP7_75t_R FILLER_156_190 ();
 DECAPx1_ASAP7_75t_R FILLER_156_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_216 ();
 DECAPx10_ASAP7_75t_R FILLER_156_223 ();
 FILLER_ASAP7_75t_R FILLER_156_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_247 ();
 DECAPx10_ASAP7_75t_R FILLER_156_251 ();
 FILLER_ASAP7_75t_R FILLER_156_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_275 ();
 DECAPx2_ASAP7_75t_R FILLER_156_279 ();
 FILLER_ASAP7_75t_R FILLER_156_285 ();
 DECAPx10_ASAP7_75t_R FILLER_156_294 ();
 DECAPx2_ASAP7_75t_R FILLER_156_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_322 ();
 DECAPx10_ASAP7_75t_R FILLER_156_331 ();
 DECAPx6_ASAP7_75t_R FILLER_156_353 ();
 FILLER_ASAP7_75t_R FILLER_156_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_381 ();
 DECAPx10_ASAP7_75t_R FILLER_156_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_411 ();
 DECAPx10_ASAP7_75t_R FILLER_156_419 ();
 DECAPx2_ASAP7_75t_R FILLER_156_441 ();
 FILLER_ASAP7_75t_R FILLER_156_447 ();
 DECAPx2_ASAP7_75t_R FILLER_156_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_461 ();
 DECAPx2_ASAP7_75t_R FILLER_156_464 ();
 FILLER_ASAP7_75t_R FILLER_156_470 ();
 DECAPx6_ASAP7_75t_R FILLER_156_485 ();
 FILLER_ASAP7_75t_R FILLER_156_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_501 ();
 DECAPx6_ASAP7_75t_R FILLER_156_531 ();
 DECAPx2_ASAP7_75t_R FILLER_156_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_551 ();
 FILLER_ASAP7_75t_R FILLER_156_561 ();
 FILLER_ASAP7_75t_R FILLER_156_584 ();
 DECAPx10_ASAP7_75t_R FILLER_156_610 ();
 DECAPx10_ASAP7_75t_R FILLER_156_632 ();
 DECAPx1_ASAP7_75t_R FILLER_156_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_658 ();
 DECAPx10_ASAP7_75t_R FILLER_156_671 ();
 DECAPx4_ASAP7_75t_R FILLER_156_693 ();
 FILLER_ASAP7_75t_R FILLER_156_703 ();
 DECAPx2_ASAP7_75t_R FILLER_156_711 ();
 FILLER_ASAP7_75t_R FILLER_156_717 ();
 DECAPx10_ASAP7_75t_R FILLER_156_725 ();
 DECAPx10_ASAP7_75t_R FILLER_156_747 ();
 DECAPx10_ASAP7_75t_R FILLER_156_769 ();
 DECAPx10_ASAP7_75t_R FILLER_156_791 ();
 DECAPx10_ASAP7_75t_R FILLER_156_813 ();
 DECAPx10_ASAP7_75t_R FILLER_156_835 ();
 DECAPx10_ASAP7_75t_R FILLER_156_857 ();
 DECAPx2_ASAP7_75t_R FILLER_156_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_885 ();
 DECAPx10_ASAP7_75t_R FILLER_156_917 ();
 DECAPx10_ASAP7_75t_R FILLER_156_939 ();
 DECAPx10_ASAP7_75t_R FILLER_156_961 ();
 DECAPx2_ASAP7_75t_R FILLER_156_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_989 ();
 DECAPx2_ASAP7_75t_R FILLER_156_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1045 ();
 FILLER_ASAP7_75t_R FILLER_156_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1080 ();
 FILLER_ASAP7_75t_R FILLER_156_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1113 ();
 FILLER_ASAP7_75t_R FILLER_156_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1136 ();
 FILLER_ASAP7_75t_R FILLER_156_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1173 ();
 FILLER_ASAP7_75t_R FILLER_156_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1225 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_157_2 ();
 DECAPx10_ASAP7_75t_R FILLER_157_24 ();
 DECAPx10_ASAP7_75t_R FILLER_157_46 ();
 DECAPx10_ASAP7_75t_R FILLER_157_68 ();
 DECAPx6_ASAP7_75t_R FILLER_157_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_104 ();
 DECAPx10_ASAP7_75t_R FILLER_157_120 ();
 DECAPx2_ASAP7_75t_R FILLER_157_142 ();
 FILLER_ASAP7_75t_R FILLER_157_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_150 ();
 DECAPx2_ASAP7_75t_R FILLER_157_164 ();
 FILLER_ASAP7_75t_R FILLER_157_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_185 ();
 FILLER_ASAP7_75t_R FILLER_157_195 ();
 DECAPx2_ASAP7_75t_R FILLER_157_212 ();
 DECAPx2_ASAP7_75t_R FILLER_157_225 ();
 FILLER_ASAP7_75t_R FILLER_157_231 ();
 DECAPx2_ASAP7_75t_R FILLER_157_259 ();
 FILLER_ASAP7_75t_R FILLER_157_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_285 ();
 FILLER_ASAP7_75t_R FILLER_157_301 ();
 FILLER_ASAP7_75t_R FILLER_157_339 ();
 DECAPx2_ASAP7_75t_R FILLER_157_355 ();
 FILLER_ASAP7_75t_R FILLER_157_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_363 ();
 FILLER_ASAP7_75t_R FILLER_157_372 ();
 DECAPx2_ASAP7_75t_R FILLER_157_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_385 ();
 DECAPx2_ASAP7_75t_R FILLER_157_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_407 ();
 DECAPx10_ASAP7_75t_R FILLER_157_414 ();
 DECAPx10_ASAP7_75t_R FILLER_157_436 ();
 DECAPx10_ASAP7_75t_R FILLER_157_458 ();
 DECAPx6_ASAP7_75t_R FILLER_157_480 ();
 DECAPx1_ASAP7_75t_R FILLER_157_494 ();
 FILLER_ASAP7_75t_R FILLER_157_544 ();
 DECAPx1_ASAP7_75t_R FILLER_157_560 ();
 DECAPx4_ASAP7_75t_R FILLER_157_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_580 ();
 FILLER_ASAP7_75t_R FILLER_157_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_589 ();
 FILLER_ASAP7_75t_R FILLER_157_598 ();
 DECAPx2_ASAP7_75t_R FILLER_157_606 ();
 FILLER_ASAP7_75t_R FILLER_157_612 ();
 DECAPx6_ASAP7_75t_R FILLER_157_622 ();
 DECAPx1_ASAP7_75t_R FILLER_157_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_640 ();
 DECAPx4_ASAP7_75t_R FILLER_157_651 ();
 DECAPx10_ASAP7_75t_R FILLER_157_667 ();
 DECAPx10_ASAP7_75t_R FILLER_157_689 ();
 DECAPx4_ASAP7_75t_R FILLER_157_711 ();
 FILLER_ASAP7_75t_R FILLER_157_721 ();
 DECAPx10_ASAP7_75t_R FILLER_157_729 ();
 DECAPx10_ASAP7_75t_R FILLER_157_751 ();
 FILLER_ASAP7_75t_R FILLER_157_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_775 ();
 DECAPx4_ASAP7_75t_R FILLER_157_797 ();
 FILLER_ASAP7_75t_R FILLER_157_807 ();
 DECAPx6_ASAP7_75t_R FILLER_157_812 ();
 FILLER_ASAP7_75t_R FILLER_157_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_828 ();
 DECAPx10_ASAP7_75t_R FILLER_157_835 ();
 DECAPx10_ASAP7_75t_R FILLER_157_857 ();
 DECAPx4_ASAP7_75t_R FILLER_157_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_889 ();
 DECAPx1_ASAP7_75t_R FILLER_157_898 ();
 DECAPx6_ASAP7_75t_R FILLER_157_905 ();
 DECAPx1_ASAP7_75t_R FILLER_157_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_923 ();
 DECAPx6_ASAP7_75t_R FILLER_157_926 ();
 FILLER_ASAP7_75t_R FILLER_157_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_942 ();
 FILLER_ASAP7_75t_R FILLER_157_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_955 ();
 DECAPx4_ASAP7_75t_R FILLER_157_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_972 ();
 DECAPx10_ASAP7_75t_R FILLER_157_979 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1001 ();
 FILLER_ASAP7_75t_R FILLER_157_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1168 ();
 FILLER_ASAP7_75t_R FILLER_157_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_158_2 ();
 DECAPx10_ASAP7_75t_R FILLER_158_24 ();
 DECAPx10_ASAP7_75t_R FILLER_158_46 ();
 DECAPx10_ASAP7_75t_R FILLER_158_68 ();
 DECAPx4_ASAP7_75t_R FILLER_158_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_100 ();
 DECAPx4_ASAP7_75t_R FILLER_158_114 ();
 DECAPx6_ASAP7_75t_R FILLER_158_131 ();
 DECAPx2_ASAP7_75t_R FILLER_158_151 ();
 DECAPx6_ASAP7_75t_R FILLER_158_163 ();
 FILLER_ASAP7_75t_R FILLER_158_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_179 ();
 DECAPx4_ASAP7_75t_R FILLER_158_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_195 ();
 DECAPx6_ASAP7_75t_R FILLER_158_204 ();
 DECAPx2_ASAP7_75t_R FILLER_158_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_224 ();
 DECAPx4_ASAP7_75t_R FILLER_158_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_249 ();
 DECAPx2_ASAP7_75t_R FILLER_158_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_272 ();
 DECAPx2_ASAP7_75t_R FILLER_158_279 ();
 FILLER_ASAP7_75t_R FILLER_158_285 ();
 DECAPx10_ASAP7_75t_R FILLER_158_300 ();
 DECAPx10_ASAP7_75t_R FILLER_158_322 ();
 DECAPx2_ASAP7_75t_R FILLER_158_376 ();
 FILLER_ASAP7_75t_R FILLER_158_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_413 ();
 DECAPx1_ASAP7_75t_R FILLER_158_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_425 ();
 FILLER_ASAP7_75t_R FILLER_158_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_437 ();
 DECAPx2_ASAP7_75t_R FILLER_158_446 ();
 FILLER_ASAP7_75t_R FILLER_158_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_461 ();
 DECAPx10_ASAP7_75t_R FILLER_158_480 ();
 DECAPx1_ASAP7_75t_R FILLER_158_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_506 ();
 DECAPx10_ASAP7_75t_R FILLER_158_558 ();
 DECAPx4_ASAP7_75t_R FILLER_158_580 ();
 FILLER_ASAP7_75t_R FILLER_158_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_592 ();
 DECAPx4_ASAP7_75t_R FILLER_158_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_609 ();
 DECAPx10_ASAP7_75t_R FILLER_158_634 ();
 DECAPx2_ASAP7_75t_R FILLER_158_656 ();
 FILLER_ASAP7_75t_R FILLER_158_662 ();
 DECAPx6_ASAP7_75t_R FILLER_158_674 ();
 DECAPx2_ASAP7_75t_R FILLER_158_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_694 ();
 DECAPx10_ASAP7_75t_R FILLER_158_703 ();
 DECAPx10_ASAP7_75t_R FILLER_158_725 ();
 DECAPx6_ASAP7_75t_R FILLER_158_747 ();
 DECAPx2_ASAP7_75t_R FILLER_158_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_767 ();
 DECAPx6_ASAP7_75t_R FILLER_158_776 ();
 DECAPx1_ASAP7_75t_R FILLER_158_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_794 ();
 FILLER_ASAP7_75t_R FILLER_158_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_821 ();
 DECAPx10_ASAP7_75t_R FILLER_158_846 ();
 DECAPx6_ASAP7_75t_R FILLER_158_868 ();
 DECAPx10_ASAP7_75t_R FILLER_158_892 ();
 DECAPx10_ASAP7_75t_R FILLER_158_914 ();
 DECAPx6_ASAP7_75t_R FILLER_158_936 ();
 DECAPx2_ASAP7_75t_R FILLER_158_950 ();
 DECAPx10_ASAP7_75t_R FILLER_158_962 ();
 DECAPx10_ASAP7_75t_R FILLER_158_984 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1034 ();
 FILLER_ASAP7_75t_R FILLER_158_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1069 ();
 FILLER_ASAP7_75t_R FILLER_158_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1122 ();
 FILLER_ASAP7_75t_R FILLER_158_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_159_2 ();
 DECAPx10_ASAP7_75t_R FILLER_159_24 ();
 DECAPx10_ASAP7_75t_R FILLER_159_46 ();
 DECAPx6_ASAP7_75t_R FILLER_159_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_82 ();
 DECAPx4_ASAP7_75t_R FILLER_159_86 ();
 FILLER_ASAP7_75t_R FILLER_159_96 ();
 DECAPx6_ASAP7_75t_R FILLER_159_116 ();
 DECAPx1_ASAP7_75t_R FILLER_159_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_134 ();
 DECAPx2_ASAP7_75t_R FILLER_159_148 ();
 FILLER_ASAP7_75t_R FILLER_159_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_156 ();
 DECAPx4_ASAP7_75t_R FILLER_159_164 ();
 FILLER_ASAP7_75t_R FILLER_159_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_176 ();
 DECAPx2_ASAP7_75t_R FILLER_159_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_192 ();
 DECAPx10_ASAP7_75t_R FILLER_159_199 ();
 DECAPx4_ASAP7_75t_R FILLER_159_239 ();
 FILLER_ASAP7_75t_R FILLER_159_249 ();
 DECAPx6_ASAP7_75t_R FILLER_159_257 ();
 FILLER_ASAP7_75t_R FILLER_159_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_285 ();
 FILLER_ASAP7_75t_R FILLER_159_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_294 ();
 DECAPx4_ASAP7_75t_R FILLER_159_298 ();
 DECAPx1_ASAP7_75t_R FILLER_159_314 ();
 DECAPx10_ASAP7_75t_R FILLER_159_325 ();
 DECAPx4_ASAP7_75t_R FILLER_159_347 ();
 FILLER_ASAP7_75t_R FILLER_159_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_359 ();
 DECAPx4_ASAP7_75t_R FILLER_159_366 ();
 FILLER_ASAP7_75t_R FILLER_159_376 ();
 DECAPx2_ASAP7_75t_R FILLER_159_391 ();
 FILLER_ASAP7_75t_R FILLER_159_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_407 ();
 DECAPx2_ASAP7_75t_R FILLER_159_415 ();
 FILLER_ASAP7_75t_R FILLER_159_421 ();
 FILLER_ASAP7_75t_R FILLER_159_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_434 ();
 DECAPx6_ASAP7_75t_R FILLER_159_480 ();
 DECAPx2_ASAP7_75t_R FILLER_159_494 ();
 DECAPx4_ASAP7_75t_R FILLER_159_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_553 ();
 FILLER_ASAP7_75t_R FILLER_159_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_564 ();
 DECAPx1_ASAP7_75t_R FILLER_159_576 ();
 DECAPx2_ASAP7_75t_R FILLER_159_587 ();
 FILLER_ASAP7_75t_R FILLER_159_593 ();
 DECAPx10_ASAP7_75t_R FILLER_159_601 ();
 DECAPx10_ASAP7_75t_R FILLER_159_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_645 ();
 DECAPx10_ASAP7_75t_R FILLER_159_652 ();
 DECAPx10_ASAP7_75t_R FILLER_159_674 ();
 DECAPx1_ASAP7_75t_R FILLER_159_696 ();
 DECAPx10_ASAP7_75t_R FILLER_159_706 ();
 DECAPx10_ASAP7_75t_R FILLER_159_728 ();
 DECAPx10_ASAP7_75t_R FILLER_159_750 ();
 DECAPx6_ASAP7_75t_R FILLER_159_772 ();
 DECAPx1_ASAP7_75t_R FILLER_159_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_790 ();
 DECAPx6_ASAP7_75t_R FILLER_159_812 ();
 DECAPx10_ASAP7_75t_R FILLER_159_834 ();
 DECAPx10_ASAP7_75t_R FILLER_159_856 ();
 DECAPx6_ASAP7_75t_R FILLER_159_878 ();
 DECAPx4_ASAP7_75t_R FILLER_159_902 ();
 DECAPx6_ASAP7_75t_R FILLER_159_926 ();
 FILLER_ASAP7_75t_R FILLER_159_940 ();
 DECAPx2_ASAP7_75t_R FILLER_159_949 ();
 DECAPx10_ASAP7_75t_R FILLER_159_961 ();
 DECAPx10_ASAP7_75t_R FILLER_159_983 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1005 ();
 FILLER_ASAP7_75t_R FILLER_159_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1013 ();
 FILLER_ASAP7_75t_R FILLER_159_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1036 ();
 FILLER_ASAP7_75t_R FILLER_159_1042 ();
 FILLER_ASAP7_75t_R FILLER_159_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1167 ();
 FILLER_ASAP7_75t_R FILLER_159_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1214 ();
 FILLER_ASAP7_75t_R FILLER_159_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_160_2 ();
 DECAPx10_ASAP7_75t_R FILLER_160_24 ();
 DECAPx10_ASAP7_75t_R FILLER_160_46 ();
 DECAPx4_ASAP7_75t_R FILLER_160_94 ();
 FILLER_ASAP7_75t_R FILLER_160_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_106 ();
 FILLER_ASAP7_75t_R FILLER_160_142 ();
 DECAPx1_ASAP7_75t_R FILLER_160_156 ();
 DECAPx10_ASAP7_75t_R FILLER_160_170 ();
 FILLER_ASAP7_75t_R FILLER_160_192 ();
 DECAPx2_ASAP7_75t_R FILLER_160_200 ();
 FILLER_ASAP7_75t_R FILLER_160_206 ();
 DECAPx6_ASAP7_75t_R FILLER_160_214 ();
 FILLER_ASAP7_75t_R FILLER_160_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_230 ();
 DECAPx2_ASAP7_75t_R FILLER_160_237 ();
 FILLER_ASAP7_75t_R FILLER_160_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_251 ();
 DECAPx10_ASAP7_75t_R FILLER_160_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_280 ();
 FILLER_ASAP7_75t_R FILLER_160_307 ();
 FILLER_ASAP7_75t_R FILLER_160_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_324 ();
 FILLER_ASAP7_75t_R FILLER_160_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_337 ();
 DECAPx10_ASAP7_75t_R FILLER_160_356 ();
 DECAPx1_ASAP7_75t_R FILLER_160_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_382 ();
 DECAPx1_ASAP7_75t_R FILLER_160_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_397 ();
 DECAPx4_ASAP7_75t_R FILLER_160_410 ();
 FILLER_ASAP7_75t_R FILLER_160_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_428 ();
 FILLER_ASAP7_75t_R FILLER_160_435 ();
 DECAPx6_ASAP7_75t_R FILLER_160_443 ();
 DECAPx1_ASAP7_75t_R FILLER_160_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_461 ();
 DECAPx10_ASAP7_75t_R FILLER_160_471 ();
 DECAPx2_ASAP7_75t_R FILLER_160_493 ();
 DECAPx2_ASAP7_75t_R FILLER_160_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_511 ();
 DECAPx10_ASAP7_75t_R FILLER_160_523 ();
 DECAPx6_ASAP7_75t_R FILLER_160_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_559 ();
 DECAPx10_ASAP7_75t_R FILLER_160_581 ();
 DECAPx10_ASAP7_75t_R FILLER_160_603 ();
 DECAPx2_ASAP7_75t_R FILLER_160_625 ();
 DECAPx4_ASAP7_75t_R FILLER_160_637 ();
 FILLER_ASAP7_75t_R FILLER_160_647 ();
 DECAPx6_ASAP7_75t_R FILLER_160_655 ();
 FILLER_ASAP7_75t_R FILLER_160_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_671 ();
 DECAPx10_ASAP7_75t_R FILLER_160_708 ();
 DECAPx1_ASAP7_75t_R FILLER_160_730 ();
 DECAPx1_ASAP7_75t_R FILLER_160_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_748 ();
 DECAPx10_ASAP7_75t_R FILLER_160_758 ();
 DECAPx10_ASAP7_75t_R FILLER_160_780 ();
 DECAPx10_ASAP7_75t_R FILLER_160_802 ();
 DECAPx10_ASAP7_75t_R FILLER_160_824 ();
 DECAPx10_ASAP7_75t_R FILLER_160_846 ();
 DECAPx10_ASAP7_75t_R FILLER_160_868 ();
 DECAPx10_ASAP7_75t_R FILLER_160_890 ();
 DECAPx10_ASAP7_75t_R FILLER_160_912 ();
 DECAPx10_ASAP7_75t_R FILLER_160_934 ();
 DECAPx6_ASAP7_75t_R FILLER_160_956 ();
 DECAPx2_ASAP7_75t_R FILLER_160_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_976 ();
 DECAPx4_ASAP7_75t_R FILLER_160_983 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1018 ();
 FILLER_ASAP7_75t_R FILLER_160_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1082 ();
 FILLER_ASAP7_75t_R FILLER_160_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1105 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1127 ();
 FILLER_ASAP7_75t_R FILLER_160_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1179 ();
 FILLER_ASAP7_75t_R FILLER_160_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1227 ();
 FILLER_ASAP7_75t_R FILLER_160_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_161_2 ();
 DECAPx10_ASAP7_75t_R FILLER_161_24 ();
 DECAPx10_ASAP7_75t_R FILLER_161_46 ();
 DECAPx10_ASAP7_75t_R FILLER_161_68 ();
 DECAPx6_ASAP7_75t_R FILLER_161_90 ();
 FILLER_ASAP7_75t_R FILLER_161_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_106 ();
 DECAPx2_ASAP7_75t_R FILLER_161_124 ();
 DECAPx6_ASAP7_75t_R FILLER_161_133 ();
 FILLER_ASAP7_75t_R FILLER_161_147 ();
 DECAPx2_ASAP7_75t_R FILLER_161_161 ();
 DECAPx10_ASAP7_75t_R FILLER_161_177 ();
 FILLER_ASAP7_75t_R FILLER_161_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_201 ();
 DECAPx2_ASAP7_75t_R FILLER_161_220 ();
 FILLER_ASAP7_75t_R FILLER_161_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_228 ();
 DECAPx2_ASAP7_75t_R FILLER_161_239 ();
 DECAPx10_ASAP7_75t_R FILLER_161_257 ();
 FILLER_ASAP7_75t_R FILLER_161_279 ();
 DECAPx10_ASAP7_75t_R FILLER_161_289 ();
 DECAPx2_ASAP7_75t_R FILLER_161_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_329 ();
 DECAPx4_ASAP7_75t_R FILLER_161_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_346 ();
 DECAPx6_ASAP7_75t_R FILLER_161_373 ();
 DECAPx2_ASAP7_75t_R FILLER_161_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_393 ();
 DECAPx6_ASAP7_75t_R FILLER_161_400 ();
 DECAPx2_ASAP7_75t_R FILLER_161_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_420 ();
 FILLER_ASAP7_75t_R FILLER_161_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_432 ();
 DECAPx10_ASAP7_75t_R FILLER_161_451 ();
 DECAPx10_ASAP7_75t_R FILLER_161_473 ();
 FILLER_ASAP7_75t_R FILLER_161_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_497 ();
 DECAPx10_ASAP7_75t_R FILLER_161_519 ();
 DECAPx1_ASAP7_75t_R FILLER_161_541 ();
 DECAPx1_ASAP7_75t_R FILLER_161_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_560 ();
 DECAPx10_ASAP7_75t_R FILLER_161_567 ();
 DECAPx2_ASAP7_75t_R FILLER_161_589 ();
 FILLER_ASAP7_75t_R FILLER_161_595 ();
 FILLER_ASAP7_75t_R FILLER_161_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_639 ();
 FILLER_ASAP7_75t_R FILLER_161_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_662 ();
 DECAPx10_ASAP7_75t_R FILLER_161_673 ();
 DECAPx1_ASAP7_75t_R FILLER_161_695 ();
 DECAPx10_ASAP7_75t_R FILLER_161_705 ();
 DECAPx4_ASAP7_75t_R FILLER_161_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_737 ();
 DECAPx4_ASAP7_75t_R FILLER_161_744 ();
 FILLER_ASAP7_75t_R FILLER_161_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_756 ();
 DECAPx10_ASAP7_75t_R FILLER_161_772 ();
 DECAPx10_ASAP7_75t_R FILLER_161_794 ();
 DECAPx10_ASAP7_75t_R FILLER_161_816 ();
 DECAPx10_ASAP7_75t_R FILLER_161_838 ();
 DECAPx1_ASAP7_75t_R FILLER_161_860 ();
 DECAPx2_ASAP7_75t_R FILLER_161_872 ();
 FILLER_ASAP7_75t_R FILLER_161_878 ();
 DECAPx6_ASAP7_75t_R FILLER_161_904 ();
 DECAPx2_ASAP7_75t_R FILLER_161_918 ();
 DECAPx6_ASAP7_75t_R FILLER_161_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_940 ();
 DECAPx4_ASAP7_75t_R FILLER_161_955 ();
 DECAPx4_ASAP7_75t_R FILLER_161_972 ();
 FILLER_ASAP7_75t_R FILLER_161_982 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_161_1073 ();
 FILLER_ASAP7_75t_R FILLER_161_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1151 ();
 FILLER_ASAP7_75t_R FILLER_161_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1195 ();
 FILLER_ASAP7_75t_R FILLER_161_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1276 ();
 FILLER_ASAP7_75t_R FILLER_161_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_162_2 ();
 DECAPx10_ASAP7_75t_R FILLER_162_24 ();
 DECAPx10_ASAP7_75t_R FILLER_162_46 ();
 DECAPx10_ASAP7_75t_R FILLER_162_68 ();
 DECAPx2_ASAP7_75t_R FILLER_162_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_96 ();
 DECAPx2_ASAP7_75t_R FILLER_162_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_115 ();
 DECAPx10_ASAP7_75t_R FILLER_162_122 ();
 FILLER_ASAP7_75t_R FILLER_162_144 ();
 DECAPx6_ASAP7_75t_R FILLER_162_154 ();
 DECAPx1_ASAP7_75t_R FILLER_162_168 ();
 DECAPx6_ASAP7_75t_R FILLER_162_198 ();
 DECAPx10_ASAP7_75t_R FILLER_162_218 ();
 DECAPx10_ASAP7_75t_R FILLER_162_240 ();
 DECAPx1_ASAP7_75t_R FILLER_162_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_266 ();
 DECAPx6_ASAP7_75t_R FILLER_162_273 ();
 FILLER_ASAP7_75t_R FILLER_162_287 ();
 DECAPx10_ASAP7_75t_R FILLER_162_295 ();
 DECAPx6_ASAP7_75t_R FILLER_162_317 ();
 DECAPx1_ASAP7_75t_R FILLER_162_331 ();
 DECAPx6_ASAP7_75t_R FILLER_162_347 ();
 DECAPx2_ASAP7_75t_R FILLER_162_364 ();
 FILLER_ASAP7_75t_R FILLER_162_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_372 ();
 DECAPx1_ASAP7_75t_R FILLER_162_385 ();
 FILLER_ASAP7_75t_R FILLER_162_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_404 ();
 DECAPx4_ASAP7_75t_R FILLER_162_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_425 ();
 DECAPx1_ASAP7_75t_R FILLER_162_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_442 ();
 DECAPx4_ASAP7_75t_R FILLER_162_449 ();
 FILLER_ASAP7_75t_R FILLER_162_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_461 ();
 DECAPx10_ASAP7_75t_R FILLER_162_464 ();
 FILLER_ASAP7_75t_R FILLER_162_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_488 ();
 DECAPx6_ASAP7_75t_R FILLER_162_507 ();
 DECAPx1_ASAP7_75t_R FILLER_162_521 ();
 FILLER_ASAP7_75t_R FILLER_162_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_535 ();
 FILLER_ASAP7_75t_R FILLER_162_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_541 ();
 FILLER_ASAP7_75t_R FILLER_162_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_550 ();
 DECAPx6_ASAP7_75t_R FILLER_162_572 ();
 FILLER_ASAP7_75t_R FILLER_162_586 ();
 DECAPx10_ASAP7_75t_R FILLER_162_594 ();
 DECAPx10_ASAP7_75t_R FILLER_162_616 ();
 DECAPx10_ASAP7_75t_R FILLER_162_638 ();
 DECAPx10_ASAP7_75t_R FILLER_162_660 ();
 DECAPx10_ASAP7_75t_R FILLER_162_682 ();
 DECAPx4_ASAP7_75t_R FILLER_162_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_714 ();
 DECAPx10_ASAP7_75t_R FILLER_162_731 ();
 DECAPx10_ASAP7_75t_R FILLER_162_753 ();
 DECAPx10_ASAP7_75t_R FILLER_162_775 ();
 DECAPx6_ASAP7_75t_R FILLER_162_797 ();
 DECAPx2_ASAP7_75t_R FILLER_162_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_817 ();
 DECAPx10_ASAP7_75t_R FILLER_162_824 ();
 DECAPx10_ASAP7_75t_R FILLER_162_846 ();
 DECAPx6_ASAP7_75t_R FILLER_162_868 ();
 DECAPx1_ASAP7_75t_R FILLER_162_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_886 ();
 DECAPx4_ASAP7_75t_R FILLER_162_895 ();
 FILLER_ASAP7_75t_R FILLER_162_905 ();
 DECAPx10_ASAP7_75t_R FILLER_162_917 ();
 DECAPx2_ASAP7_75t_R FILLER_162_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_945 ();
 DECAPx6_ASAP7_75t_R FILLER_162_953 ();
 DECAPx1_ASAP7_75t_R FILLER_162_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1014 ();
 FILLER_ASAP7_75t_R FILLER_162_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1055 ();
 FILLER_ASAP7_75t_R FILLER_162_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1081 ();
 FILLER_ASAP7_75t_R FILLER_162_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1129 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1151 ();
 FILLER_ASAP7_75t_R FILLER_162_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1200 ();
 FILLER_ASAP7_75t_R FILLER_162_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1281 ();
 FILLER_ASAP7_75t_R FILLER_162_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_163_2 ();
 DECAPx10_ASAP7_75t_R FILLER_163_24 ();
 DECAPx10_ASAP7_75t_R FILLER_163_46 ();
 DECAPx1_ASAP7_75t_R FILLER_163_68 ();
 DECAPx4_ASAP7_75t_R FILLER_163_98 ();
 FILLER_ASAP7_75t_R FILLER_163_108 ();
 FILLER_ASAP7_75t_R FILLER_163_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_126 ();
 FILLER_ASAP7_75t_R FILLER_163_136 ();
 DECAPx2_ASAP7_75t_R FILLER_163_146 ();
 DECAPx4_ASAP7_75t_R FILLER_163_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_190 ();
 DECAPx2_ASAP7_75t_R FILLER_163_202 ();
 FILLER_ASAP7_75t_R FILLER_163_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_210 ();
 DECAPx2_ASAP7_75t_R FILLER_163_237 ();
 DECAPx1_ASAP7_75t_R FILLER_163_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_261 ();
 DECAPx1_ASAP7_75t_R FILLER_163_275 ();
 FILLER_ASAP7_75t_R FILLER_163_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_289 ();
 DECAPx2_ASAP7_75t_R FILLER_163_293 ();
 DECAPx10_ASAP7_75t_R FILLER_163_305 ();
 DECAPx2_ASAP7_75t_R FILLER_163_327 ();
 FILLER_ASAP7_75t_R FILLER_163_333 ();
 DECAPx1_ASAP7_75t_R FILLER_163_345 ();
 DECAPx10_ASAP7_75t_R FILLER_163_355 ();
 DECAPx2_ASAP7_75t_R FILLER_163_377 ();
 FILLER_ASAP7_75t_R FILLER_163_383 ();
 DECAPx6_ASAP7_75t_R FILLER_163_392 ();
 FILLER_ASAP7_75t_R FILLER_163_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_408 ();
 DECAPx2_ASAP7_75t_R FILLER_163_423 ();
 FILLER_ASAP7_75t_R FILLER_163_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_431 ();
 DECAPx4_ASAP7_75t_R FILLER_163_439 ();
 DECAPx6_ASAP7_75t_R FILLER_163_494 ();
 FILLER_ASAP7_75t_R FILLER_163_508 ();
 DECAPx10_ASAP7_75t_R FILLER_163_539 ();
 DECAPx6_ASAP7_75t_R FILLER_163_561 ();
 DECAPx1_ASAP7_75t_R FILLER_163_575 ();
 DECAPx6_ASAP7_75t_R FILLER_163_586 ();
 FILLER_ASAP7_75t_R FILLER_163_600 ();
 DECAPx1_ASAP7_75t_R FILLER_163_610 ();
 DECAPx6_ASAP7_75t_R FILLER_163_617 ();
 FILLER_ASAP7_75t_R FILLER_163_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_633 ();
 DECAPx10_ASAP7_75t_R FILLER_163_642 ();
 DECAPx6_ASAP7_75t_R FILLER_163_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_678 ();
 DECAPx6_ASAP7_75t_R FILLER_163_685 ();
 FILLER_ASAP7_75t_R FILLER_163_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_701 ();
 DECAPx1_ASAP7_75t_R FILLER_163_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_718 ();
 DECAPx6_ASAP7_75t_R FILLER_163_734 ();
 DECAPx2_ASAP7_75t_R FILLER_163_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_754 ();
 DECAPx1_ASAP7_75t_R FILLER_163_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_765 ();
 DECAPx10_ASAP7_75t_R FILLER_163_772 ();
 DECAPx10_ASAP7_75t_R FILLER_163_794 ();
 DECAPx1_ASAP7_75t_R FILLER_163_816 ();
 DECAPx2_ASAP7_75t_R FILLER_163_826 ();
 FILLER_ASAP7_75t_R FILLER_163_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_834 ();
 DECAPx10_ASAP7_75t_R FILLER_163_854 ();
 DECAPx1_ASAP7_75t_R FILLER_163_876 ();
 DECAPx6_ASAP7_75t_R FILLER_163_886 ();
 FILLER_ASAP7_75t_R FILLER_163_900 ();
 DECAPx6_ASAP7_75t_R FILLER_163_926 ();
 DECAPx1_ASAP7_75t_R FILLER_163_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_944 ();
 DECAPx6_ASAP7_75t_R FILLER_163_959 ();
 DECAPx1_ASAP7_75t_R FILLER_163_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_977 ();
 DECAPx1_ASAP7_75t_R FILLER_163_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_992 ();
 DECAPx6_ASAP7_75t_R FILLER_163_999 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1026 ();
 FILLER_ASAP7_75t_R FILLER_163_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1083 ();
 FILLER_ASAP7_75t_R FILLER_163_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1105 ();
 FILLER_ASAP7_75t_R FILLER_163_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1184 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1195 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_164_2 ();
 DECAPx10_ASAP7_75t_R FILLER_164_24 ();
 DECAPx10_ASAP7_75t_R FILLER_164_46 ();
 DECAPx6_ASAP7_75t_R FILLER_164_68 ();
 DECAPx1_ASAP7_75t_R FILLER_164_82 ();
 DECAPx10_ASAP7_75t_R FILLER_164_89 ();
 DECAPx2_ASAP7_75t_R FILLER_164_111 ();
 FILLER_ASAP7_75t_R FILLER_164_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_119 ();
 DECAPx10_ASAP7_75t_R FILLER_164_131 ();
 DECAPx10_ASAP7_75t_R FILLER_164_153 ();
 DECAPx1_ASAP7_75t_R FILLER_164_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_179 ();
 DECAPx1_ASAP7_75t_R FILLER_164_192 ();
 DECAPx2_ASAP7_75t_R FILLER_164_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_212 ();
 DECAPx1_ASAP7_75t_R FILLER_164_221 ();
 DECAPx2_ASAP7_75t_R FILLER_164_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_234 ();
 DECAPx6_ASAP7_75t_R FILLER_164_261 ();
 DECAPx4_ASAP7_75t_R FILLER_164_301 ();
 DECAPx1_ASAP7_75t_R FILLER_164_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_318 ();
 DECAPx4_ASAP7_75t_R FILLER_164_331 ();
 DECAPx2_ASAP7_75t_R FILLER_164_347 ();
 FILLER_ASAP7_75t_R FILLER_164_353 ();
 DECAPx2_ASAP7_75t_R FILLER_164_358 ();
 DECAPx6_ASAP7_75t_R FILLER_164_370 ();
 FILLER_ASAP7_75t_R FILLER_164_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_386 ();
 DECAPx4_ASAP7_75t_R FILLER_164_393 ();
 FILLER_ASAP7_75t_R FILLER_164_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_405 ();
 DECAPx1_ASAP7_75t_R FILLER_164_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_420 ();
 FILLER_ASAP7_75t_R FILLER_164_433 ();
 DECAPx2_ASAP7_75t_R FILLER_164_454 ();
 FILLER_ASAP7_75t_R FILLER_164_460 ();
 DECAPx10_ASAP7_75t_R FILLER_164_464 ();
 DECAPx6_ASAP7_75t_R FILLER_164_486 ();
 DECAPx2_ASAP7_75t_R FILLER_164_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_506 ();
 DECAPx2_ASAP7_75t_R FILLER_164_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_528 ();
 DECAPx10_ASAP7_75t_R FILLER_164_535 ();
 FILLER_ASAP7_75t_R FILLER_164_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_559 ();
 DECAPx1_ASAP7_75t_R FILLER_164_568 ();
 FILLER_ASAP7_75t_R FILLER_164_575 ();
 DECAPx1_ASAP7_75t_R FILLER_164_591 ();
 DECAPx10_ASAP7_75t_R FILLER_164_619 ();
 DECAPx10_ASAP7_75t_R FILLER_164_647 ();
 DECAPx6_ASAP7_75t_R FILLER_164_669 ();
 DECAPx10_ASAP7_75t_R FILLER_164_689 ();
 DECAPx10_ASAP7_75t_R FILLER_164_711 ();
 DECAPx4_ASAP7_75t_R FILLER_164_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_743 ();
 DECAPx10_ASAP7_75t_R FILLER_164_753 ();
 DECAPx10_ASAP7_75t_R FILLER_164_775 ();
 DECAPx6_ASAP7_75t_R FILLER_164_797 ();
 DECAPx1_ASAP7_75t_R FILLER_164_811 ();
 DECAPx10_ASAP7_75t_R FILLER_164_825 ();
 DECAPx4_ASAP7_75t_R FILLER_164_847 ();
 FILLER_ASAP7_75t_R FILLER_164_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_859 ();
 DECAPx10_ASAP7_75t_R FILLER_164_870 ();
 DECAPx10_ASAP7_75t_R FILLER_164_892 ();
 DECAPx10_ASAP7_75t_R FILLER_164_914 ();
 DECAPx10_ASAP7_75t_R FILLER_164_936 ();
 DECAPx10_ASAP7_75t_R FILLER_164_958 ();
 FILLER_ASAP7_75t_R FILLER_164_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_982 ();
 DECAPx6_ASAP7_75t_R FILLER_164_993 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1268 ();
 FILLER_ASAP7_75t_R FILLER_164_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_165_2 ();
 DECAPx10_ASAP7_75t_R FILLER_165_24 ();
 DECAPx6_ASAP7_75t_R FILLER_165_46 ();
 DECAPx2_ASAP7_75t_R FILLER_165_60 ();
 DECAPx6_ASAP7_75t_R FILLER_165_104 ();
 DECAPx6_ASAP7_75t_R FILLER_165_127 ();
 DECAPx1_ASAP7_75t_R FILLER_165_141 ();
 DECAPx10_ASAP7_75t_R FILLER_165_151 ();
 DECAPx4_ASAP7_75t_R FILLER_165_173 ();
 FILLER_ASAP7_75t_R FILLER_165_183 ();
 DECAPx6_ASAP7_75t_R FILLER_165_191 ();
 FILLER_ASAP7_75t_R FILLER_165_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_213 ();
 DECAPx2_ASAP7_75t_R FILLER_165_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_230 ();
 FILLER_ASAP7_75t_R FILLER_165_247 ();
 DECAPx2_ASAP7_75t_R FILLER_165_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_268 ();
 DECAPx2_ASAP7_75t_R FILLER_165_279 ();
 FILLER_ASAP7_75t_R FILLER_165_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_334 ();
 FILLER_ASAP7_75t_R FILLER_165_383 ();
 DECAPx6_ASAP7_75t_R FILLER_165_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_406 ();
 DECAPx6_ASAP7_75t_R FILLER_165_417 ();
 DECAPx1_ASAP7_75t_R FILLER_165_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_435 ();
 DECAPx4_ASAP7_75t_R FILLER_165_442 ();
 DECAPx10_ASAP7_75t_R FILLER_165_464 ();
 DECAPx6_ASAP7_75t_R FILLER_165_486 ();
 DECAPx1_ASAP7_75t_R FILLER_165_500 ();
 DECAPx6_ASAP7_75t_R FILLER_165_536 ();
 DECAPx1_ASAP7_75t_R FILLER_165_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_576 ();
 DECAPx10_ASAP7_75t_R FILLER_165_598 ();
 DECAPx6_ASAP7_75t_R FILLER_165_620 ();
 FILLER_ASAP7_75t_R FILLER_165_634 ();
 DECAPx1_ASAP7_75t_R FILLER_165_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_658 ();
 DECAPx2_ASAP7_75t_R FILLER_165_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_681 ();
 FILLER_ASAP7_75t_R FILLER_165_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_690 ();
 DECAPx2_ASAP7_75t_R FILLER_165_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_703 ();
 DECAPx10_ASAP7_75t_R FILLER_165_718 ();
 DECAPx2_ASAP7_75t_R FILLER_165_740 ();
 FILLER_ASAP7_75t_R FILLER_165_746 ();
 DECAPx10_ASAP7_75t_R FILLER_165_763 ();
 DECAPx10_ASAP7_75t_R FILLER_165_785 ();
 DECAPx2_ASAP7_75t_R FILLER_165_807 ();
 DECAPx10_ASAP7_75t_R FILLER_165_821 ();
 DECAPx10_ASAP7_75t_R FILLER_165_843 ();
 DECAPx10_ASAP7_75t_R FILLER_165_865 ();
 DECAPx10_ASAP7_75t_R FILLER_165_887 ();
 DECAPx6_ASAP7_75t_R FILLER_165_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_923 ();
 DECAPx10_ASAP7_75t_R FILLER_165_926 ();
 DECAPx10_ASAP7_75t_R FILLER_165_948 ();
 DECAPx10_ASAP7_75t_R FILLER_165_970 ();
 FILLER_ASAP7_75t_R FILLER_165_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_994 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1027 ();
 FILLER_ASAP7_75t_R FILLER_165_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1147 ();
 FILLER_ASAP7_75t_R FILLER_165_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1168 ();
 FILLER_ASAP7_75t_R FILLER_165_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_166_2 ();
 DECAPx10_ASAP7_75t_R FILLER_166_24 ();
 DECAPx10_ASAP7_75t_R FILLER_166_46 ();
 DECAPx10_ASAP7_75t_R FILLER_166_68 ();
 DECAPx6_ASAP7_75t_R FILLER_166_90 ();
 DECAPx2_ASAP7_75t_R FILLER_166_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_110 ();
 DECAPx2_ASAP7_75t_R FILLER_166_136 ();
 FILLER_ASAP7_75t_R FILLER_166_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_144 ();
 DECAPx10_ASAP7_75t_R FILLER_166_153 ();
 FILLER_ASAP7_75t_R FILLER_166_175 ();
 DECAPx4_ASAP7_75t_R FILLER_166_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_203 ();
 DECAPx2_ASAP7_75t_R FILLER_166_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_216 ();
 DECAPx1_ASAP7_75t_R FILLER_166_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_227 ();
 DECAPx2_ASAP7_75t_R FILLER_166_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_240 ();
 DECAPx6_ASAP7_75t_R FILLER_166_248 ();
 DECAPx6_ASAP7_75t_R FILLER_166_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_288 ();
 DECAPx10_ASAP7_75t_R FILLER_166_299 ();
 DECAPx2_ASAP7_75t_R FILLER_166_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_327 ();
 DECAPx2_ASAP7_75t_R FILLER_166_334 ();
 DECAPx2_ASAP7_75t_R FILLER_166_352 ();
 DECAPx10_ASAP7_75t_R FILLER_166_370 ();
 DECAPx10_ASAP7_75t_R FILLER_166_392 ();
 DECAPx10_ASAP7_75t_R FILLER_166_414 ();
 FILLER_ASAP7_75t_R FILLER_166_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_438 ();
 DECAPx6_ASAP7_75t_R FILLER_166_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_461 ();
 DECAPx10_ASAP7_75t_R FILLER_166_464 ();
 DECAPx10_ASAP7_75t_R FILLER_166_486 ();
 DECAPx6_ASAP7_75t_R FILLER_166_508 ();
 DECAPx1_ASAP7_75t_R FILLER_166_522 ();
 DECAPx10_ASAP7_75t_R FILLER_166_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_554 ();
 DECAPx10_ASAP7_75t_R FILLER_166_561 ();
 DECAPx10_ASAP7_75t_R FILLER_166_583 ();
 DECAPx10_ASAP7_75t_R FILLER_166_605 ();
 DECAPx10_ASAP7_75t_R FILLER_166_627 ();
 DECAPx10_ASAP7_75t_R FILLER_166_649 ();
 DECAPx10_ASAP7_75t_R FILLER_166_671 ();
 DECAPx10_ASAP7_75t_R FILLER_166_693 ();
 DECAPx10_ASAP7_75t_R FILLER_166_715 ();
 DECAPx10_ASAP7_75t_R FILLER_166_737 ();
 DECAPx10_ASAP7_75t_R FILLER_166_759 ();
 DECAPx10_ASAP7_75t_R FILLER_166_781 ();
 DECAPx2_ASAP7_75t_R FILLER_166_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_809 ();
 DECAPx10_ASAP7_75t_R FILLER_166_820 ();
 DECAPx10_ASAP7_75t_R FILLER_166_842 ();
 DECAPx10_ASAP7_75t_R FILLER_166_864 ();
 DECAPx10_ASAP7_75t_R FILLER_166_886 ();
 DECAPx6_ASAP7_75t_R FILLER_166_908 ();
 DECAPx1_ASAP7_75t_R FILLER_166_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_926 ();
 FILLER_ASAP7_75t_R FILLER_166_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_955 ();
 DECAPx10_ASAP7_75t_R FILLER_166_962 ();
 DECAPx6_ASAP7_75t_R FILLER_166_984 ();
 DECAPx2_ASAP7_75t_R FILLER_166_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1142 ();
 FILLER_ASAP7_75t_R FILLER_166_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_167_2 ();
 DECAPx10_ASAP7_75t_R FILLER_167_24 ();
 DECAPx10_ASAP7_75t_R FILLER_167_46 ();
 DECAPx10_ASAP7_75t_R FILLER_167_68 ();
 FILLER_ASAP7_75t_R FILLER_167_90 ();
 FILLER_ASAP7_75t_R FILLER_167_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_106 ();
 DECAPx10_ASAP7_75t_R FILLER_167_116 ();
 DECAPx6_ASAP7_75t_R FILLER_167_138 ();
 FILLER_ASAP7_75t_R FILLER_167_152 ();
 DECAPx2_ASAP7_75t_R FILLER_167_176 ();
 FILLER_ASAP7_75t_R FILLER_167_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_184 ();
 DECAPx10_ASAP7_75t_R FILLER_167_194 ();
 DECAPx6_ASAP7_75t_R FILLER_167_216 ();
 DECAPx2_ASAP7_75t_R FILLER_167_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_236 ();
 DECAPx10_ASAP7_75t_R FILLER_167_243 ();
 DECAPx6_ASAP7_75t_R FILLER_167_265 ();
 DECAPx2_ASAP7_75t_R FILLER_167_279 ();
 DECAPx10_ASAP7_75t_R FILLER_167_299 ();
 DECAPx2_ASAP7_75t_R FILLER_167_321 ();
 FILLER_ASAP7_75t_R FILLER_167_327 ();
 DECAPx10_ASAP7_75t_R FILLER_167_339 ();
 DECAPx2_ASAP7_75t_R FILLER_167_361 ();
 FILLER_ASAP7_75t_R FILLER_167_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_369 ();
 DECAPx4_ASAP7_75t_R FILLER_167_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_393 ();
 DECAPx10_ASAP7_75t_R FILLER_167_400 ();
 DECAPx4_ASAP7_75t_R FILLER_167_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_432 ();
 FILLER_ASAP7_75t_R FILLER_167_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_442 ();
 DECAPx10_ASAP7_75t_R FILLER_167_449 ();
 FILLER_ASAP7_75t_R FILLER_167_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_473 ();
 DECAPx10_ASAP7_75t_R FILLER_167_484 ();
 DECAPx4_ASAP7_75t_R FILLER_167_506 ();
 FILLER_ASAP7_75t_R FILLER_167_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_518 ();
 DECAPx1_ASAP7_75t_R FILLER_167_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_534 ();
 DECAPx10_ASAP7_75t_R FILLER_167_556 ();
 DECAPx6_ASAP7_75t_R FILLER_167_578 ();
 DECAPx2_ASAP7_75t_R FILLER_167_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_598 ();
 DECAPx10_ASAP7_75t_R FILLER_167_607 ();
 DECAPx10_ASAP7_75t_R FILLER_167_629 ();
 DECAPx10_ASAP7_75t_R FILLER_167_651 ();
 DECAPx10_ASAP7_75t_R FILLER_167_673 ();
 DECAPx10_ASAP7_75t_R FILLER_167_695 ();
 DECAPx10_ASAP7_75t_R FILLER_167_717 ();
 DECAPx10_ASAP7_75t_R FILLER_167_739 ();
 DECAPx10_ASAP7_75t_R FILLER_167_761 ();
 DECAPx10_ASAP7_75t_R FILLER_167_783 ();
 DECAPx10_ASAP7_75t_R FILLER_167_805 ();
 DECAPx10_ASAP7_75t_R FILLER_167_827 ();
 DECAPx4_ASAP7_75t_R FILLER_167_849 ();
 FILLER_ASAP7_75t_R FILLER_167_859 ();
 DECAPx10_ASAP7_75t_R FILLER_167_891 ();
 DECAPx4_ASAP7_75t_R FILLER_167_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_923 ();
 DECAPx2_ASAP7_75t_R FILLER_167_933 ();
 DECAPx6_ASAP7_75t_R FILLER_167_945 ();
 DECAPx10_ASAP7_75t_R FILLER_167_965 ();
 DECAPx10_ASAP7_75t_R FILLER_167_987 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1045 ();
 FILLER_ASAP7_75t_R FILLER_167_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1093 ();
 FILLER_ASAP7_75t_R FILLER_167_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1118 ();
 FILLER_ASAP7_75t_R FILLER_167_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1175 ();
 FILLER_ASAP7_75t_R FILLER_167_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1194 ();
 FILLER_ASAP7_75t_R FILLER_167_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1220 ();
 FILLER_ASAP7_75t_R FILLER_167_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_168_2 ();
 DECAPx10_ASAP7_75t_R FILLER_168_24 ();
 DECAPx10_ASAP7_75t_R FILLER_168_46 ();
 DECAPx10_ASAP7_75t_R FILLER_168_68 ();
 DECAPx4_ASAP7_75t_R FILLER_168_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_113 ();
 DECAPx2_ASAP7_75t_R FILLER_168_121 ();
 FILLER_ASAP7_75t_R FILLER_168_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_136 ();
 FILLER_ASAP7_75t_R FILLER_168_146 ();
 FILLER_ASAP7_75t_R FILLER_168_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_163 ();
 FILLER_ASAP7_75t_R FILLER_168_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_172 ();
 DECAPx10_ASAP7_75t_R FILLER_168_185 ();
 DECAPx6_ASAP7_75t_R FILLER_168_207 ();
 DECAPx1_ASAP7_75t_R FILLER_168_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_225 ();
 DECAPx2_ASAP7_75t_R FILLER_168_232 ();
 FILLER_ASAP7_75t_R FILLER_168_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_240 ();
 DECAPx10_ASAP7_75t_R FILLER_168_247 ();
 DECAPx10_ASAP7_75t_R FILLER_168_269 ();
 FILLER_ASAP7_75t_R FILLER_168_291 ();
 DECAPx2_ASAP7_75t_R FILLER_168_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_312 ();
 DECAPx10_ASAP7_75t_R FILLER_168_319 ();
 DECAPx6_ASAP7_75t_R FILLER_168_341 ();
 DECAPx1_ASAP7_75t_R FILLER_168_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_359 ();
 FILLER_ASAP7_75t_R FILLER_168_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_383 ();
 DECAPx4_ASAP7_75t_R FILLER_168_390 ();
 FILLER_ASAP7_75t_R FILLER_168_400 ();
 DECAPx2_ASAP7_75t_R FILLER_168_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_415 ();
 FILLER_ASAP7_75t_R FILLER_168_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_461 ();
 DECAPx4_ASAP7_75t_R FILLER_168_464 ();
 FILLER_ASAP7_75t_R FILLER_168_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_485 ();
 DECAPx6_ASAP7_75t_R FILLER_168_494 ();
 FILLER_ASAP7_75t_R FILLER_168_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_510 ();
 DECAPx4_ASAP7_75t_R FILLER_168_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_542 ();
 DECAPx2_ASAP7_75t_R FILLER_168_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_560 ();
 DECAPx6_ASAP7_75t_R FILLER_168_575 ();
 DECAPx1_ASAP7_75t_R FILLER_168_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_593 ();
 DECAPx2_ASAP7_75t_R FILLER_168_618 ();
 FILLER_ASAP7_75t_R FILLER_168_624 ();
 DECAPx1_ASAP7_75t_R FILLER_168_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_636 ();
 DECAPx4_ASAP7_75t_R FILLER_168_643 ();
 FILLER_ASAP7_75t_R FILLER_168_653 ();
 DECAPx10_ASAP7_75t_R FILLER_168_661 ();
 DECAPx4_ASAP7_75t_R FILLER_168_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_693 ();
 DECAPx1_ASAP7_75t_R FILLER_168_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_723 ();
 DECAPx10_ASAP7_75t_R FILLER_168_730 ();
 DECAPx4_ASAP7_75t_R FILLER_168_752 ();
 DECAPx6_ASAP7_75t_R FILLER_168_769 ();
 DECAPx2_ASAP7_75t_R FILLER_168_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_789 ();
 DECAPx10_ASAP7_75t_R FILLER_168_804 ();
 DECAPx10_ASAP7_75t_R FILLER_168_826 ();
 DECAPx1_ASAP7_75t_R FILLER_168_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_852 ();
 DECAPx10_ASAP7_75t_R FILLER_168_869 ();
 DECAPx1_ASAP7_75t_R FILLER_168_891 ();
 DECAPx10_ASAP7_75t_R FILLER_168_905 ();
 DECAPx10_ASAP7_75t_R FILLER_168_927 ();
 DECAPx6_ASAP7_75t_R FILLER_168_949 ();
 FILLER_ASAP7_75t_R FILLER_168_963 ();
 DECAPx10_ASAP7_75t_R FILLER_168_977 ();
 DECAPx6_ASAP7_75t_R FILLER_168_999 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1049 ();
 FILLER_ASAP7_75t_R FILLER_168_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1084 ();
 FILLER_ASAP7_75t_R FILLER_168_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1102 ();
 FILLER_ASAP7_75t_R FILLER_168_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1170 ();
 FILLER_ASAP7_75t_R FILLER_168_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1176 ();
 FILLER_ASAP7_75t_R FILLER_168_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_169_2 ();
 DECAPx10_ASAP7_75t_R FILLER_169_24 ();
 DECAPx10_ASAP7_75t_R FILLER_169_46 ();
 DECAPx10_ASAP7_75t_R FILLER_169_68 ();
 DECAPx6_ASAP7_75t_R FILLER_169_90 ();
 FILLER_ASAP7_75t_R FILLER_169_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_106 ();
 DECAPx4_ASAP7_75t_R FILLER_169_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_124 ();
 DECAPx10_ASAP7_75t_R FILLER_169_132 ();
 FILLER_ASAP7_75t_R FILLER_169_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_156 ();
 FILLER_ASAP7_75t_R FILLER_169_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_178 ();
 FILLER_ASAP7_75t_R FILLER_169_197 ();
 DECAPx6_ASAP7_75t_R FILLER_169_211 ();
 FILLER_ASAP7_75t_R FILLER_169_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_227 ();
 DECAPx10_ASAP7_75t_R FILLER_169_234 ();
 DECAPx6_ASAP7_75t_R FILLER_169_256 ();
 DECAPx1_ASAP7_75t_R FILLER_169_270 ();
 DECAPx1_ASAP7_75t_R FILLER_169_280 ();
 DECAPx6_ASAP7_75t_R FILLER_169_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_312 ();
 DECAPx4_ASAP7_75t_R FILLER_169_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_331 ();
 FILLER_ASAP7_75t_R FILLER_169_338 ();
 DECAPx4_ASAP7_75t_R FILLER_169_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_356 ();
 FILLER_ASAP7_75t_R FILLER_169_378 ();
 FILLER_ASAP7_75t_R FILLER_169_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_434 ();
 FILLER_ASAP7_75t_R FILLER_169_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_488 ();
 DECAPx10_ASAP7_75t_R FILLER_169_513 ();
 DECAPx2_ASAP7_75t_R FILLER_169_535 ();
 FILLER_ASAP7_75t_R FILLER_169_541 ();
 FILLER_ASAP7_75t_R FILLER_169_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_551 ();
 DECAPx1_ASAP7_75t_R FILLER_169_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_596 ();
 DECAPx10_ASAP7_75t_R FILLER_169_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_625 ();
 DECAPx10_ASAP7_75t_R FILLER_169_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_684 ();
 DECAPx1_ASAP7_75t_R FILLER_169_697 ();
 DECAPx10_ASAP7_75t_R FILLER_169_713 ();
 DECAPx10_ASAP7_75t_R FILLER_169_735 ();
 DECAPx10_ASAP7_75t_R FILLER_169_757 ();
 DECAPx10_ASAP7_75t_R FILLER_169_779 ();
 DECAPx10_ASAP7_75t_R FILLER_169_801 ();
 DECAPx10_ASAP7_75t_R FILLER_169_823 ();
 DECAPx10_ASAP7_75t_R FILLER_169_845 ();
 DECAPx10_ASAP7_75t_R FILLER_169_867 ();
 DECAPx2_ASAP7_75t_R FILLER_169_889 ();
 DECAPx10_ASAP7_75t_R FILLER_169_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_923 ();
 DECAPx10_ASAP7_75t_R FILLER_169_926 ();
 DECAPx10_ASAP7_75t_R FILLER_169_948 ();
 DECAPx10_ASAP7_75t_R FILLER_169_970 ();
 DECAPx10_ASAP7_75t_R FILLER_169_992 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1089 ();
 FILLER_ASAP7_75t_R FILLER_169_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1143 ();
 FILLER_ASAP7_75t_R FILLER_169_1154 ();
 FILLER_ASAP7_75t_R FILLER_169_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_170_2 ();
 DECAPx10_ASAP7_75t_R FILLER_170_24 ();
 DECAPx10_ASAP7_75t_R FILLER_170_46 ();
 DECAPx10_ASAP7_75t_R FILLER_170_68 ();
 DECAPx6_ASAP7_75t_R FILLER_170_90 ();
 DECAPx1_ASAP7_75t_R FILLER_170_104 ();
 FILLER_ASAP7_75t_R FILLER_170_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_150 ();
 DECAPx6_ASAP7_75t_R FILLER_170_157 ();
 DECAPx2_ASAP7_75t_R FILLER_170_171 ();
 DECAPx10_ASAP7_75t_R FILLER_170_190 ();
 DECAPx4_ASAP7_75t_R FILLER_170_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_222 ();
 FILLER_ASAP7_75t_R FILLER_170_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_237 ();
 DECAPx2_ASAP7_75t_R FILLER_170_261 ();
 FILLER_ASAP7_75t_R FILLER_170_267 ();
 DECAPx6_ASAP7_75t_R FILLER_170_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_297 ();
 DECAPx2_ASAP7_75t_R FILLER_170_306 ();
 DECAPx10_ASAP7_75t_R FILLER_170_318 ();
 DECAPx6_ASAP7_75t_R FILLER_170_340 ();
 DECAPx2_ASAP7_75t_R FILLER_170_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_360 ();
 DECAPx2_ASAP7_75t_R FILLER_170_373 ();
 FILLER_ASAP7_75t_R FILLER_170_379 ();
 DECAPx1_ASAP7_75t_R FILLER_170_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_410 ();
 DECAPx6_ASAP7_75t_R FILLER_170_421 ();
 DECAPx1_ASAP7_75t_R FILLER_170_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_439 ();
 DECAPx4_ASAP7_75t_R FILLER_170_452 ();
 DECAPx2_ASAP7_75t_R FILLER_170_464 ();
 DECAPx10_ASAP7_75t_R FILLER_170_476 ();
 DECAPx1_ASAP7_75t_R FILLER_170_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_502 ();
 DECAPx4_ASAP7_75t_R FILLER_170_527 ();
 FILLER_ASAP7_75t_R FILLER_170_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_539 ();
 DECAPx10_ASAP7_75t_R FILLER_170_546 ();
 FILLER_ASAP7_75t_R FILLER_170_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_570 ();
 DECAPx6_ASAP7_75t_R FILLER_170_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_588 ();
 DECAPx10_ASAP7_75t_R FILLER_170_595 ();
 DECAPx6_ASAP7_75t_R FILLER_170_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_631 ();
 DECAPx6_ASAP7_75t_R FILLER_170_672 ();
 DECAPx2_ASAP7_75t_R FILLER_170_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_692 ();
 DECAPx10_ASAP7_75t_R FILLER_170_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_721 ();
 DECAPx10_ASAP7_75t_R FILLER_170_732 ();
 DECAPx1_ASAP7_75t_R FILLER_170_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_758 ();
 DECAPx10_ASAP7_75t_R FILLER_170_767 ();
 DECAPx10_ASAP7_75t_R FILLER_170_789 ();
 DECAPx2_ASAP7_75t_R FILLER_170_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_817 ();
 DECAPx10_ASAP7_75t_R FILLER_170_824 ();
 DECAPx6_ASAP7_75t_R FILLER_170_846 ();
 DECAPx10_ASAP7_75t_R FILLER_170_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_888 ();
 DECAPx1_ASAP7_75t_R FILLER_170_895 ();
 DECAPx6_ASAP7_75t_R FILLER_170_907 ();
 FILLER_ASAP7_75t_R FILLER_170_941 ();
 DECAPx10_ASAP7_75t_R FILLER_170_951 ();
 DECAPx6_ASAP7_75t_R FILLER_170_973 ();
 DECAPx1_ASAP7_75t_R FILLER_170_987 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1027 ();
 FILLER_ASAP7_75t_R FILLER_170_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1156 ();
 FILLER_ASAP7_75t_R FILLER_170_1167 ();
 FILLER_ASAP7_75t_R FILLER_170_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_171_2 ();
 DECAPx10_ASAP7_75t_R FILLER_171_24 ();
 DECAPx10_ASAP7_75t_R FILLER_171_46 ();
 DECAPx10_ASAP7_75t_R FILLER_171_68 ();
 DECAPx6_ASAP7_75t_R FILLER_171_90 ();
 DECAPx2_ASAP7_75t_R FILLER_171_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_117 ();
 DECAPx4_ASAP7_75t_R FILLER_171_135 ();
 FILLER_ASAP7_75t_R FILLER_171_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_154 ();
 FILLER_ASAP7_75t_R FILLER_171_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_163 ();
 DECAPx2_ASAP7_75t_R FILLER_171_232 ();
 DECAPx2_ASAP7_75t_R FILLER_171_247 ();
 FILLER_ASAP7_75t_R FILLER_171_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_255 ();
 DECAPx10_ASAP7_75t_R FILLER_171_273 ();
 DECAPx10_ASAP7_75t_R FILLER_171_295 ();
 FILLER_ASAP7_75t_R FILLER_171_317 ();
 DECAPx6_ASAP7_75t_R FILLER_171_350 ();
 FILLER_ASAP7_75t_R FILLER_171_364 ();
 DECAPx4_ASAP7_75t_R FILLER_171_372 ();
 DECAPx4_ASAP7_75t_R FILLER_171_389 ();
 DECAPx10_ASAP7_75t_R FILLER_171_405 ();
 DECAPx10_ASAP7_75t_R FILLER_171_427 ();
 DECAPx10_ASAP7_75t_R FILLER_171_449 ();
 DECAPx10_ASAP7_75t_R FILLER_171_471 ();
 DECAPx2_ASAP7_75t_R FILLER_171_493 ();
 FILLER_ASAP7_75t_R FILLER_171_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_501 ();
 DECAPx4_ASAP7_75t_R FILLER_171_518 ();
 FILLER_ASAP7_75t_R FILLER_171_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_530 ();
 DECAPx1_ASAP7_75t_R FILLER_171_539 ();
 DECAPx10_ASAP7_75t_R FILLER_171_572 ();
 DECAPx10_ASAP7_75t_R FILLER_171_594 ();
 DECAPx10_ASAP7_75t_R FILLER_171_626 ();
 DECAPx1_ASAP7_75t_R FILLER_171_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_652 ();
 DECAPx2_ASAP7_75t_R FILLER_171_663 ();
 DECAPx10_ASAP7_75t_R FILLER_171_675 ();
 DECAPx10_ASAP7_75t_R FILLER_171_697 ();
 DECAPx10_ASAP7_75t_R FILLER_171_719 ();
 DECAPx4_ASAP7_75t_R FILLER_171_741 ();
 DECAPx10_ASAP7_75t_R FILLER_171_771 ();
 DECAPx10_ASAP7_75t_R FILLER_171_793 ();
 DECAPx2_ASAP7_75t_R FILLER_171_815 ();
 DECAPx10_ASAP7_75t_R FILLER_171_827 ();
 DECAPx10_ASAP7_75t_R FILLER_171_849 ();
 DECAPx10_ASAP7_75t_R FILLER_171_871 ();
 DECAPx10_ASAP7_75t_R FILLER_171_893 ();
 DECAPx2_ASAP7_75t_R FILLER_171_915 ();
 FILLER_ASAP7_75t_R FILLER_171_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_923 ();
 DECAPx10_ASAP7_75t_R FILLER_171_926 ();
 DECAPx4_ASAP7_75t_R FILLER_171_948 ();
 FILLER_ASAP7_75t_R FILLER_171_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_978 ();
 DECAPx4_ASAP7_75t_R FILLER_171_993 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1011 ();
 FILLER_ASAP7_75t_R FILLER_171_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1032 ();
 FILLER_ASAP7_75t_R FILLER_171_1042 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1066 ();
 FILLER_ASAP7_75t_R FILLER_171_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1089 ();
 FILLER_ASAP7_75t_R FILLER_171_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_172_2 ();
 DECAPx10_ASAP7_75t_R FILLER_172_24 ();
 DECAPx10_ASAP7_75t_R FILLER_172_46 ();
 DECAPx10_ASAP7_75t_R FILLER_172_68 ();
 DECAPx6_ASAP7_75t_R FILLER_172_90 ();
 FILLER_ASAP7_75t_R FILLER_172_104 ();
 DECAPx10_ASAP7_75t_R FILLER_172_120 ();
 DECAPx6_ASAP7_75t_R FILLER_172_142 ();
 FILLER_ASAP7_75t_R FILLER_172_156 ();
 DECAPx10_ASAP7_75t_R FILLER_172_192 ();
 FILLER_ASAP7_75t_R FILLER_172_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_216 ();
 DECAPx2_ASAP7_75t_R FILLER_172_234 ();
 DECAPx1_ASAP7_75t_R FILLER_172_253 ();
 DECAPx10_ASAP7_75t_R FILLER_172_293 ();
 DECAPx10_ASAP7_75t_R FILLER_172_315 ();
 DECAPx1_ASAP7_75t_R FILLER_172_337 ();
 DECAPx4_ASAP7_75t_R FILLER_172_347 ();
 FILLER_ASAP7_75t_R FILLER_172_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_367 ();
 DECAPx10_ASAP7_75t_R FILLER_172_375 ();
 DECAPx10_ASAP7_75t_R FILLER_172_397 ();
 DECAPx6_ASAP7_75t_R FILLER_172_419 ();
 FILLER_ASAP7_75t_R FILLER_172_433 ();
 FILLER_ASAP7_75t_R FILLER_172_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_455 ();
 DECAPx6_ASAP7_75t_R FILLER_172_464 ();
 DECAPx2_ASAP7_75t_R FILLER_172_478 ();
 DECAPx4_ASAP7_75t_R FILLER_172_496 ();
 FILLER_ASAP7_75t_R FILLER_172_506 ();
 DECAPx6_ASAP7_75t_R FILLER_172_514 ();
 DECAPx2_ASAP7_75t_R FILLER_172_528 ();
 FILLER_ASAP7_75t_R FILLER_172_541 ();
 DECAPx6_ASAP7_75t_R FILLER_172_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_560 ();
 FILLER_ASAP7_75t_R FILLER_172_569 ();
 FILLER_ASAP7_75t_R FILLER_172_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_576 ();
 FILLER_ASAP7_75t_R FILLER_172_592 ();
 FILLER_ASAP7_75t_R FILLER_172_603 ();
 DECAPx10_ASAP7_75t_R FILLER_172_616 ();
 FILLER_ASAP7_75t_R FILLER_172_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_648 ();
 DECAPx10_ASAP7_75t_R FILLER_172_655 ();
 DECAPx6_ASAP7_75t_R FILLER_172_677 ();
 DECAPx1_ASAP7_75t_R FILLER_172_691 ();
 DECAPx1_ASAP7_75t_R FILLER_172_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_705 ();
 DECAPx2_ASAP7_75t_R FILLER_172_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_718 ();
 DECAPx1_ASAP7_75t_R FILLER_172_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_730 ();
 DECAPx10_ASAP7_75t_R FILLER_172_745 ();
 DECAPx10_ASAP7_75t_R FILLER_172_767 ();
 DECAPx10_ASAP7_75t_R FILLER_172_789 ();
 DECAPx10_ASAP7_75t_R FILLER_172_811 ();
 DECAPx10_ASAP7_75t_R FILLER_172_843 ();
 DECAPx4_ASAP7_75t_R FILLER_172_865 ();
 FILLER_ASAP7_75t_R FILLER_172_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_877 ();
 DECAPx6_ASAP7_75t_R FILLER_172_903 ();
 FILLER_ASAP7_75t_R FILLER_172_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_919 ();
 DECAPx1_ASAP7_75t_R FILLER_172_926 ();
 DECAPx10_ASAP7_75t_R FILLER_172_942 ();
 DECAPx10_ASAP7_75t_R FILLER_172_964 ();
 DECAPx10_ASAP7_75t_R FILLER_172_986 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1030 ();
 FILLER_ASAP7_75t_R FILLER_172_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1045 ();
 FILLER_ASAP7_75t_R FILLER_172_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1116 ();
 FILLER_ASAP7_75t_R FILLER_172_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1192 ();
 FILLER_ASAP7_75t_R FILLER_172_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1269 ();
 FILLER_ASAP7_75t_R FILLER_172_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_173_2 ();
 DECAPx10_ASAP7_75t_R FILLER_173_24 ();
 DECAPx10_ASAP7_75t_R FILLER_173_46 ();
 DECAPx10_ASAP7_75t_R FILLER_173_68 ();
 DECAPx10_ASAP7_75t_R FILLER_173_90 ();
 DECAPx10_ASAP7_75t_R FILLER_173_112 ();
 DECAPx10_ASAP7_75t_R FILLER_173_134 ();
 FILLER_ASAP7_75t_R FILLER_173_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_158 ();
 DECAPx10_ASAP7_75t_R FILLER_173_181 ();
 FILLER_ASAP7_75t_R FILLER_173_203 ();
 FILLER_ASAP7_75t_R FILLER_173_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_213 ();
 DECAPx1_ASAP7_75t_R FILLER_173_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_230 ();
 FILLER_ASAP7_75t_R FILLER_173_241 ();
 DECAPx2_ASAP7_75t_R FILLER_173_259 ();
 FILLER_ASAP7_75t_R FILLER_173_265 ();
 DECAPx2_ASAP7_75t_R FILLER_173_273 ();
 FILLER_ASAP7_75t_R FILLER_173_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_281 ();
 FILLER_ASAP7_75t_R FILLER_173_289 ();
 DECAPx2_ASAP7_75t_R FILLER_173_310 ();
 FILLER_ASAP7_75t_R FILLER_173_316 ();
 DECAPx2_ASAP7_75t_R FILLER_173_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_330 ();
 FILLER_ASAP7_75t_R FILLER_173_337 ();
 DECAPx6_ASAP7_75t_R FILLER_173_352 ();
 FILLER_ASAP7_75t_R FILLER_173_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_368 ();
 FILLER_ASAP7_75t_R FILLER_173_376 ();
 DECAPx1_ASAP7_75t_R FILLER_173_396 ();
 DECAPx10_ASAP7_75t_R FILLER_173_408 ();
 FILLER_ASAP7_75t_R FILLER_173_430 ();
 DECAPx6_ASAP7_75t_R FILLER_173_456 ();
 DECAPx2_ASAP7_75t_R FILLER_173_470 ();
 DECAPx1_ASAP7_75t_R FILLER_173_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_507 ();
 DECAPx4_ASAP7_75t_R FILLER_173_514 ();
 FILLER_ASAP7_75t_R FILLER_173_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_548 ();
 FILLER_ASAP7_75t_R FILLER_173_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_600 ();
 DECAPx4_ASAP7_75t_R FILLER_173_622 ();
 FILLER_ASAP7_75t_R FILLER_173_632 ();
 DECAPx2_ASAP7_75t_R FILLER_173_646 ();
 DECAPx4_ASAP7_75t_R FILLER_173_658 ();
 FILLER_ASAP7_75t_R FILLER_173_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_678 ();
 DECAPx4_ASAP7_75t_R FILLER_173_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_695 ();
 DECAPx1_ASAP7_75t_R FILLER_173_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_724 ();
 DECAPx10_ASAP7_75t_R FILLER_173_732 ();
 DECAPx10_ASAP7_75t_R FILLER_173_754 ();
 DECAPx10_ASAP7_75t_R FILLER_173_776 ();
 DECAPx10_ASAP7_75t_R FILLER_173_798 ();
 DECAPx10_ASAP7_75t_R FILLER_173_820 ();
 DECAPx10_ASAP7_75t_R FILLER_173_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_864 ();
 DECAPx1_ASAP7_75t_R FILLER_173_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_875 ();
 DECAPx4_ASAP7_75t_R FILLER_173_882 ();
 DECAPx10_ASAP7_75t_R FILLER_173_899 ();
 FILLER_ASAP7_75t_R FILLER_173_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_923 ();
 DECAPx6_ASAP7_75t_R FILLER_173_926 ();
 FILLER_ASAP7_75t_R FILLER_173_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_942 ();
 DECAPx2_ASAP7_75t_R FILLER_173_956 ();
 DECAPx2_ASAP7_75t_R FILLER_173_972 ();
 DECAPx10_ASAP7_75t_R FILLER_173_984 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1050 ();
 FILLER_ASAP7_75t_R FILLER_173_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1128 ();
 FILLER_ASAP7_75t_R FILLER_173_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1195 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_174_2 ();
 DECAPx10_ASAP7_75t_R FILLER_174_24 ();
 DECAPx10_ASAP7_75t_R FILLER_174_46 ();
 DECAPx10_ASAP7_75t_R FILLER_174_68 ();
 DECAPx10_ASAP7_75t_R FILLER_174_90 ();
 DECAPx6_ASAP7_75t_R FILLER_174_112 ();
 DECAPx2_ASAP7_75t_R FILLER_174_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_132 ();
 DECAPx6_ASAP7_75t_R FILLER_174_151 ();
 FILLER_ASAP7_75t_R FILLER_174_165 ();
 DECAPx10_ASAP7_75t_R FILLER_174_173 ();
 DECAPx10_ASAP7_75t_R FILLER_174_195 ();
 DECAPx1_ASAP7_75t_R FILLER_174_217 ();
 DECAPx6_ASAP7_75t_R FILLER_174_232 ();
 DECAPx2_ASAP7_75t_R FILLER_174_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_252 ();
 DECAPx2_ASAP7_75t_R FILLER_174_259 ();
 FILLER_ASAP7_75t_R FILLER_174_265 ();
 DECAPx2_ASAP7_75t_R FILLER_174_275 ();
 DECAPx4_ASAP7_75t_R FILLER_174_307 ();
 FILLER_ASAP7_75t_R FILLER_174_323 ();
 DECAPx1_ASAP7_75t_R FILLER_174_331 ();
 DECAPx1_ASAP7_75t_R FILLER_174_341 ();
 DECAPx1_ASAP7_75t_R FILLER_174_354 ();
 DECAPx6_ASAP7_75t_R FILLER_174_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_379 ();
 DECAPx4_ASAP7_75t_R FILLER_174_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_420 ();
 DECAPx10_ASAP7_75t_R FILLER_174_431 ();
 DECAPx4_ASAP7_75t_R FILLER_174_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_474 ();
 DECAPx10_ASAP7_75t_R FILLER_174_484 ();
 DECAPx2_ASAP7_75t_R FILLER_174_506 ();
 DECAPx6_ASAP7_75t_R FILLER_174_518 ();
 FILLER_ASAP7_75t_R FILLER_174_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_534 ();
 DECAPx10_ASAP7_75t_R FILLER_174_542 ();
 DECAPx10_ASAP7_75t_R FILLER_174_564 ();
 DECAPx10_ASAP7_75t_R FILLER_174_586 ();
 DECAPx10_ASAP7_75t_R FILLER_174_608 ();
 DECAPx10_ASAP7_75t_R FILLER_174_630 ();
 DECAPx4_ASAP7_75t_R FILLER_174_652 ();
 FILLER_ASAP7_75t_R FILLER_174_662 ();
 DECAPx1_ASAP7_75t_R FILLER_174_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_674 ();
 DECAPx10_ASAP7_75t_R FILLER_174_690 ();
 DECAPx6_ASAP7_75t_R FILLER_174_712 ();
 FILLER_ASAP7_75t_R FILLER_174_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_728 ();
 DECAPx10_ASAP7_75t_R FILLER_174_736 ();
 DECAPx10_ASAP7_75t_R FILLER_174_758 ();
 DECAPx10_ASAP7_75t_R FILLER_174_780 ();
 DECAPx10_ASAP7_75t_R FILLER_174_802 ();
 DECAPx10_ASAP7_75t_R FILLER_174_824 ();
 DECAPx10_ASAP7_75t_R FILLER_174_846 ();
 DECAPx10_ASAP7_75t_R FILLER_174_868 ();
 DECAPx10_ASAP7_75t_R FILLER_174_890 ();
 DECAPx10_ASAP7_75t_R FILLER_174_912 ();
 DECAPx10_ASAP7_75t_R FILLER_174_934 ();
 DECAPx1_ASAP7_75t_R FILLER_174_956 ();
 DECAPx10_ASAP7_75t_R FILLER_174_966 ();
 DECAPx2_ASAP7_75t_R FILLER_174_988 ();
 FILLER_ASAP7_75t_R FILLER_174_994 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1096 ();
 FILLER_ASAP7_75t_R FILLER_174_1102 ();
 FILLER_ASAP7_75t_R FILLER_174_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1155 ();
 FILLER_ASAP7_75t_R FILLER_174_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_175_2 ();
 DECAPx10_ASAP7_75t_R FILLER_175_24 ();
 DECAPx10_ASAP7_75t_R FILLER_175_46 ();
 DECAPx10_ASAP7_75t_R FILLER_175_68 ();
 DECAPx6_ASAP7_75t_R FILLER_175_90 ();
 DECAPx2_ASAP7_75t_R FILLER_175_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_110 ();
 DECAPx10_ASAP7_75t_R FILLER_175_151 ();
 DECAPx10_ASAP7_75t_R FILLER_175_173 ();
 DECAPx10_ASAP7_75t_R FILLER_175_195 ();
 FILLER_ASAP7_75t_R FILLER_175_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_219 ();
 DECAPx10_ASAP7_75t_R FILLER_175_236 ();
 DECAPx6_ASAP7_75t_R FILLER_175_258 ();
 DECAPx4_ASAP7_75t_R FILLER_175_284 ();
 FILLER_ASAP7_75t_R FILLER_175_294 ();
 DECAPx1_ASAP7_75t_R FILLER_175_311 ();
 DECAPx2_ASAP7_75t_R FILLER_175_324 ();
 FILLER_ASAP7_75t_R FILLER_175_330 ();
 DECAPx10_ASAP7_75t_R FILLER_175_344 ();
 DECAPx6_ASAP7_75t_R FILLER_175_366 ();
 FILLER_ASAP7_75t_R FILLER_175_380 ();
 FILLER_ASAP7_75t_R FILLER_175_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_390 ();
 DECAPx1_ASAP7_75t_R FILLER_175_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_408 ();
 DECAPx10_ASAP7_75t_R FILLER_175_421 ();
 DECAPx1_ASAP7_75t_R FILLER_175_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_447 ();
 DECAPx1_ASAP7_75t_R FILLER_175_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_458 ();
 DECAPx10_ASAP7_75t_R FILLER_175_474 ();
 DECAPx6_ASAP7_75t_R FILLER_175_496 ();
 DECAPx1_ASAP7_75t_R FILLER_175_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_514 ();
 FILLER_ASAP7_75t_R FILLER_175_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_536 ();
 DECAPx10_ASAP7_75t_R FILLER_175_548 ();
 DECAPx10_ASAP7_75t_R FILLER_175_570 ();
 DECAPx1_ASAP7_75t_R FILLER_175_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_596 ();
 DECAPx10_ASAP7_75t_R FILLER_175_603 ();
 DECAPx2_ASAP7_75t_R FILLER_175_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_631 ();
 DECAPx4_ASAP7_75t_R FILLER_175_640 ();
 DECAPx10_ASAP7_75t_R FILLER_175_658 ();
 DECAPx10_ASAP7_75t_R FILLER_175_680 ();
 DECAPx10_ASAP7_75t_R FILLER_175_702 ();
 DECAPx10_ASAP7_75t_R FILLER_175_724 ();
 DECAPx10_ASAP7_75t_R FILLER_175_746 ();
 DECAPx2_ASAP7_75t_R FILLER_175_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_774 ();
 DECAPx6_ASAP7_75t_R FILLER_175_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_812 ();
 DECAPx10_ASAP7_75t_R FILLER_175_816 ();
 DECAPx10_ASAP7_75t_R FILLER_175_838 ();
 DECAPx10_ASAP7_75t_R FILLER_175_860 ();
 DECAPx10_ASAP7_75t_R FILLER_175_882 ();
 DECAPx6_ASAP7_75t_R FILLER_175_904 ();
 DECAPx2_ASAP7_75t_R FILLER_175_918 ();
 DECAPx6_ASAP7_75t_R FILLER_175_926 ();
 FILLER_ASAP7_75t_R FILLER_175_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_942 ();
 DECAPx10_ASAP7_75t_R FILLER_175_949 ();
 DECAPx2_ASAP7_75t_R FILLER_175_971 ();
 FILLER_ASAP7_75t_R FILLER_175_977 ();
 DECAPx6_ASAP7_75t_R FILLER_175_985 ();
 FILLER_ASAP7_75t_R FILLER_175_999 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_175_1083 ();
 FILLER_ASAP7_75t_R FILLER_175_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1285 ();
 FILLER_ASAP7_75t_R FILLER_175_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_176_2 ();
 DECAPx10_ASAP7_75t_R FILLER_176_24 ();
 DECAPx10_ASAP7_75t_R FILLER_176_46 ();
 DECAPx10_ASAP7_75t_R FILLER_176_68 ();
 DECAPx10_ASAP7_75t_R FILLER_176_90 ();
 DECAPx6_ASAP7_75t_R FILLER_176_112 ();
 DECAPx2_ASAP7_75t_R FILLER_176_126 ();
 DECAPx2_ASAP7_75t_R FILLER_176_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_156 ();
 DECAPx6_ASAP7_75t_R FILLER_176_169 ();
 DECAPx2_ASAP7_75t_R FILLER_176_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_195 ();
 DECAPx6_ASAP7_75t_R FILLER_176_208 ();
 DECAPx2_ASAP7_75t_R FILLER_176_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_228 ();
 DECAPx10_ASAP7_75t_R FILLER_176_233 ();
 DECAPx6_ASAP7_75t_R FILLER_176_255 ();
 FILLER_ASAP7_75t_R FILLER_176_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_271 ();
 DECAPx2_ASAP7_75t_R FILLER_176_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_290 ();
 DECAPx1_ASAP7_75t_R FILLER_176_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_311 ();
 DECAPx10_ASAP7_75t_R FILLER_176_319 ();
 DECAPx6_ASAP7_75t_R FILLER_176_341 ();
 DECAPx2_ASAP7_75t_R FILLER_176_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_361 ();
 DECAPx4_ASAP7_75t_R FILLER_176_371 ();
 FILLER_ASAP7_75t_R FILLER_176_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_383 ();
 DECAPx2_ASAP7_75t_R FILLER_176_396 ();
 DECAPx4_ASAP7_75t_R FILLER_176_412 ();
 FILLER_ASAP7_75t_R FILLER_176_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_446 ();
 DECAPx6_ASAP7_75t_R FILLER_176_479 ();
 DECAPx2_ASAP7_75t_R FILLER_176_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_520 ();
 DECAPx10_ASAP7_75t_R FILLER_176_550 ();
 DECAPx1_ASAP7_75t_R FILLER_176_572 ();
 FILLER_ASAP7_75t_R FILLER_176_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_581 ();
 DECAPx10_ASAP7_75t_R FILLER_176_592 ();
 DECAPx6_ASAP7_75t_R FILLER_176_614 ();
 DECAPx2_ASAP7_75t_R FILLER_176_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_634 ();
 DECAPx10_ASAP7_75t_R FILLER_176_647 ();
 DECAPx10_ASAP7_75t_R FILLER_176_669 ();
 DECAPx4_ASAP7_75t_R FILLER_176_691 ();
 DECAPx2_ASAP7_75t_R FILLER_176_707 ();
 DECAPx10_ASAP7_75t_R FILLER_176_719 ();
 DECAPx4_ASAP7_75t_R FILLER_176_741 ();
 FILLER_ASAP7_75t_R FILLER_176_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_753 ();
 DECAPx10_ASAP7_75t_R FILLER_176_764 ();
 DECAPx6_ASAP7_75t_R FILLER_176_786 ();
 DECAPx2_ASAP7_75t_R FILLER_176_821 ();
 DECAPx6_ASAP7_75t_R FILLER_176_833 ();
 DECAPx1_ASAP7_75t_R FILLER_176_847 ();
 DECAPx4_ASAP7_75t_R FILLER_176_861 ();
 FILLER_ASAP7_75t_R FILLER_176_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_873 ();
 DECAPx10_ASAP7_75t_R FILLER_176_880 ();
 DECAPx10_ASAP7_75t_R FILLER_176_902 ();
 DECAPx1_ASAP7_75t_R FILLER_176_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_928 ();
 DECAPx2_ASAP7_75t_R FILLER_176_935 ();
 FILLER_ASAP7_75t_R FILLER_176_941 ();
 DECAPx4_ASAP7_75t_R FILLER_176_951 ();
 FILLER_ASAP7_75t_R FILLER_176_961 ();
 DECAPx4_ASAP7_75t_R FILLER_176_970 ();
 FILLER_ASAP7_75t_R FILLER_176_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_982 ();
 DECAPx4_ASAP7_75t_R FILLER_176_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1016 ();
 FILLER_ASAP7_75t_R FILLER_176_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1060 ();
 FILLER_ASAP7_75t_R FILLER_176_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_177_2 ();
 DECAPx10_ASAP7_75t_R FILLER_177_24 ();
 DECAPx10_ASAP7_75t_R FILLER_177_46 ();
 DECAPx10_ASAP7_75t_R FILLER_177_68 ();
 DECAPx10_ASAP7_75t_R FILLER_177_90 ();
 DECAPx6_ASAP7_75t_R FILLER_177_112 ();
 DECAPx2_ASAP7_75t_R FILLER_177_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_132 ();
 FILLER_ASAP7_75t_R FILLER_177_139 ();
 DECAPx10_ASAP7_75t_R FILLER_177_147 ();
 DECAPx10_ASAP7_75t_R FILLER_177_169 ();
 DECAPx1_ASAP7_75t_R FILLER_177_191 ();
 DECAPx10_ASAP7_75t_R FILLER_177_207 ();
 DECAPx4_ASAP7_75t_R FILLER_177_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_239 ();
 DECAPx4_ASAP7_75t_R FILLER_177_252 ();
 DECAPx1_ASAP7_75t_R FILLER_177_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_290 ();
 DECAPx6_ASAP7_75t_R FILLER_177_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_312 ();
 DECAPx6_ASAP7_75t_R FILLER_177_318 ();
 DECAPx2_ASAP7_75t_R FILLER_177_332 ();
 FILLER_ASAP7_75t_R FILLER_177_350 ();
 DECAPx10_ASAP7_75t_R FILLER_177_363 ();
 DECAPx10_ASAP7_75t_R FILLER_177_385 ();
 DECAPx6_ASAP7_75t_R FILLER_177_407 ();
 FILLER_ASAP7_75t_R FILLER_177_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_423 ();
 DECAPx4_ASAP7_75t_R FILLER_177_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_446 ();
 DECAPx2_ASAP7_75t_R FILLER_177_453 ();
 FILLER_ASAP7_75t_R FILLER_177_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_461 ();
 DECAPx10_ASAP7_75t_R FILLER_177_471 ();
 FILLER_ASAP7_75t_R FILLER_177_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_495 ();
 DECAPx10_ASAP7_75t_R FILLER_177_517 ();
 DECAPx4_ASAP7_75t_R FILLER_177_539 ();
 FILLER_ASAP7_75t_R FILLER_177_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_559 ();
 FILLER_ASAP7_75t_R FILLER_177_563 ();
 FILLER_ASAP7_75t_R FILLER_177_586 ();
 FILLER_ASAP7_75t_R FILLER_177_610 ();
 DECAPx4_ASAP7_75t_R FILLER_177_639 ();
 FILLER_ASAP7_75t_R FILLER_177_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_651 ();
 DECAPx4_ASAP7_75t_R FILLER_177_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_668 ();
 DECAPx6_ASAP7_75t_R FILLER_177_675 ();
 FILLER_ASAP7_75t_R FILLER_177_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_691 ();
 DECAPx2_ASAP7_75t_R FILLER_177_713 ();
 FILLER_ASAP7_75t_R FILLER_177_725 ();
 DECAPx10_ASAP7_75t_R FILLER_177_737 ();
 DECAPx10_ASAP7_75t_R FILLER_177_759 ();
 DECAPx10_ASAP7_75t_R FILLER_177_781 ();
 DECAPx10_ASAP7_75t_R FILLER_177_803 ();
 DECAPx4_ASAP7_75t_R FILLER_177_831 ();
 DECAPx10_ASAP7_75t_R FILLER_177_853 ();
 DECAPx6_ASAP7_75t_R FILLER_177_875 ();
 DECAPx4_ASAP7_75t_R FILLER_177_896 ();
 FILLER_ASAP7_75t_R FILLER_177_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_908 ();
 FILLER_ASAP7_75t_R FILLER_177_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_923 ();
 FILLER_ASAP7_75t_R FILLER_177_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_938 ();
 DECAPx4_ASAP7_75t_R FILLER_177_948 ();
 FILLER_ASAP7_75t_R FILLER_177_958 ();
 DECAPx4_ASAP7_75t_R FILLER_177_968 ();
 FILLER_ASAP7_75t_R FILLER_177_978 ();
 DECAPx10_ASAP7_75t_R FILLER_177_986 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1183 ();
 FILLER_ASAP7_75t_R FILLER_177_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_178_2 ();
 DECAPx10_ASAP7_75t_R FILLER_178_24 ();
 DECAPx10_ASAP7_75t_R FILLER_178_46 ();
 DECAPx10_ASAP7_75t_R FILLER_178_68 ();
 DECAPx10_ASAP7_75t_R FILLER_178_90 ();
 DECAPx10_ASAP7_75t_R FILLER_178_112 ();
 DECAPx1_ASAP7_75t_R FILLER_178_134 ();
 DECAPx10_ASAP7_75t_R FILLER_178_144 ();
 DECAPx6_ASAP7_75t_R FILLER_178_166 ();
 DECAPx4_ASAP7_75t_R FILLER_178_198 ();
 FILLER_ASAP7_75t_R FILLER_178_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_213 ();
 FILLER_ASAP7_75t_R FILLER_178_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_226 ();
 DECAPx1_ASAP7_75t_R FILLER_178_239 ();
 DECAPx6_ASAP7_75t_R FILLER_178_250 ();
 DECAPx1_ASAP7_75t_R FILLER_178_264 ();
 DECAPx10_ASAP7_75t_R FILLER_178_280 ();
 DECAPx10_ASAP7_75t_R FILLER_178_302 ();
 DECAPx6_ASAP7_75t_R FILLER_178_324 ();
 FILLER_ASAP7_75t_R FILLER_178_338 ();
 FILLER_ASAP7_75t_R FILLER_178_358 ();
 DECAPx1_ASAP7_75t_R FILLER_178_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_371 ();
 DECAPx1_ASAP7_75t_R FILLER_178_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_391 ();
 FILLER_ASAP7_75t_R FILLER_178_399 ();
 DECAPx10_ASAP7_75t_R FILLER_178_407 ();
 DECAPx6_ASAP7_75t_R FILLER_178_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_443 ();
 DECAPx2_ASAP7_75t_R FILLER_178_454 ();
 FILLER_ASAP7_75t_R FILLER_178_460 ();
 FILLER_ASAP7_75t_R FILLER_178_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_472 ();
 DECAPx10_ASAP7_75t_R FILLER_178_480 ();
 DECAPx2_ASAP7_75t_R FILLER_178_502 ();
 FILLER_ASAP7_75t_R FILLER_178_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_521 ();
 DECAPx6_ASAP7_75t_R FILLER_178_530 ();
 FILLER_ASAP7_75t_R FILLER_178_544 ();
 DECAPx1_ASAP7_75t_R FILLER_178_567 ();
 DECAPx1_ASAP7_75t_R FILLER_178_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_607 ();
 DECAPx6_ASAP7_75t_R FILLER_178_619 ();
 FILLER_ASAP7_75t_R FILLER_178_633 ();
 DECAPx2_ASAP7_75t_R FILLER_178_641 ();
 DECAPx4_ASAP7_75t_R FILLER_178_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_669 ();
 FILLER_ASAP7_75t_R FILLER_178_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_684 ();
 DECAPx10_ASAP7_75t_R FILLER_178_697 ();
 DECAPx10_ASAP7_75t_R FILLER_178_719 ();
 FILLER_ASAP7_75t_R FILLER_178_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_743 ();
 DECAPx1_ASAP7_75t_R FILLER_178_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_760 ();
 DECAPx10_ASAP7_75t_R FILLER_178_773 ();
 DECAPx10_ASAP7_75t_R FILLER_178_795 ();
 DECAPx10_ASAP7_75t_R FILLER_178_817 ();
 DECAPx10_ASAP7_75t_R FILLER_178_839 ();
 FILLER_ASAP7_75t_R FILLER_178_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_863 ();
 DECAPx2_ASAP7_75t_R FILLER_178_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_885 ();
 DECAPx10_ASAP7_75t_R FILLER_178_892 ();
 DECAPx4_ASAP7_75t_R FILLER_178_914 ();
 DECAPx10_ASAP7_75t_R FILLER_178_926 ();
 DECAPx10_ASAP7_75t_R FILLER_178_948 ();
 DECAPx4_ASAP7_75t_R FILLER_178_970 ();
 FILLER_ASAP7_75t_R FILLER_178_980 ();
 DECAPx10_ASAP7_75t_R FILLER_178_988 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1010 ();
 FILLER_ASAP7_75t_R FILLER_178_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1028 ();
 FILLER_ASAP7_75t_R FILLER_178_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1040 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1059 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1076 ();
 FILLER_ASAP7_75t_R FILLER_178_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1189 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_179_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_182 ();
 FILLER_ASAP7_75t_R FILLER_179_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_188 ();
 DECAPx2_ASAP7_75t_R FILLER_179_201 ();
 DECAPx1_ASAP7_75t_R FILLER_179_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_247 ();
 DECAPx1_ASAP7_75t_R FILLER_179_260 ();
 DECAPx2_ASAP7_75t_R FILLER_179_273 ();
 FILLER_ASAP7_75t_R FILLER_179_285 ();
 DECAPx10_ASAP7_75t_R FILLER_179_293 ();
 DECAPx2_ASAP7_75t_R FILLER_179_315 ();
 DECAPx6_ASAP7_75t_R FILLER_179_327 ();
 FILLER_ASAP7_75t_R FILLER_179_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_351 ();
 DECAPx10_ASAP7_75t_R FILLER_179_375 ();
 FILLER_ASAP7_75t_R FILLER_179_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_399 ();
 DECAPx10_ASAP7_75t_R FILLER_179_406 ();
 DECAPx6_ASAP7_75t_R FILLER_179_428 ();
 DECAPx2_ASAP7_75t_R FILLER_179_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_448 ();
 DECAPx10_ASAP7_75t_R FILLER_179_455 ();
 DECAPx10_ASAP7_75t_R FILLER_179_477 ();
 DECAPx2_ASAP7_75t_R FILLER_179_499 ();
 FILLER_ASAP7_75t_R FILLER_179_505 ();
 DECAPx6_ASAP7_75t_R FILLER_179_513 ();
 DECAPx1_ASAP7_75t_R FILLER_179_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_546 ();
 DECAPx6_ASAP7_75t_R FILLER_179_553 ();
 DECAPx4_ASAP7_75t_R FILLER_179_573 ();
 DECAPx10_ASAP7_75t_R FILLER_179_589 ();
 DECAPx10_ASAP7_75t_R FILLER_179_611 ();
 DECAPx6_ASAP7_75t_R FILLER_179_633 ();
 DECAPx2_ASAP7_75t_R FILLER_179_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_653 ();
 DECAPx1_ASAP7_75t_R FILLER_179_660 ();
 DECAPx10_ASAP7_75t_R FILLER_179_670 ();
 DECAPx2_ASAP7_75t_R FILLER_179_692 ();
 FILLER_ASAP7_75t_R FILLER_179_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_700 ();
 DECAPx10_ASAP7_75t_R FILLER_179_707 ();
 DECAPx10_ASAP7_75t_R FILLER_179_729 ();
 DECAPx10_ASAP7_75t_R FILLER_179_751 ();
 DECAPx10_ASAP7_75t_R FILLER_179_773 ();
 DECAPx6_ASAP7_75t_R FILLER_179_795 ();
 FILLER_ASAP7_75t_R FILLER_179_809 ();
 DECAPx10_ASAP7_75t_R FILLER_179_815 ();
 DECAPx2_ASAP7_75t_R FILLER_179_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_843 ();
 DECAPx10_ASAP7_75t_R FILLER_179_851 ();
 DECAPx10_ASAP7_75t_R FILLER_179_873 ();
 DECAPx10_ASAP7_75t_R FILLER_179_895 ();
 DECAPx10_ASAP7_75t_R FILLER_179_917 ();
 DECAPx10_ASAP7_75t_R FILLER_179_939 ();
 DECAPx10_ASAP7_75t_R FILLER_179_961 ();
 DECAPx4_ASAP7_75t_R FILLER_179_983 ();
 FILLER_ASAP7_75t_R FILLER_179_993 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1280 ();
 FILLER_ASAP7_75t_R FILLER_179_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_180_172 ();
 FILLER_ASAP7_75t_R FILLER_180_178 ();
 DECAPx6_ASAP7_75t_R FILLER_180_196 ();
 FILLER_ASAP7_75t_R FILLER_180_210 ();
 DECAPx6_ASAP7_75t_R FILLER_180_221 ();
 DECAPx2_ASAP7_75t_R FILLER_180_250 ();
 FILLER_ASAP7_75t_R FILLER_180_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_258 ();
 DECAPx2_ASAP7_75t_R FILLER_180_278 ();
 FILLER_ASAP7_75t_R FILLER_180_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_286 ();
 DECAPx2_ASAP7_75t_R FILLER_180_295 ();
 FILLER_ASAP7_75t_R FILLER_180_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_303 ();
 DECAPx10_ASAP7_75t_R FILLER_180_310 ();
 DECAPx6_ASAP7_75t_R FILLER_180_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_346 ();
 DECAPx2_ASAP7_75t_R FILLER_180_359 ();
 FILLER_ASAP7_75t_R FILLER_180_365 ();
 DECAPx6_ASAP7_75t_R FILLER_180_374 ();
 FILLER_ASAP7_75t_R FILLER_180_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_390 ();
 DECAPx2_ASAP7_75t_R FILLER_180_419 ();
 FILLER_ASAP7_75t_R FILLER_180_425 ();
 DECAPx2_ASAP7_75t_R FILLER_180_439 ();
 DECAPx10_ASAP7_75t_R FILLER_180_478 ();
 DECAPx2_ASAP7_75t_R FILLER_180_500 ();
 FILLER_ASAP7_75t_R FILLER_180_506 ();
 DECAPx4_ASAP7_75t_R FILLER_180_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_524 ();
 DECAPx2_ASAP7_75t_R FILLER_180_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_539 ();
 DECAPx10_ASAP7_75t_R FILLER_180_549 ();
 DECAPx10_ASAP7_75t_R FILLER_180_571 ();
 DECAPx6_ASAP7_75t_R FILLER_180_593 ();
 FILLER_ASAP7_75t_R FILLER_180_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_609 ();
 DECAPx4_ASAP7_75t_R FILLER_180_620 ();
 FILLER_ASAP7_75t_R FILLER_180_630 ();
 DECAPx2_ASAP7_75t_R FILLER_180_634 ();
 DECAPx10_ASAP7_75t_R FILLER_180_647 ();
 DECAPx6_ASAP7_75t_R FILLER_180_675 ();
 DECAPx1_ASAP7_75t_R FILLER_180_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_693 ();
 DECAPx10_ASAP7_75t_R FILLER_180_700 ();
 DECAPx10_ASAP7_75t_R FILLER_180_722 ();
 DECAPx10_ASAP7_75t_R FILLER_180_744 ();
 DECAPx2_ASAP7_75t_R FILLER_180_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_772 ();
 DECAPx10_ASAP7_75t_R FILLER_180_781 ();
 DECAPx1_ASAP7_75t_R FILLER_180_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_828 ();
 DECAPx10_ASAP7_75t_R FILLER_180_847 ();
 DECAPx10_ASAP7_75t_R FILLER_180_869 ();
 DECAPx10_ASAP7_75t_R FILLER_180_891 ();
 DECAPx4_ASAP7_75t_R FILLER_180_913 ();
 DECAPx10_ASAP7_75t_R FILLER_180_935 ();
 DECAPx6_ASAP7_75t_R FILLER_180_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_971 ();
 DECAPx2_ASAP7_75t_R FILLER_180_984 ();
 FILLER_ASAP7_75t_R FILLER_180_990 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1007 ();
 FILLER_ASAP7_75t_R FILLER_180_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1122 ();
 FILLER_ASAP7_75t_R FILLER_180_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1133 ();
 FILLER_ASAP7_75t_R FILLER_180_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1172 ();
 FILLER_ASAP7_75t_R FILLER_180_1182 ();
 FILLER_ASAP7_75t_R FILLER_180_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_181_172 ();
 FILLER_ASAP7_75t_R FILLER_181_186 ();
 DECAPx6_ASAP7_75t_R FILLER_181_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_214 ();
 DECAPx2_ASAP7_75t_R FILLER_181_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_235 ();
 DECAPx6_ASAP7_75t_R FILLER_181_242 ();
 DECAPx1_ASAP7_75t_R FILLER_181_262 ();
 DECAPx6_ASAP7_75t_R FILLER_181_282 ();
 DECAPx1_ASAP7_75t_R FILLER_181_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_308 ();
 DECAPx10_ASAP7_75t_R FILLER_181_324 ();
 DECAPx10_ASAP7_75t_R FILLER_181_346 ();
 DECAPx2_ASAP7_75t_R FILLER_181_368 ();
 FILLER_ASAP7_75t_R FILLER_181_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_376 ();
 DECAPx6_ASAP7_75t_R FILLER_181_408 ();
 DECAPx2_ASAP7_75t_R FILLER_181_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_434 ();
 DECAPx2_ASAP7_75t_R FILLER_181_454 ();
 FILLER_ASAP7_75t_R FILLER_181_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_462 ();
 DECAPx10_ASAP7_75t_R FILLER_181_470 ();
 DECAPx1_ASAP7_75t_R FILLER_181_492 ();
 DECAPx1_ASAP7_75t_R FILLER_181_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_551 ();
 DECAPx2_ASAP7_75t_R FILLER_181_555 ();
 FILLER_ASAP7_75t_R FILLER_181_561 ();
 DECAPx2_ASAP7_75t_R FILLER_181_571 ();
 DECAPx6_ASAP7_75t_R FILLER_181_580 ();
 FILLER_ASAP7_75t_R FILLER_181_594 ();
 DECAPx4_ASAP7_75t_R FILLER_181_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_612 ();
 DECAPx10_ASAP7_75t_R FILLER_181_624 ();
 DECAPx1_ASAP7_75t_R FILLER_181_646 ();
 DECAPx6_ASAP7_75t_R FILLER_181_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_674 ();
 DECAPx10_ASAP7_75t_R FILLER_181_695 ();
 DECAPx10_ASAP7_75t_R FILLER_181_717 ();
 DECAPx10_ASAP7_75t_R FILLER_181_739 ();
 DECAPx6_ASAP7_75t_R FILLER_181_761 ();
 DECAPx1_ASAP7_75t_R FILLER_181_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_779 ();
 DECAPx4_ASAP7_75t_R FILLER_181_794 ();
 FILLER_ASAP7_75t_R FILLER_181_804 ();
 DECAPx10_ASAP7_75t_R FILLER_181_813 ();
 DECAPx10_ASAP7_75t_R FILLER_181_835 ();
 DECAPx6_ASAP7_75t_R FILLER_181_857 ();
 DECAPx2_ASAP7_75t_R FILLER_181_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_877 ();
 DECAPx10_ASAP7_75t_R FILLER_181_892 ();
 FILLER_ASAP7_75t_R FILLER_181_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_916 ();
 DECAPx6_ASAP7_75t_R FILLER_181_943 ();
 DECAPx2_ASAP7_75t_R FILLER_181_957 ();
 DECAPx10_ASAP7_75t_R FILLER_181_975 ();
 DECAPx10_ASAP7_75t_R FILLER_181_997 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1039 ();
 FILLER_ASAP7_75t_R FILLER_181_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1096 ();
 FILLER_ASAP7_75t_R FILLER_181_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1155 ();
 FILLER_ASAP7_75t_R FILLER_181_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1277 ();
 FILLER_ASAP7_75t_R FILLER_181_1291 ();
 DECAPx4_ASAP7_75t_R FILLER_182_172 ();
 DECAPx6_ASAP7_75t_R FILLER_182_194 ();
 DECAPx1_ASAP7_75t_R FILLER_182_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_212 ();
 DECAPx1_ASAP7_75t_R FILLER_182_228 ();
 DECAPx6_ASAP7_75t_R FILLER_182_239 ();
 DECAPx10_ASAP7_75t_R FILLER_182_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_282 ();
 DECAPx2_ASAP7_75t_R FILLER_182_291 ();
 FILLER_ASAP7_75t_R FILLER_182_297 ();
 DECAPx10_ASAP7_75t_R FILLER_182_312 ();
 DECAPx2_ASAP7_75t_R FILLER_182_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_350 ();
 DECAPx10_ASAP7_75t_R FILLER_182_364 ();
 DECAPx10_ASAP7_75t_R FILLER_182_386 ();
 DECAPx6_ASAP7_75t_R FILLER_182_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_422 ();
 FILLER_ASAP7_75t_R FILLER_182_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_443 ();
 DECAPx6_ASAP7_75t_R FILLER_182_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_461 ();
 DECAPx10_ASAP7_75t_R FILLER_182_472 ();
 DECAPx2_ASAP7_75t_R FILLER_182_494 ();
 FILLER_ASAP7_75t_R FILLER_182_500 ();
 DECAPx4_ASAP7_75t_R FILLER_182_523 ();
 FILLER_ASAP7_75t_R FILLER_182_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_535 ();
 FILLER_ASAP7_75t_R FILLER_182_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_559 ();
 DECAPx1_ASAP7_75t_R FILLER_182_581 ();
 DECAPx6_ASAP7_75t_R FILLER_182_593 ();
 FILLER_ASAP7_75t_R FILLER_182_607 ();
 FILLER_ASAP7_75t_R FILLER_182_630 ();
 DECAPx10_ASAP7_75t_R FILLER_182_634 ();
 DECAPx10_ASAP7_75t_R FILLER_182_656 ();
 DECAPx4_ASAP7_75t_R FILLER_182_678 ();
 FILLER_ASAP7_75t_R FILLER_182_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_690 ();
 DECAPx6_ASAP7_75t_R FILLER_182_697 ();
 FILLER_ASAP7_75t_R FILLER_182_711 ();
 DECAPx4_ASAP7_75t_R FILLER_182_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_731 ();
 DECAPx6_ASAP7_75t_R FILLER_182_740 ();
 FILLER_ASAP7_75t_R FILLER_182_754 ();
 FILLER_ASAP7_75t_R FILLER_182_762 ();
 DECAPx10_ASAP7_75t_R FILLER_182_774 ();
 DECAPx10_ASAP7_75t_R FILLER_182_796 ();
 DECAPx10_ASAP7_75t_R FILLER_182_818 ();
 DECAPx10_ASAP7_75t_R FILLER_182_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_862 ();
 DECAPx6_ASAP7_75t_R FILLER_182_869 ();
 DECAPx1_ASAP7_75t_R FILLER_182_883 ();
 DECAPx10_ASAP7_75t_R FILLER_182_893 ();
 DECAPx4_ASAP7_75t_R FILLER_182_915 ();
 FILLER_ASAP7_75t_R FILLER_182_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_942 ();
 DECAPx6_ASAP7_75t_R FILLER_182_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_965 ();
 DECAPx10_ASAP7_75t_R FILLER_182_974 ();
 DECAPx6_ASAP7_75t_R FILLER_182_996 ();
 FILLER_ASAP7_75t_R FILLER_182_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1027 ();
 FILLER_ASAP7_75t_R FILLER_182_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1045 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1157 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1185 ();
 FILLER_ASAP7_75t_R FILLER_182_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1269 ();
 FILLER_ASAP7_75t_R FILLER_182_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_183_172 ();
 FILLER_ASAP7_75t_R FILLER_183_186 ();
 DECAPx2_ASAP7_75t_R FILLER_183_200 ();
 FILLER_ASAP7_75t_R FILLER_183_206 ();
 FILLER_ASAP7_75t_R FILLER_183_214 ();
 DECAPx1_ASAP7_75t_R FILLER_183_224 ();
 DECAPx1_ASAP7_75t_R FILLER_183_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_238 ();
 DECAPx10_ASAP7_75t_R FILLER_183_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_285 ();
 DECAPx2_ASAP7_75t_R FILLER_183_298 ();
 FILLER_ASAP7_75t_R FILLER_183_304 ();
 DECAPx4_ASAP7_75t_R FILLER_183_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_354 ();
 FILLER_ASAP7_75t_R FILLER_183_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_371 ();
 FILLER_ASAP7_75t_R FILLER_183_379 ();
 FILLER_ASAP7_75t_R FILLER_183_392 ();
 FILLER_ASAP7_75t_R FILLER_183_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_403 ();
 DECAPx10_ASAP7_75t_R FILLER_183_410 ();
 DECAPx10_ASAP7_75t_R FILLER_183_432 ();
 DECAPx10_ASAP7_75t_R FILLER_183_454 ();
 DECAPx10_ASAP7_75t_R FILLER_183_476 ();
 DECAPx10_ASAP7_75t_R FILLER_183_498 ();
 DECAPx10_ASAP7_75t_R FILLER_183_520 ();
 DECAPx6_ASAP7_75t_R FILLER_183_542 ();
 FILLER_ASAP7_75t_R FILLER_183_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_558 ();
 DECAPx2_ASAP7_75t_R FILLER_183_565 ();
 FILLER_ASAP7_75t_R FILLER_183_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_573 ();
 FILLER_ASAP7_75t_R FILLER_183_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_598 ();
 DECAPx10_ASAP7_75t_R FILLER_183_602 ();
 DECAPx6_ASAP7_75t_R FILLER_183_624 ();
 DECAPx1_ASAP7_75t_R FILLER_183_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_642 ();
 DECAPx10_ASAP7_75t_R FILLER_183_675 ();
 DECAPx1_ASAP7_75t_R FILLER_183_707 ();
 DECAPx10_ASAP7_75t_R FILLER_183_721 ();
 DECAPx10_ASAP7_75t_R FILLER_183_743 ();
 DECAPx10_ASAP7_75t_R FILLER_183_765 ();
 DECAPx6_ASAP7_75t_R FILLER_183_787 ();
 DECAPx1_ASAP7_75t_R FILLER_183_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_805 ();
 DECAPx1_ASAP7_75t_R FILLER_183_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_818 ();
 DECAPx4_ASAP7_75t_R FILLER_183_822 ();
 DECAPx10_ASAP7_75t_R FILLER_183_840 ();
 DECAPx10_ASAP7_75t_R FILLER_183_862 ();
 DECAPx10_ASAP7_75t_R FILLER_183_884 ();
 DECAPx10_ASAP7_75t_R FILLER_183_906 ();
 DECAPx10_ASAP7_75t_R FILLER_183_928 ();
 FILLER_ASAP7_75t_R FILLER_183_950 ();
 DECAPx4_ASAP7_75t_R FILLER_183_970 ();
 FILLER_ASAP7_75t_R FILLER_183_980 ();
 DECAPx1_ASAP7_75t_R FILLER_183_988 ();
 DECAPx2_ASAP7_75t_R FILLER_183_998 ();
 FILLER_ASAP7_75t_R FILLER_183_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1043 ();
 FILLER_ASAP7_75t_R FILLER_183_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1093 ();
 FILLER_ASAP7_75t_R FILLER_183_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_183_1104 ();
 FILLER_ASAP7_75t_R FILLER_183_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_184_172 ();
 FILLER_ASAP7_75t_R FILLER_184_182 ();
 DECAPx6_ASAP7_75t_R FILLER_184_206 ();
 FILLER_ASAP7_75t_R FILLER_184_228 ();
 DECAPx10_ASAP7_75t_R FILLER_184_242 ();
 DECAPx1_ASAP7_75t_R FILLER_184_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_272 ();
 DECAPx10_ASAP7_75t_R FILLER_184_276 ();
 DECAPx10_ASAP7_75t_R FILLER_184_298 ();
 DECAPx10_ASAP7_75t_R FILLER_184_320 ();
 DECAPx6_ASAP7_75t_R FILLER_184_342 ();
 DECAPx2_ASAP7_75t_R FILLER_184_356 ();
 DECAPx2_ASAP7_75t_R FILLER_184_378 ();
 FILLER_ASAP7_75t_R FILLER_184_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_402 ();
 DECAPx6_ASAP7_75t_R FILLER_184_410 ();
 DECAPx2_ASAP7_75t_R FILLER_184_424 ();
 DECAPx1_ASAP7_75t_R FILLER_184_467 ();
 FILLER_ASAP7_75t_R FILLER_184_483 ();
 DECAPx2_ASAP7_75t_R FILLER_184_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_500 ();
 DECAPx2_ASAP7_75t_R FILLER_184_511 ();
 FILLER_ASAP7_75t_R FILLER_184_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_519 ();
 FILLER_ASAP7_75t_R FILLER_184_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_530 ();
 DECAPx10_ASAP7_75t_R FILLER_184_534 ();
 DECAPx10_ASAP7_75t_R FILLER_184_556 ();
 DECAPx1_ASAP7_75t_R FILLER_184_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_582 ();
 DECAPx10_ASAP7_75t_R FILLER_184_604 ();
 DECAPx2_ASAP7_75t_R FILLER_184_626 ();
 DECAPx2_ASAP7_75t_R FILLER_184_634 ();
 FILLER_ASAP7_75t_R FILLER_184_640 ();
 DECAPx10_ASAP7_75t_R FILLER_184_652 ();
 DECAPx10_ASAP7_75t_R FILLER_184_674 ();
 DECAPx10_ASAP7_75t_R FILLER_184_696 ();
 DECAPx10_ASAP7_75t_R FILLER_184_718 ();
 DECAPx10_ASAP7_75t_R FILLER_184_740 ();
 DECAPx6_ASAP7_75t_R FILLER_184_762 ();
 FILLER_ASAP7_75t_R FILLER_184_776 ();
 DECAPx6_ASAP7_75t_R FILLER_184_786 ();
 FILLER_ASAP7_75t_R FILLER_184_800 ();
 DECAPx10_ASAP7_75t_R FILLER_184_823 ();
 DECAPx10_ASAP7_75t_R FILLER_184_845 ();
 DECAPx10_ASAP7_75t_R FILLER_184_867 ();
 DECAPx10_ASAP7_75t_R FILLER_184_889 ();
 DECAPx10_ASAP7_75t_R FILLER_184_911 ();
 DECAPx10_ASAP7_75t_R FILLER_184_933 ();
 DECAPx10_ASAP7_75t_R FILLER_184_955 ();
 FILLER_ASAP7_75t_R FILLER_184_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_979 ();
 FILLER_ASAP7_75t_R FILLER_184_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_988 ();
 DECAPx10_ASAP7_75t_R FILLER_184_999 ();
 FILLER_ASAP7_75t_R FILLER_184_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1029 ();
 FILLER_ASAP7_75t_R FILLER_184_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1085 ();
 FILLER_ASAP7_75t_R FILLER_184_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1093 ();
 FILLER_ASAP7_75t_R FILLER_184_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1190 ();
 FILLER_ASAP7_75t_R FILLER_184_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_185_172 ();
 DECAPx1_ASAP7_75t_R FILLER_185_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_198 ();
 DECAPx4_ASAP7_75t_R FILLER_185_205 ();
 FILLER_ASAP7_75t_R FILLER_185_221 ();
 DECAPx2_ASAP7_75t_R FILLER_185_229 ();
 DECAPx6_ASAP7_75t_R FILLER_185_245 ();
 FILLER_ASAP7_75t_R FILLER_185_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_261 ();
 DECAPx4_ASAP7_75t_R FILLER_185_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_290 ();
 DECAPx2_ASAP7_75t_R FILLER_185_294 ();
 FILLER_ASAP7_75t_R FILLER_185_300 ();
 DECAPx10_ASAP7_75t_R FILLER_185_349 ();
 DECAPx2_ASAP7_75t_R FILLER_185_379 ();
 DECAPx10_ASAP7_75t_R FILLER_185_405 ();
 DECAPx1_ASAP7_75t_R FILLER_185_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_465 ();
 FILLER_ASAP7_75t_R FILLER_185_473 ();
 FILLER_ASAP7_75t_R FILLER_185_485 ();
 DECAPx1_ASAP7_75t_R FILLER_185_496 ();
 DECAPx1_ASAP7_75t_R FILLER_185_512 ();
 DECAPx1_ASAP7_75t_R FILLER_185_537 ();
 DECAPx1_ASAP7_75t_R FILLER_185_549 ();
 DECAPx2_ASAP7_75t_R FILLER_185_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_571 ();
 DECAPx10_ASAP7_75t_R FILLER_185_575 ();
 DECAPx1_ASAP7_75t_R FILLER_185_597 ();
 DECAPx6_ASAP7_75t_R FILLER_185_622 ();
 DECAPx2_ASAP7_75t_R FILLER_185_636 ();
 DECAPx10_ASAP7_75t_R FILLER_185_652 ();
 DECAPx4_ASAP7_75t_R FILLER_185_674 ();
 FILLER_ASAP7_75t_R FILLER_185_684 ();
 DECAPx6_ASAP7_75t_R FILLER_185_692 ();
 FILLER_ASAP7_75t_R FILLER_185_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_708 ();
 DECAPx10_ASAP7_75t_R FILLER_185_721 ();
 DECAPx10_ASAP7_75t_R FILLER_185_743 ();
 DECAPx10_ASAP7_75t_R FILLER_185_765 ();
 DECAPx10_ASAP7_75t_R FILLER_185_787 ();
 DECAPx10_ASAP7_75t_R FILLER_185_809 ();
 DECAPx10_ASAP7_75t_R FILLER_185_831 ();
 DECAPx10_ASAP7_75t_R FILLER_185_853 ();
 DECAPx4_ASAP7_75t_R FILLER_185_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_885 ();
 DECAPx10_ASAP7_75t_R FILLER_185_897 ();
 DECAPx4_ASAP7_75t_R FILLER_185_919 ();
 FILLER_ASAP7_75t_R FILLER_185_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_931 ();
 DECAPx10_ASAP7_75t_R FILLER_185_942 ();
 DECAPx10_ASAP7_75t_R FILLER_185_964 ();
 DECAPx10_ASAP7_75t_R FILLER_185_986 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1008 ();
 FILLER_ASAP7_75t_R FILLER_185_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1082 ();
 FILLER_ASAP7_75t_R FILLER_185_1092 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1096 ();
 FILLER_ASAP7_75t_R FILLER_185_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1170 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1192 ();
 FILLER_ASAP7_75t_R FILLER_185_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1269 ();
 FILLER_ASAP7_75t_R FILLER_185_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_186_172 ();
 FILLER_ASAP7_75t_R FILLER_186_186 ();
 DECAPx4_ASAP7_75t_R FILLER_186_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_212 ();
 DECAPx10_ASAP7_75t_R FILLER_186_216 ();
 DECAPx6_ASAP7_75t_R FILLER_186_238 ();
 DECAPx2_ASAP7_75t_R FILLER_186_252 ();
 FILLER_ASAP7_75t_R FILLER_186_265 ();
 DECAPx2_ASAP7_75t_R FILLER_186_270 ();
 DECAPx2_ASAP7_75t_R FILLER_186_285 ();
 FILLER_ASAP7_75t_R FILLER_186_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_293 ();
 DECAPx10_ASAP7_75t_R FILLER_186_303 ();
 DECAPx2_ASAP7_75t_R FILLER_186_325 ();
 DECAPx10_ASAP7_75t_R FILLER_186_338 ();
 DECAPx10_ASAP7_75t_R FILLER_186_360 ();
 DECAPx6_ASAP7_75t_R FILLER_186_382 ();
 DECAPx1_ASAP7_75t_R FILLER_186_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_400 ();
 DECAPx6_ASAP7_75t_R FILLER_186_407 ();
 DECAPx2_ASAP7_75t_R FILLER_186_421 ();
 DECAPx10_ASAP7_75t_R FILLER_186_449 ();
 DECAPx1_ASAP7_75t_R FILLER_186_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_475 ();
 DECAPx10_ASAP7_75t_R FILLER_186_485 ();
 DECAPx4_ASAP7_75t_R FILLER_186_507 ();
 DECAPx4_ASAP7_75t_R FILLER_186_523 ();
 FILLER_ASAP7_75t_R FILLER_186_533 ();
 FILLER_ASAP7_75t_R FILLER_186_556 ();
 DECAPx2_ASAP7_75t_R FILLER_186_579 ();
 FILLER_ASAP7_75t_R FILLER_186_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_604 ();
 FILLER_ASAP7_75t_R FILLER_186_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_615 ();
 DECAPx4_ASAP7_75t_R FILLER_186_619 ();
 FILLER_ASAP7_75t_R FILLER_186_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_631 ();
 DECAPx4_ASAP7_75t_R FILLER_186_634 ();
 DECAPx10_ASAP7_75t_R FILLER_186_662 ();
 DECAPx1_ASAP7_75t_R FILLER_186_684 ();
 DECAPx10_ASAP7_75t_R FILLER_186_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_716 ();
 DECAPx10_ASAP7_75t_R FILLER_186_723 ();
 DECAPx6_ASAP7_75t_R FILLER_186_745 ();
 FILLER_ASAP7_75t_R FILLER_186_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_761 ();
 DECAPx10_ASAP7_75t_R FILLER_186_772 ();
 DECAPx10_ASAP7_75t_R FILLER_186_794 ();
 DECAPx10_ASAP7_75t_R FILLER_186_816 ();
 DECAPx10_ASAP7_75t_R FILLER_186_838 ();
 DECAPx10_ASAP7_75t_R FILLER_186_860 ();
 DECAPx1_ASAP7_75t_R FILLER_186_882 ();
 DECAPx10_ASAP7_75t_R FILLER_186_892 ();
 DECAPx1_ASAP7_75t_R FILLER_186_914 ();
 DECAPx10_ASAP7_75t_R FILLER_186_938 ();
 FILLER_ASAP7_75t_R FILLER_186_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_962 ();
 DECAPx1_ASAP7_75t_R FILLER_186_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_973 ();
 DECAPx6_ASAP7_75t_R FILLER_186_980 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1000 ();
 FILLER_ASAP7_75t_R FILLER_186_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1016 ();
 FILLER_ASAP7_75t_R FILLER_186_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1063 ();
 FILLER_ASAP7_75t_R FILLER_186_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_187_172 ();
 FILLER_ASAP7_75t_R FILLER_187_178 ();
 DECAPx4_ASAP7_75t_R FILLER_187_204 ();
 FILLER_ASAP7_75t_R FILLER_187_214 ();
 FILLER_ASAP7_75t_R FILLER_187_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_224 ();
 DECAPx6_ASAP7_75t_R FILLER_187_235 ();
 DECAPx2_ASAP7_75t_R FILLER_187_249 ();
 DECAPx1_ASAP7_75t_R FILLER_187_277 ();
 DECAPx2_ASAP7_75t_R FILLER_187_284 ();
 DECAPx10_ASAP7_75t_R FILLER_187_299 ();
 DECAPx6_ASAP7_75t_R FILLER_187_321 ();
 DECAPx4_ASAP7_75t_R FILLER_187_342 ();
 FILLER_ASAP7_75t_R FILLER_187_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_354 ();
 DECAPx1_ASAP7_75t_R FILLER_187_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_382 ();
 DECAPx6_ASAP7_75t_R FILLER_187_389 ();
 FILLER_ASAP7_75t_R FILLER_187_403 ();
 DECAPx6_ASAP7_75t_R FILLER_187_415 ();
 FILLER_ASAP7_75t_R FILLER_187_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_431 ();
 DECAPx10_ASAP7_75t_R FILLER_187_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_464 ();
 DECAPx10_ASAP7_75t_R FILLER_187_474 ();
 DECAPx10_ASAP7_75t_R FILLER_187_496 ();
 DECAPx6_ASAP7_75t_R FILLER_187_518 ();
 DECAPx2_ASAP7_75t_R FILLER_187_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_538 ();
 DECAPx1_ASAP7_75t_R FILLER_187_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_557 ();
 DECAPx6_ASAP7_75t_R FILLER_187_564 ();
 DECAPx1_ASAP7_75t_R FILLER_187_599 ();
 FILLER_ASAP7_75t_R FILLER_187_609 ();
 DECAPx6_ASAP7_75t_R FILLER_187_619 ();
 DECAPx10_ASAP7_75t_R FILLER_187_636 ();
 DECAPx6_ASAP7_75t_R FILLER_187_658 ();
 DECAPx1_ASAP7_75t_R FILLER_187_672 ();
 DECAPx2_ASAP7_75t_R FILLER_187_682 ();
 FILLER_ASAP7_75t_R FILLER_187_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_690 ();
 FILLER_ASAP7_75t_R FILLER_187_697 ();
 DECAPx2_ASAP7_75t_R FILLER_187_711 ();
 FILLER_ASAP7_75t_R FILLER_187_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_719 ();
 DECAPx2_ASAP7_75t_R FILLER_187_726 ();
 DECAPx10_ASAP7_75t_R FILLER_187_746 ();
 DECAPx10_ASAP7_75t_R FILLER_187_768 ();
 DECAPx2_ASAP7_75t_R FILLER_187_790 ();
 DECAPx10_ASAP7_75t_R FILLER_187_802 ();
 DECAPx2_ASAP7_75t_R FILLER_187_824 ();
 DECAPx4_ASAP7_75t_R FILLER_187_836 ();
 DECAPx2_ASAP7_75t_R FILLER_187_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_869 ();
 DECAPx10_ASAP7_75t_R FILLER_187_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_908 ();
 DECAPx10_ASAP7_75t_R FILLER_187_919 ();
 DECAPx6_ASAP7_75t_R FILLER_187_941 ();
 FILLER_ASAP7_75t_R FILLER_187_955 ();
 DECAPx4_ASAP7_75t_R FILLER_187_984 ();
 FILLER_ASAP7_75t_R FILLER_187_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_996 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1014 ();
 FILLER_ASAP7_75t_R FILLER_187_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1042 ();
 FILLER_ASAP7_75t_R FILLER_187_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_188_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_186 ();
 DECAPx2_ASAP7_75t_R FILLER_188_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_212 ();
 FILLER_ASAP7_75t_R FILLER_188_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_244 ();
 DECAPx10_ASAP7_75t_R FILLER_188_257 ();
 DECAPx4_ASAP7_75t_R FILLER_188_279 ();
 DECAPx4_ASAP7_75t_R FILLER_188_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_311 ();
 FILLER_ASAP7_75t_R FILLER_188_318 ();
 DECAPx1_ASAP7_75t_R FILLER_188_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_344 ();
 DECAPx4_ASAP7_75t_R FILLER_188_373 ();
 DECAPx10_ASAP7_75t_R FILLER_188_391 ();
 DECAPx4_ASAP7_75t_R FILLER_188_413 ();
 FILLER_ASAP7_75t_R FILLER_188_423 ();
 DECAPx4_ASAP7_75t_R FILLER_188_447 ();
 FILLER_ASAP7_75t_R FILLER_188_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_459 ();
 DECAPx2_ASAP7_75t_R FILLER_188_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_499 ();
 DECAPx1_ASAP7_75t_R FILLER_188_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_520 ();
 DECAPx6_ASAP7_75t_R FILLER_188_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_538 ();
 DECAPx4_ASAP7_75t_R FILLER_188_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_579 ();
 DECAPx6_ASAP7_75t_R FILLER_188_586 ();
 DECAPx2_ASAP7_75t_R FILLER_188_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_606 ();
 DECAPx1_ASAP7_75t_R FILLER_188_628 ();
 DECAPx4_ASAP7_75t_R FILLER_188_634 ();
 DECAPx6_ASAP7_75t_R FILLER_188_678 ();
 DECAPx1_ASAP7_75t_R FILLER_188_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_696 ();
 DECAPx10_ASAP7_75t_R FILLER_188_700 ();
 DECAPx10_ASAP7_75t_R FILLER_188_722 ();
 DECAPx10_ASAP7_75t_R FILLER_188_744 ();
 DECAPx4_ASAP7_75t_R FILLER_188_766 ();
 FILLER_ASAP7_75t_R FILLER_188_776 ();
 DECAPx2_ASAP7_75t_R FILLER_188_785 ();
 DECAPx1_ASAP7_75t_R FILLER_188_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_801 ();
 DECAPx6_ASAP7_75t_R FILLER_188_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_828 ();
 DECAPx6_ASAP7_75t_R FILLER_188_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_849 ();
 DECAPx10_ASAP7_75t_R FILLER_188_856 ();
 DECAPx4_ASAP7_75t_R FILLER_188_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_888 ();
 DECAPx10_ASAP7_75t_R FILLER_188_913 ();
 DECAPx4_ASAP7_75t_R FILLER_188_935 ();
 DECAPx10_ASAP7_75t_R FILLER_188_952 ();
 DECAPx6_ASAP7_75t_R FILLER_188_974 ();
 FILLER_ASAP7_75t_R FILLER_188_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_990 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1169 ();
 FILLER_ASAP7_75t_R FILLER_188_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_189_172 ();
 DECAPx4_ASAP7_75t_R FILLER_189_200 ();
 FILLER_ASAP7_75t_R FILLER_189_210 ();
 DECAPx4_ASAP7_75t_R FILLER_189_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_229 ();
 DECAPx6_ASAP7_75t_R FILLER_189_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_267 ();
 FILLER_ASAP7_75t_R FILLER_189_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_280 ();
 DECAPx6_ASAP7_75t_R FILLER_189_302 ();
 FILLER_ASAP7_75t_R FILLER_189_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_318 ();
 DECAPx10_ASAP7_75t_R FILLER_189_335 ();
 DECAPx6_ASAP7_75t_R FILLER_189_369 ();
 DECAPx1_ASAP7_75t_R FILLER_189_383 ();
 DECAPx10_ASAP7_75t_R FILLER_189_401 ();
 DECAPx2_ASAP7_75t_R FILLER_189_423 ();
 DECAPx4_ASAP7_75t_R FILLER_189_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_459 ();
 DECAPx4_ASAP7_75t_R FILLER_189_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_478 ();
 FILLER_ASAP7_75t_R FILLER_189_493 ();
 DECAPx2_ASAP7_75t_R FILLER_189_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_507 ();
 DECAPx4_ASAP7_75t_R FILLER_189_529 ();
 DECAPx1_ASAP7_75t_R FILLER_189_570 ();
 FILLER_ASAP7_75t_R FILLER_189_577 ();
 DECAPx1_ASAP7_75t_R FILLER_189_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_590 ();
 DECAPx10_ASAP7_75t_R FILLER_189_621 ();
 DECAPx6_ASAP7_75t_R FILLER_189_643 ();
 DECAPx1_ASAP7_75t_R FILLER_189_657 ();
 DECAPx10_ASAP7_75t_R FILLER_189_667 ();
 FILLER_ASAP7_75t_R FILLER_189_689 ();
 DECAPx6_ASAP7_75t_R FILLER_189_712 ();
 DECAPx2_ASAP7_75t_R FILLER_189_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_732 ();
 DECAPx6_ASAP7_75t_R FILLER_189_741 ();
 FILLER_ASAP7_75t_R FILLER_189_755 ();
 DECAPx10_ASAP7_75t_R FILLER_189_763 ();
 DECAPx10_ASAP7_75t_R FILLER_189_785 ();
 DECAPx10_ASAP7_75t_R FILLER_189_807 ();
 DECAPx10_ASAP7_75t_R FILLER_189_829 ();
 DECAPx10_ASAP7_75t_R FILLER_189_851 ();
 DECAPx6_ASAP7_75t_R FILLER_189_873 ();
 DECAPx1_ASAP7_75t_R FILLER_189_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_891 ();
 DECAPx2_ASAP7_75t_R FILLER_189_900 ();
 DECAPx10_ASAP7_75t_R FILLER_189_912 ();
 FILLER_ASAP7_75t_R FILLER_189_941 ();
 DECAPx10_ASAP7_75t_R FILLER_189_949 ();
 FILLER_ASAP7_75t_R FILLER_189_971 ();
 DECAPx4_ASAP7_75t_R FILLER_189_979 ();
 DECAPx10_ASAP7_75t_R FILLER_189_997 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_189_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1100 ();
 FILLER_ASAP7_75t_R FILLER_189_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_189_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_189_1180 ();
 FILLER_ASAP7_75t_R FILLER_189_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_190_172 ();
 FILLER_ASAP7_75t_R FILLER_190_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_184 ();
 DECAPx10_ASAP7_75t_R FILLER_190_197 ();
 DECAPx6_ASAP7_75t_R FILLER_190_219 ();
 FILLER_ASAP7_75t_R FILLER_190_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_235 ();
 FILLER_ASAP7_75t_R FILLER_190_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_249 ();
 FILLER_ASAP7_75t_R FILLER_190_271 ();
 DECAPx1_ASAP7_75t_R FILLER_190_279 ();
 DECAPx1_ASAP7_75t_R FILLER_190_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_295 ();
 DECAPx1_ASAP7_75t_R FILLER_190_302 ();
 DECAPx6_ASAP7_75t_R FILLER_190_319 ();
 DECAPx2_ASAP7_75t_R FILLER_190_333 ();
 DECAPx6_ASAP7_75t_R FILLER_190_344 ();
 FILLER_ASAP7_75t_R FILLER_190_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_360 ();
 DECAPx10_ASAP7_75t_R FILLER_190_385 ();
 DECAPx10_ASAP7_75t_R FILLER_190_407 ();
 DECAPx10_ASAP7_75t_R FILLER_190_429 ();
 DECAPx6_ASAP7_75t_R FILLER_190_451 ();
 DECAPx2_ASAP7_75t_R FILLER_190_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_471 ();
 DECAPx2_ASAP7_75t_R FILLER_190_500 ();
 FILLER_ASAP7_75t_R FILLER_190_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_508 ();
 DECAPx6_ASAP7_75t_R FILLER_190_515 ();
 DECAPx2_ASAP7_75t_R FILLER_190_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_535 ();
 DECAPx1_ASAP7_75t_R FILLER_190_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_582 ();
 FILLER_ASAP7_75t_R FILLER_190_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_623 ();
 DECAPx10_ASAP7_75t_R FILLER_190_634 ();
 DECAPx1_ASAP7_75t_R FILLER_190_656 ();
 DECAPx2_ASAP7_75t_R FILLER_190_666 ();
 FILLER_ASAP7_75t_R FILLER_190_672 ();
 DECAPx10_ASAP7_75t_R FILLER_190_680 ();
 DECAPx10_ASAP7_75t_R FILLER_190_702 ();
 DECAPx2_ASAP7_75t_R FILLER_190_724 ();
 FILLER_ASAP7_75t_R FILLER_190_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_732 ();
 DECAPx10_ASAP7_75t_R FILLER_190_739 ();
 DECAPx10_ASAP7_75t_R FILLER_190_761 ();
 DECAPx10_ASAP7_75t_R FILLER_190_783 ();
 DECAPx10_ASAP7_75t_R FILLER_190_805 ();
 DECAPx10_ASAP7_75t_R FILLER_190_827 ();
 DECAPx2_ASAP7_75t_R FILLER_190_849 ();
 FILLER_ASAP7_75t_R FILLER_190_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_857 ();
 DECAPx2_ASAP7_75t_R FILLER_190_882 ();
 DECAPx4_ASAP7_75t_R FILLER_190_895 ();
 FILLER_ASAP7_75t_R FILLER_190_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_907 ();
 DECAPx1_ASAP7_75t_R FILLER_190_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_919 ();
 FILLER_ASAP7_75t_R FILLER_190_933 ();
 DECAPx10_ASAP7_75t_R FILLER_190_941 ();
 DECAPx4_ASAP7_75t_R FILLER_190_963 ();
 FILLER_ASAP7_75t_R FILLER_190_973 ();
 DECAPx2_ASAP7_75t_R FILLER_190_981 ();
 FILLER_ASAP7_75t_R FILLER_190_987 ();
 DECAPx6_ASAP7_75t_R FILLER_190_997 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1121 ();
 FILLER_ASAP7_75t_R FILLER_190_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1157 ();
 FILLER_ASAP7_75t_R FILLER_190_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1191 ();
 FILLER_ASAP7_75t_R FILLER_190_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_191_172 ();
 FILLER_ASAP7_75t_R FILLER_191_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_180 ();
 DECAPx10_ASAP7_75t_R FILLER_191_195 ();
 DECAPx6_ASAP7_75t_R FILLER_191_217 ();
 DECAPx2_ASAP7_75t_R FILLER_191_231 ();
 DECAPx6_ASAP7_75t_R FILLER_191_245 ();
 DECAPx2_ASAP7_75t_R FILLER_191_259 ();
 DECAPx10_ASAP7_75t_R FILLER_191_271 ();
 DECAPx4_ASAP7_75t_R FILLER_191_293 ();
 FILLER_ASAP7_75t_R FILLER_191_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_305 ();
 DECAPx2_ASAP7_75t_R FILLER_191_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_326 ();
 DECAPx4_ASAP7_75t_R FILLER_191_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_368 ();
 DECAPx10_ASAP7_75t_R FILLER_191_375 ();
 FILLER_ASAP7_75t_R FILLER_191_397 ();
 DECAPx10_ASAP7_75t_R FILLER_191_409 ();
 DECAPx10_ASAP7_75t_R FILLER_191_431 ();
 DECAPx2_ASAP7_75t_R FILLER_191_453 ();
 FILLER_ASAP7_75t_R FILLER_191_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_461 ();
 DECAPx6_ASAP7_75t_R FILLER_191_490 ();
 DECAPx1_ASAP7_75t_R FILLER_191_504 ();
 DECAPx4_ASAP7_75t_R FILLER_191_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_526 ();
 DECAPx2_ASAP7_75t_R FILLER_191_530 ();
 FILLER_ASAP7_75t_R FILLER_191_536 ();
 DECAPx10_ASAP7_75t_R FILLER_191_549 ();
 DECAPx4_ASAP7_75t_R FILLER_191_571 ();
 FILLER_ASAP7_75t_R FILLER_191_581 ();
 DECAPx2_ASAP7_75t_R FILLER_191_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_610 ();
 FILLER_ASAP7_75t_R FILLER_191_614 ();
 DECAPx2_ASAP7_75t_R FILLER_191_630 ();
 FILLER_ASAP7_75t_R FILLER_191_636 ();
 DECAPx10_ASAP7_75t_R FILLER_191_656 ();
 DECAPx10_ASAP7_75t_R FILLER_191_678 ();
 FILLER_ASAP7_75t_R FILLER_191_700 ();
 DECAPx6_ASAP7_75t_R FILLER_191_720 ();
 DECAPx1_ASAP7_75t_R FILLER_191_734 ();
 DECAPx10_ASAP7_75t_R FILLER_191_748 ();
 FILLER_ASAP7_75t_R FILLER_191_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_772 ();
 DECAPx10_ASAP7_75t_R FILLER_191_781 ();
 DECAPx10_ASAP7_75t_R FILLER_191_803 ();
 DECAPx1_ASAP7_75t_R FILLER_191_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_829 ();
 FILLER_ASAP7_75t_R FILLER_191_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_838 ();
 DECAPx4_ASAP7_75t_R FILLER_191_857 ();
 DECAPx10_ASAP7_75t_R FILLER_191_875 ();
 DECAPx10_ASAP7_75t_R FILLER_191_897 ();
 DECAPx10_ASAP7_75t_R FILLER_191_919 ();
 DECAPx6_ASAP7_75t_R FILLER_191_941 ();
 DECAPx2_ASAP7_75t_R FILLER_191_955 ();
 DECAPx10_ASAP7_75t_R FILLER_191_977 ();
 DECAPx2_ASAP7_75t_R FILLER_191_999 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1013 ();
 DECAPx4_ASAP7_75t_R FILLER_191_1035 ();
 FILLER_ASAP7_75t_R FILLER_191_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1053 ();
 FILLER_ASAP7_75t_R FILLER_191_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_191_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_192_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_182 ();
 DECAPx2_ASAP7_75t_R FILLER_192_203 ();
 DECAPx4_ASAP7_75t_R FILLER_192_216 ();
 DECAPx2_ASAP7_75t_R FILLER_192_240 ();
 DECAPx10_ASAP7_75t_R FILLER_192_257 ();
 DECAPx1_ASAP7_75t_R FILLER_192_279 ();
 DECAPx2_ASAP7_75t_R FILLER_192_304 ();
 DECAPx6_ASAP7_75t_R FILLER_192_316 ();
 DECAPx2_ASAP7_75t_R FILLER_192_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_336 ();
 DECAPx10_ASAP7_75t_R FILLER_192_340 ();
 DECAPx4_ASAP7_75t_R FILLER_192_362 ();
 FILLER_ASAP7_75t_R FILLER_192_372 ();
 FILLER_ASAP7_75t_R FILLER_192_380 ();
 FILLER_ASAP7_75t_R FILLER_192_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_392 ();
 DECAPx2_ASAP7_75t_R FILLER_192_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_405 ();
 DECAPx4_ASAP7_75t_R FILLER_192_412 ();
 FILLER_ASAP7_75t_R FILLER_192_422 ();
 DECAPx4_ASAP7_75t_R FILLER_192_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_452 ();
 DECAPx2_ASAP7_75t_R FILLER_192_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_479 ();
 DECAPx1_ASAP7_75t_R FILLER_192_487 ();
 DECAPx2_ASAP7_75t_R FILLER_192_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_512 ();
 FILLER_ASAP7_75t_R FILLER_192_549 ();
 DECAPx10_ASAP7_75t_R FILLER_192_557 ();
 DECAPx4_ASAP7_75t_R FILLER_192_579 ();
 FILLER_ASAP7_75t_R FILLER_192_589 ();
 DECAPx2_ASAP7_75t_R FILLER_192_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_611 ();
 DECAPx1_ASAP7_75t_R FILLER_192_620 ();
 DECAPx10_ASAP7_75t_R FILLER_192_634 ();
 DECAPx10_ASAP7_75t_R FILLER_192_656 ();
 DECAPx10_ASAP7_75t_R FILLER_192_678 ();
 DECAPx10_ASAP7_75t_R FILLER_192_700 ();
 DECAPx10_ASAP7_75t_R FILLER_192_722 ();
 DECAPx10_ASAP7_75t_R FILLER_192_744 ();
 DECAPx10_ASAP7_75t_R FILLER_192_766 ();
 DECAPx10_ASAP7_75t_R FILLER_192_788 ();
 DECAPx10_ASAP7_75t_R FILLER_192_810 ();
 DECAPx10_ASAP7_75t_R FILLER_192_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_854 ();
 DECAPx10_ASAP7_75t_R FILLER_192_861 ();
 DECAPx10_ASAP7_75t_R FILLER_192_883 ();
 DECAPx10_ASAP7_75t_R FILLER_192_905 ();
 DECAPx10_ASAP7_75t_R FILLER_192_927 ();
 DECAPx10_ASAP7_75t_R FILLER_192_949 ();
 DECAPx10_ASAP7_75t_R FILLER_192_971 ();
 FILLER_ASAP7_75t_R FILLER_192_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1002 ();
 FILLER_ASAP7_75t_R FILLER_192_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_193_172 ();
 DECAPx1_ASAP7_75t_R FILLER_193_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_196 ();
 DECAPx4_ASAP7_75t_R FILLER_193_203 ();
 FILLER_ASAP7_75t_R FILLER_193_213 ();
 FILLER_ASAP7_75t_R FILLER_193_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_254 ();
 DECAPx1_ASAP7_75t_R FILLER_193_261 ();
 FILLER_ASAP7_75t_R FILLER_193_272 ();
 DECAPx4_ASAP7_75t_R FILLER_193_282 ();
 DECAPx10_ASAP7_75t_R FILLER_193_307 ();
 DECAPx2_ASAP7_75t_R FILLER_193_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_335 ();
 FILLER_ASAP7_75t_R FILLER_193_345 ();
 FILLER_ASAP7_75t_R FILLER_193_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_381 ();
 DECAPx4_ASAP7_75t_R FILLER_193_388 ();
 FILLER_ASAP7_75t_R FILLER_193_398 ();
 DECAPx4_ASAP7_75t_R FILLER_193_406 ();
 FILLER_ASAP7_75t_R FILLER_193_422 ();
 DECAPx4_ASAP7_75t_R FILLER_193_446 ();
 FILLER_ASAP7_75t_R FILLER_193_456 ();
 DECAPx2_ASAP7_75t_R FILLER_193_474 ();
 DECAPx1_ASAP7_75t_R FILLER_193_486 ();
 DECAPx2_ASAP7_75t_R FILLER_193_568 ();
 DECAPx2_ASAP7_75t_R FILLER_193_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_591 ();
 DECAPx4_ASAP7_75t_R FILLER_193_622 ();
 DECAPx10_ASAP7_75t_R FILLER_193_644 ();
 DECAPx2_ASAP7_75t_R FILLER_193_666 ();
 FILLER_ASAP7_75t_R FILLER_193_678 ();
 DECAPx10_ASAP7_75t_R FILLER_193_686 ();
 DECAPx10_ASAP7_75t_R FILLER_193_708 ();
 DECAPx10_ASAP7_75t_R FILLER_193_730 ();
 DECAPx10_ASAP7_75t_R FILLER_193_752 ();
 DECAPx10_ASAP7_75t_R FILLER_193_774 ();
 FILLER_ASAP7_75t_R FILLER_193_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_808 ();
 DECAPx10_ASAP7_75t_R FILLER_193_815 ();
 DECAPx10_ASAP7_75t_R FILLER_193_837 ();
 DECAPx4_ASAP7_75t_R FILLER_193_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_869 ();
 DECAPx10_ASAP7_75t_R FILLER_193_876 ();
 DECAPx10_ASAP7_75t_R FILLER_193_898 ();
 DECAPx4_ASAP7_75t_R FILLER_193_920 ();
 FILLER_ASAP7_75t_R FILLER_193_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_944 ();
 DECAPx10_ASAP7_75t_R FILLER_193_955 ();
 DECAPx2_ASAP7_75t_R FILLER_193_977 ();
 FILLER_ASAP7_75t_R FILLER_193_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_985 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1002 ();
 FILLER_ASAP7_75t_R FILLER_193_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_193_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1110 ();
 FILLER_ASAP7_75t_R FILLER_193_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_194_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_182 ();
 DECAPx4_ASAP7_75t_R FILLER_194_202 ();
 FILLER_ASAP7_75t_R FILLER_194_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_214 ();
 DECAPx1_ASAP7_75t_R FILLER_194_227 ();
 DECAPx10_ASAP7_75t_R FILLER_194_247 ();
 DECAPx4_ASAP7_75t_R FILLER_194_269 ();
 FILLER_ASAP7_75t_R FILLER_194_279 ();
 DECAPx10_ASAP7_75t_R FILLER_194_312 ();
 DECAPx10_ASAP7_75t_R FILLER_194_334 ();
 DECAPx6_ASAP7_75t_R FILLER_194_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_370 ();
 FILLER_ASAP7_75t_R FILLER_194_383 ();
 DECAPx1_ASAP7_75t_R FILLER_194_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_397 ();
 DECAPx6_ASAP7_75t_R FILLER_194_404 ();
 FILLER_ASAP7_75t_R FILLER_194_418 ();
 FILLER_ASAP7_75t_R FILLER_194_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_434 ();
 DECAPx6_ASAP7_75t_R FILLER_194_442 ();
 DECAPx2_ASAP7_75t_R FILLER_194_456 ();
 DECAPx6_ASAP7_75t_R FILLER_194_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_500 ();
 FILLER_ASAP7_75t_R FILLER_194_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_510 ();
 FILLER_ASAP7_75t_R FILLER_194_567 ();
 DECAPx10_ASAP7_75t_R FILLER_194_590 ();
 DECAPx6_ASAP7_75t_R FILLER_194_612 ();
 DECAPx2_ASAP7_75t_R FILLER_194_626 ();
 DECAPx6_ASAP7_75t_R FILLER_194_634 ();
 FILLER_ASAP7_75t_R FILLER_194_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_650 ();
 DECAPx2_ASAP7_75t_R FILLER_194_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_681 ();
 DECAPx2_ASAP7_75t_R FILLER_194_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_711 ();
 DECAPx10_ASAP7_75t_R FILLER_194_731 ();
 DECAPx10_ASAP7_75t_R FILLER_194_753 ();
 DECAPx10_ASAP7_75t_R FILLER_194_775 ();
 DECAPx10_ASAP7_75t_R FILLER_194_797 ();
 DECAPx10_ASAP7_75t_R FILLER_194_819 ();
 DECAPx10_ASAP7_75t_R FILLER_194_841 ();
 DECAPx6_ASAP7_75t_R FILLER_194_863 ();
 DECAPx1_ASAP7_75t_R FILLER_194_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_881 ();
 DECAPx6_ASAP7_75t_R FILLER_194_888 ();
 DECAPx2_ASAP7_75t_R FILLER_194_902 ();
 DECAPx2_ASAP7_75t_R FILLER_194_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_924 ();
 DECAPx6_ASAP7_75t_R FILLER_194_931 ();
 DECAPx2_ASAP7_75t_R FILLER_194_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_972 ();
 DECAPx10_ASAP7_75t_R FILLER_194_979 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1039 ();
 FILLER_ASAP7_75t_R FILLER_194_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1093 ();
 FILLER_ASAP7_75t_R FILLER_194_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1139 ();
 FILLER_ASAP7_75t_R FILLER_194_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1172 ();
 FILLER_ASAP7_75t_R FILLER_194_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_194_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_195_172 ();
 FILLER_ASAP7_75t_R FILLER_195_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_187 ();
 DECAPx10_ASAP7_75t_R FILLER_195_191 ();
 DECAPx6_ASAP7_75t_R FILLER_195_213 ();
 FILLER_ASAP7_75t_R FILLER_195_227 ();
 DECAPx10_ASAP7_75t_R FILLER_195_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_265 ();
 DECAPx2_ASAP7_75t_R FILLER_195_272 ();
 FILLER_ASAP7_75t_R FILLER_195_278 ();
 DECAPx2_ASAP7_75t_R FILLER_195_288 ();
 FILLER_ASAP7_75t_R FILLER_195_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_316 ();
 DECAPx10_ASAP7_75t_R FILLER_195_348 ();
 DECAPx10_ASAP7_75t_R FILLER_195_370 ();
 DECAPx1_ASAP7_75t_R FILLER_195_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_396 ();
 FILLER_ASAP7_75t_R FILLER_195_407 ();
 DECAPx6_ASAP7_75t_R FILLER_195_419 ();
 DECAPx2_ASAP7_75t_R FILLER_195_433 ();
 FILLER_ASAP7_75t_R FILLER_195_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_453 ();
 DECAPx10_ASAP7_75t_R FILLER_195_471 ();
 DECAPx10_ASAP7_75t_R FILLER_195_493 ();
 DECAPx4_ASAP7_75t_R FILLER_195_515 ();
 FILLER_ASAP7_75t_R FILLER_195_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_527 ();
 DECAPx2_ASAP7_75t_R FILLER_195_538 ();
 DECAPx6_ASAP7_75t_R FILLER_195_552 ();
 DECAPx1_ASAP7_75t_R FILLER_195_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_570 ();
 FILLER_ASAP7_75t_R FILLER_195_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_587 ();
 DECAPx6_ASAP7_75t_R FILLER_195_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_608 ();
 DECAPx6_ASAP7_75t_R FILLER_195_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_631 ();
 DECAPx10_ASAP7_75t_R FILLER_195_661 ();
 DECAPx4_ASAP7_75t_R FILLER_195_683 ();
 FILLER_ASAP7_75t_R FILLER_195_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_695 ();
 DECAPx10_ASAP7_75t_R FILLER_195_723 ();
 DECAPx4_ASAP7_75t_R FILLER_195_745 ();
 DECAPx10_ASAP7_75t_R FILLER_195_763 ();
 FILLER_ASAP7_75t_R FILLER_195_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_787 ();
 DECAPx10_ASAP7_75t_R FILLER_195_799 ();
 DECAPx2_ASAP7_75t_R FILLER_195_821 ();
 FILLER_ASAP7_75t_R FILLER_195_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_829 ();
 DECAPx10_ASAP7_75t_R FILLER_195_838 ();
 DECAPx10_ASAP7_75t_R FILLER_195_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_882 ();
 DECAPx6_ASAP7_75t_R FILLER_195_889 ();
 FILLER_ASAP7_75t_R FILLER_195_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_905 ();
 DECAPx2_ASAP7_75t_R FILLER_195_922 ();
 DECAPx6_ASAP7_75t_R FILLER_195_934 ();
 FILLER_ASAP7_75t_R FILLER_195_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_950 ();
 DECAPx10_ASAP7_75t_R FILLER_195_957 ();
 DECAPx10_ASAP7_75t_R FILLER_195_979 ();
 FILLER_ASAP7_75t_R FILLER_195_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_196_172 ();
 FILLER_ASAP7_75t_R FILLER_196_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_226 ();
 FILLER_ASAP7_75t_R FILLER_196_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_235 ();
 DECAPx6_ASAP7_75t_R FILLER_196_242 ();
 DECAPx1_ASAP7_75t_R FILLER_196_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_274 ();
 DECAPx1_ASAP7_75t_R FILLER_196_291 ();
 DECAPx2_ASAP7_75t_R FILLER_196_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_307 ();
 DECAPx1_ASAP7_75t_R FILLER_196_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_338 ();
 FILLER_ASAP7_75t_R FILLER_196_342 ();
 DECAPx2_ASAP7_75t_R FILLER_196_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_359 ();
 DECAPx10_ASAP7_75t_R FILLER_196_371 ();
 DECAPx10_ASAP7_75t_R FILLER_196_393 ();
 DECAPx2_ASAP7_75t_R FILLER_196_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_421 ();
 DECAPx6_ASAP7_75t_R FILLER_196_428 ();
 FILLER_ASAP7_75t_R FILLER_196_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_444 ();
 DECAPx10_ASAP7_75t_R FILLER_196_484 ();
 DECAPx10_ASAP7_75t_R FILLER_196_506 ();
 DECAPx2_ASAP7_75t_R FILLER_196_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_534 ();
 DECAPx10_ASAP7_75t_R FILLER_196_542 ();
 DECAPx6_ASAP7_75t_R FILLER_196_564 ();
 DECAPx2_ASAP7_75t_R FILLER_196_578 ();
 DECAPx10_ASAP7_75t_R FILLER_196_592 ();
 DECAPx6_ASAP7_75t_R FILLER_196_614 ();
 DECAPx1_ASAP7_75t_R FILLER_196_628 ();
 DECAPx4_ASAP7_75t_R FILLER_196_634 ();
 FILLER_ASAP7_75t_R FILLER_196_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_646 ();
 DECAPx10_ASAP7_75t_R FILLER_196_657 ();
 DECAPx2_ASAP7_75t_R FILLER_196_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_685 ();
 DECAPx10_ASAP7_75t_R FILLER_196_692 ();
 DECAPx6_ASAP7_75t_R FILLER_196_714 ();
 FILLER_ASAP7_75t_R FILLER_196_728 ();
 DECAPx10_ASAP7_75t_R FILLER_196_748 ();
 DECAPx4_ASAP7_75t_R FILLER_196_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_780 ();
 DECAPx10_ASAP7_75t_R FILLER_196_802 ();
 DECAPx1_ASAP7_75t_R FILLER_196_824 ();
 DECAPx2_ASAP7_75t_R FILLER_196_837 ();
 DECAPx4_ASAP7_75t_R FILLER_196_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_866 ();
 DECAPx10_ASAP7_75t_R FILLER_196_884 ();
 DECAPx10_ASAP7_75t_R FILLER_196_906 ();
 DECAPx10_ASAP7_75t_R FILLER_196_928 ();
 DECAPx1_ASAP7_75t_R FILLER_196_950 ();
 FILLER_ASAP7_75t_R FILLER_196_960 ();
 DECAPx10_ASAP7_75t_R FILLER_196_970 ();
 DECAPx4_ASAP7_75t_R FILLER_196_992 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1173 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_197_172 ();
 FILLER_ASAP7_75t_R FILLER_197_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_180 ();
 DECAPx4_ASAP7_75t_R FILLER_197_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_213 ();
 DECAPx4_ASAP7_75t_R FILLER_197_221 ();
 FILLER_ASAP7_75t_R FILLER_197_231 ();
 DECAPx2_ASAP7_75t_R FILLER_197_241 ();
 FILLER_ASAP7_75t_R FILLER_197_247 ();
 DECAPx2_ASAP7_75t_R FILLER_197_261 ();
 DECAPx10_ASAP7_75t_R FILLER_197_280 ();
 DECAPx6_ASAP7_75t_R FILLER_197_302 ();
 FILLER_ASAP7_75t_R FILLER_197_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_324 ();
 DECAPx10_ASAP7_75t_R FILLER_197_338 ();
 DECAPx1_ASAP7_75t_R FILLER_197_360 ();
 DECAPx10_ASAP7_75t_R FILLER_197_388 ();
 DECAPx10_ASAP7_75t_R FILLER_197_410 ();
 DECAPx10_ASAP7_75t_R FILLER_197_432 ();
 DECAPx2_ASAP7_75t_R FILLER_197_454 ();
 FILLER_ASAP7_75t_R FILLER_197_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_462 ();
 DECAPx1_ASAP7_75t_R FILLER_197_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_473 ();
 DECAPx2_ASAP7_75t_R FILLER_197_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_520 ();
 DECAPx1_ASAP7_75t_R FILLER_197_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_533 ();
 DECAPx6_ASAP7_75t_R FILLER_197_549 ();
 DECAPx10_ASAP7_75t_R FILLER_197_571 ();
 DECAPx10_ASAP7_75t_R FILLER_197_593 ();
 DECAPx4_ASAP7_75t_R FILLER_197_615 ();
 FILLER_ASAP7_75t_R FILLER_197_625 ();
 DECAPx10_ASAP7_75t_R FILLER_197_648 ();
 DECAPx1_ASAP7_75t_R FILLER_197_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_674 ();
 DECAPx10_ASAP7_75t_R FILLER_197_684 ();
 DECAPx10_ASAP7_75t_R FILLER_197_706 ();
 DECAPx10_ASAP7_75t_R FILLER_197_728 ();
 DECAPx6_ASAP7_75t_R FILLER_197_750 ();
 FILLER_ASAP7_75t_R FILLER_197_764 ();
 DECAPx10_ASAP7_75t_R FILLER_197_774 ();
 DECAPx4_ASAP7_75t_R FILLER_197_796 ();
 FILLER_ASAP7_75t_R FILLER_197_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_808 ();
 DECAPx4_ASAP7_75t_R FILLER_197_817 ();
 DECAPx6_ASAP7_75t_R FILLER_197_848 ();
 DECAPx2_ASAP7_75t_R FILLER_197_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_868 ();
 DECAPx4_ASAP7_75t_R FILLER_197_886 ();
 DECAPx4_ASAP7_75t_R FILLER_197_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_917 ();
 DECAPx4_ASAP7_75t_R FILLER_197_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_936 ();
 DECAPx10_ASAP7_75t_R FILLER_197_947 ();
 DECAPx6_ASAP7_75t_R FILLER_197_969 ();
 DECAPx4_ASAP7_75t_R FILLER_197_989 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1045 ();
 FILLER_ASAP7_75t_R FILLER_197_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1102 ();
 FILLER_ASAP7_75t_R FILLER_197_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1150 ();
 FILLER_ASAP7_75t_R FILLER_197_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1165 ();
 FILLER_ASAP7_75t_R FILLER_197_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1173 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1188 ();
 FILLER_ASAP7_75t_R FILLER_197_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_198_172 ();
 DECAPx1_ASAP7_75t_R FILLER_198_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_190 ();
 DECAPx4_ASAP7_75t_R FILLER_198_198 ();
 FILLER_ASAP7_75t_R FILLER_198_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_210 ();
 DECAPx4_ASAP7_75t_R FILLER_198_217 ();
 FILLER_ASAP7_75t_R FILLER_198_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_229 ();
 DECAPx6_ASAP7_75t_R FILLER_198_237 ();
 DECAPx2_ASAP7_75t_R FILLER_198_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_257 ();
 DECAPx1_ASAP7_75t_R FILLER_198_270 ();
 DECAPx10_ASAP7_75t_R FILLER_198_287 ();
 DECAPx10_ASAP7_75t_R FILLER_198_309 ();
 DECAPx10_ASAP7_75t_R FILLER_198_331 ();
 DECAPx10_ASAP7_75t_R FILLER_198_353 ();
 DECAPx1_ASAP7_75t_R FILLER_198_375 ();
 DECAPx10_ASAP7_75t_R FILLER_198_391 ();
 DECAPx10_ASAP7_75t_R FILLER_198_413 ();
 DECAPx2_ASAP7_75t_R FILLER_198_435 ();
 DECAPx2_ASAP7_75t_R FILLER_198_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_457 ();
 DECAPx10_ASAP7_75t_R FILLER_198_485 ();
 DECAPx2_ASAP7_75t_R FILLER_198_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_513 ();
 DECAPx2_ASAP7_75t_R FILLER_198_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_523 ();
 DECAPx1_ASAP7_75t_R FILLER_198_532 ();
 DECAPx1_ASAP7_75t_R FILLER_198_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_547 ();
 FILLER_ASAP7_75t_R FILLER_198_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_558 ();
 DECAPx6_ASAP7_75t_R FILLER_198_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_585 ();
 FILLER_ASAP7_75t_R FILLER_198_589 ();
 FILLER_ASAP7_75t_R FILLER_198_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_599 ();
 DECAPx2_ASAP7_75t_R FILLER_198_608 ();
 FILLER_ASAP7_75t_R FILLER_198_614 ();
 DECAPx4_ASAP7_75t_R FILLER_198_620 ();
 FILLER_ASAP7_75t_R FILLER_198_630 ();
 DECAPx10_ASAP7_75t_R FILLER_198_634 ();
 DECAPx4_ASAP7_75t_R FILLER_198_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_666 ();
 DECAPx10_ASAP7_75t_R FILLER_198_685 ();
 DECAPx6_ASAP7_75t_R FILLER_198_707 ();
 DECAPx1_ASAP7_75t_R FILLER_198_721 ();
 DECAPx10_ASAP7_75t_R FILLER_198_735 ();
 DECAPx10_ASAP7_75t_R FILLER_198_757 ();
 DECAPx10_ASAP7_75t_R FILLER_198_779 ();
 DECAPx4_ASAP7_75t_R FILLER_198_801 ();
 FILLER_ASAP7_75t_R FILLER_198_811 ();
 DECAPx10_ASAP7_75t_R FILLER_198_821 ();
 DECAPx10_ASAP7_75t_R FILLER_198_843 ();
 FILLER_ASAP7_75t_R FILLER_198_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_867 ();
 FILLER_ASAP7_75t_R FILLER_198_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_880 ();
 DECAPx10_ASAP7_75t_R FILLER_198_887 ();
 DECAPx2_ASAP7_75t_R FILLER_198_909 ();
 FILLER_ASAP7_75t_R FILLER_198_915 ();
 DECAPx10_ASAP7_75t_R FILLER_198_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_945 ();
 DECAPx1_ASAP7_75t_R FILLER_198_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_962 ();
 DECAPx1_ASAP7_75t_R FILLER_198_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_977 ();
 DECAPx10_ASAP7_75t_R FILLER_198_984 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1037 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1097 ();
 FILLER_ASAP7_75t_R FILLER_198_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1105 ();
 FILLER_ASAP7_75t_R FILLER_198_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1186 ();
 FILLER_ASAP7_75t_R FILLER_198_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1276 ();
 FILLER_ASAP7_75t_R FILLER_198_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_199_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_194 ();
 DECAPx4_ASAP7_75t_R FILLER_199_202 ();
 FILLER_ASAP7_75t_R FILLER_199_212 ();
 DECAPx2_ASAP7_75t_R FILLER_199_222 ();
 FILLER_ASAP7_75t_R FILLER_199_228 ();
 DECAPx2_ASAP7_75t_R FILLER_199_237 ();
 DECAPx10_ASAP7_75t_R FILLER_199_252 ();
 DECAPx1_ASAP7_75t_R FILLER_199_274 ();
 DECAPx6_ASAP7_75t_R FILLER_199_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_300 ();
 DECAPx10_ASAP7_75t_R FILLER_199_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_331 ();
 DECAPx6_ASAP7_75t_R FILLER_199_348 ();
 FILLER_ASAP7_75t_R FILLER_199_362 ();
 DECAPx4_ASAP7_75t_R FILLER_199_375 ();
 FILLER_ASAP7_75t_R FILLER_199_385 ();
 DECAPx10_ASAP7_75t_R FILLER_199_390 ();
 DECAPx2_ASAP7_75t_R FILLER_199_412 ();
 FILLER_ASAP7_75t_R FILLER_199_418 ();
 DECAPx6_ASAP7_75t_R FILLER_199_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_457 ();
 DECAPx6_ASAP7_75t_R FILLER_199_483 ();
 DECAPx2_ASAP7_75t_R FILLER_199_497 ();
 DECAPx6_ASAP7_75t_R FILLER_199_524 ();
 FILLER_ASAP7_75t_R FILLER_199_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_540 ();
 FILLER_ASAP7_75t_R FILLER_199_570 ();
 DECAPx1_ASAP7_75t_R FILLER_199_593 ();
 DECAPx6_ASAP7_75t_R FILLER_199_618 ();
 DECAPx1_ASAP7_75t_R FILLER_199_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_636 ();
 DECAPx10_ASAP7_75t_R FILLER_199_659 ();
 DECAPx10_ASAP7_75t_R FILLER_199_681 ();
 DECAPx10_ASAP7_75t_R FILLER_199_703 ();
 DECAPx2_ASAP7_75t_R FILLER_199_725 ();
 FILLER_ASAP7_75t_R FILLER_199_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_733 ();
 DECAPx10_ASAP7_75t_R FILLER_199_740 ();
 DECAPx10_ASAP7_75t_R FILLER_199_762 ();
 DECAPx2_ASAP7_75t_R FILLER_199_784 ();
 FILLER_ASAP7_75t_R FILLER_199_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_792 ();
 DECAPx10_ASAP7_75t_R FILLER_199_803 ();
 DECAPx10_ASAP7_75t_R FILLER_199_825 ();
 DECAPx10_ASAP7_75t_R FILLER_199_847 ();
 DECAPx10_ASAP7_75t_R FILLER_199_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_891 ();
 DECAPx10_ASAP7_75t_R FILLER_199_898 ();
 DECAPx10_ASAP7_75t_R FILLER_199_920 ();
 DECAPx10_ASAP7_75t_R FILLER_199_942 ();
 DECAPx6_ASAP7_75t_R FILLER_199_964 ();
 DECAPx2_ASAP7_75t_R FILLER_199_978 ();
 DECAPx2_ASAP7_75t_R FILLER_199_992 ();
 FILLER_ASAP7_75t_R FILLER_199_998 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1021 ();
 FILLER_ASAP7_75t_R FILLER_199_1031 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1039 ();
 FILLER_ASAP7_75t_R FILLER_199_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1141 ();
 FILLER_ASAP7_75t_R FILLER_199_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1279 ();
 DECAPx6_ASAP7_75t_R FILLER_200_172 ();
 FILLER_ASAP7_75t_R FILLER_200_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_188 ();
 FILLER_ASAP7_75t_R FILLER_200_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_203 ();
 DECAPx6_ASAP7_75t_R FILLER_200_218 ();
 FILLER_ASAP7_75t_R FILLER_200_232 ();
 FILLER_ASAP7_75t_R FILLER_200_242 ();
 DECAPx2_ASAP7_75t_R FILLER_200_250 ();
 FILLER_ASAP7_75t_R FILLER_200_256 ();
 FILLER_ASAP7_75t_R FILLER_200_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_268 ();
 DECAPx4_ASAP7_75t_R FILLER_200_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_286 ();
 DECAPx6_ASAP7_75t_R FILLER_200_295 ();
 DECAPx2_ASAP7_75t_R FILLER_200_309 ();
 DECAPx1_ASAP7_75t_R FILLER_200_339 ();
 FILLER_ASAP7_75t_R FILLER_200_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_348 ();
 DECAPx10_ASAP7_75t_R FILLER_200_358 ();
 DECAPx2_ASAP7_75t_R FILLER_200_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_386 ();
 DECAPx2_ASAP7_75t_R FILLER_200_396 ();
 FILLER_ASAP7_75t_R FILLER_200_402 ();
 FILLER_ASAP7_75t_R FILLER_200_410 ();
 DECAPx2_ASAP7_75t_R FILLER_200_418 ();
 DECAPx6_ASAP7_75t_R FILLER_200_432 ();
 FILLER_ASAP7_75t_R FILLER_200_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_448 ();
 DECAPx10_ASAP7_75t_R FILLER_200_473 ();
 DECAPx10_ASAP7_75t_R FILLER_200_495 ();
 DECAPx10_ASAP7_75t_R FILLER_200_517 ();
 DECAPx10_ASAP7_75t_R FILLER_200_539 ();
 DECAPx4_ASAP7_75t_R FILLER_200_561 ();
 FILLER_ASAP7_75t_R FILLER_200_571 ();
 DECAPx10_ASAP7_75t_R FILLER_200_586 ();
 DECAPx10_ASAP7_75t_R FILLER_200_608 ();
 FILLER_ASAP7_75t_R FILLER_200_630 ();
 DECAPx4_ASAP7_75t_R FILLER_200_634 ();
 FILLER_ASAP7_75t_R FILLER_200_644 ();
 DECAPx6_ASAP7_75t_R FILLER_200_662 ();
 DECAPx1_ASAP7_75t_R FILLER_200_676 ();
 DECAPx10_ASAP7_75t_R FILLER_200_694 ();
 DECAPx6_ASAP7_75t_R FILLER_200_716 ();
 DECAPx1_ASAP7_75t_R FILLER_200_730 ();
 DECAPx6_ASAP7_75t_R FILLER_200_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_754 ();
 DECAPx6_ASAP7_75t_R FILLER_200_762 ();
 DECAPx1_ASAP7_75t_R FILLER_200_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_780 ();
 DECAPx10_ASAP7_75t_R FILLER_200_801 ();
 DECAPx2_ASAP7_75t_R FILLER_200_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_852 ();
 DECAPx10_ASAP7_75t_R FILLER_200_865 ();
 DECAPx4_ASAP7_75t_R FILLER_200_887 ();
 FILLER_ASAP7_75t_R FILLER_200_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_899 ();
 DECAPx2_ASAP7_75t_R FILLER_200_908 ();
 FILLER_ASAP7_75t_R FILLER_200_924 ();
 DECAPx10_ASAP7_75t_R FILLER_200_936 ();
 DECAPx1_ASAP7_75t_R FILLER_200_967 ();
 DECAPx10_ASAP7_75t_R FILLER_200_981 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1039 ();
 FILLER_ASAP7_75t_R FILLER_200_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1098 ();
 FILLER_ASAP7_75t_R FILLER_200_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_201_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_204 ();
 DECAPx1_ASAP7_75t_R FILLER_201_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_227 ();
 DECAPx1_ASAP7_75t_R FILLER_201_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_262 ();
 DECAPx2_ASAP7_75t_R FILLER_201_282 ();
 FILLER_ASAP7_75t_R FILLER_201_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_290 ();
 DECAPx4_ASAP7_75t_R FILLER_201_303 ();
 FILLER_ASAP7_75t_R FILLER_201_313 ();
 DECAPx6_ASAP7_75t_R FILLER_201_330 ();
 FILLER_ASAP7_75t_R FILLER_201_344 ();
 DECAPx1_ASAP7_75t_R FILLER_201_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_360 ();
 DECAPx6_ASAP7_75t_R FILLER_201_388 ();
 DECAPx1_ASAP7_75t_R FILLER_201_402 ();
 DECAPx2_ASAP7_75t_R FILLER_201_418 ();
 FILLER_ASAP7_75t_R FILLER_201_424 ();
 DECAPx4_ASAP7_75t_R FILLER_201_432 ();
 DECAPx6_ASAP7_75t_R FILLER_201_459 ();
 FILLER_ASAP7_75t_R FILLER_201_473 ();
 DECAPx4_ASAP7_75t_R FILLER_201_482 ();
 FILLER_ASAP7_75t_R FILLER_201_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_494 ();
 DECAPx4_ASAP7_75t_R FILLER_201_502 ();
 DECAPx10_ASAP7_75t_R FILLER_201_536 ();
 DECAPx2_ASAP7_75t_R FILLER_201_558 ();
 FILLER_ASAP7_75t_R FILLER_201_564 ();
 DECAPx10_ASAP7_75t_R FILLER_201_577 ();
 DECAPx2_ASAP7_75t_R FILLER_201_599 ();
 DECAPx10_ASAP7_75t_R FILLER_201_629 ();
 DECAPx6_ASAP7_75t_R FILLER_201_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_665 ();
 DECAPx10_ASAP7_75t_R FILLER_201_675 ();
 DECAPx10_ASAP7_75t_R FILLER_201_697 ();
 DECAPx10_ASAP7_75t_R FILLER_201_719 ();
 DECAPx10_ASAP7_75t_R FILLER_201_741 ();
 DECAPx10_ASAP7_75t_R FILLER_201_763 ();
 DECAPx6_ASAP7_75t_R FILLER_201_785 ();
 DECAPx10_ASAP7_75t_R FILLER_201_805 ();
 DECAPx10_ASAP7_75t_R FILLER_201_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_849 ();
 DECAPx2_ASAP7_75t_R FILLER_201_862 ();
 FILLER_ASAP7_75t_R FILLER_201_868 ();
 DECAPx10_ASAP7_75t_R FILLER_201_886 ();
 DECAPx6_ASAP7_75t_R FILLER_201_908 ();
 DECAPx1_ASAP7_75t_R FILLER_201_922 ();
 FILLER_ASAP7_75t_R FILLER_201_932 ();
 DECAPx10_ASAP7_75t_R FILLER_201_940 ();
 DECAPx10_ASAP7_75t_R FILLER_201_962 ();
 DECAPx6_ASAP7_75t_R FILLER_201_984 ();
 FILLER_ASAP7_75t_R FILLER_201_998 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1006 ();
 FILLER_ASAP7_75t_R FILLER_201_1012 ();
 FILLER_ASAP7_75t_R FILLER_201_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1033 ();
 FILLER_ASAP7_75t_R FILLER_201_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1062 ();
 FILLER_ASAP7_75t_R FILLER_201_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1074 ();
 FILLER_ASAP7_75t_R FILLER_201_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1134 ();
 FILLER_ASAP7_75t_R FILLER_201_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_202_172 ();
 DECAPx4_ASAP7_75t_R FILLER_202_194 ();
 FILLER_ASAP7_75t_R FILLER_202_204 ();
 DECAPx10_ASAP7_75t_R FILLER_202_209 ();
 FILLER_ASAP7_75t_R FILLER_202_231 ();
 FILLER_ASAP7_75t_R FILLER_202_236 ();
 DECAPx10_ASAP7_75t_R FILLER_202_250 ();
 FILLER_ASAP7_75t_R FILLER_202_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_274 ();
 DECAPx2_ASAP7_75t_R FILLER_202_287 ();
 DECAPx10_ASAP7_75t_R FILLER_202_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_324 ();
 DECAPx2_ASAP7_75t_R FILLER_202_334 ();
 FILLER_ASAP7_75t_R FILLER_202_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_342 ();
 DECAPx10_ASAP7_75t_R FILLER_202_361 ();
 DECAPx2_ASAP7_75t_R FILLER_202_383 ();
 FILLER_ASAP7_75t_R FILLER_202_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_391 ();
 DECAPx10_ASAP7_75t_R FILLER_202_413 ();
 DECAPx4_ASAP7_75t_R FILLER_202_435 ();
 DECAPx4_ASAP7_75t_R FILLER_202_453 ();
 DECAPx2_ASAP7_75t_R FILLER_202_469 ();
 FILLER_ASAP7_75t_R FILLER_202_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_477 ();
 DECAPx1_ASAP7_75t_R FILLER_202_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_504 ();
 FILLER_ASAP7_75t_R FILLER_202_515 ();
 DECAPx6_ASAP7_75t_R FILLER_202_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_539 ();
 DECAPx2_ASAP7_75t_R FILLER_202_548 ();
 FILLER_ASAP7_75t_R FILLER_202_557 ();
 DECAPx1_ASAP7_75t_R FILLER_202_580 ();
 FILLER_ASAP7_75t_R FILLER_202_598 ();
 DECAPx10_ASAP7_75t_R FILLER_202_603 ();
 DECAPx2_ASAP7_75t_R FILLER_202_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_631 ();
 DECAPx10_ASAP7_75t_R FILLER_202_634 ();
 DECAPx10_ASAP7_75t_R FILLER_202_656 ();
 DECAPx2_ASAP7_75t_R FILLER_202_678 ();
 FILLER_ASAP7_75t_R FILLER_202_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_686 ();
 DECAPx10_ASAP7_75t_R FILLER_202_693 ();
 DECAPx1_ASAP7_75t_R FILLER_202_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_719 ();
 DECAPx4_ASAP7_75t_R FILLER_202_734 ();
 DECAPx6_ASAP7_75t_R FILLER_202_753 ();
 FILLER_ASAP7_75t_R FILLER_202_767 ();
 DECAPx10_ASAP7_75t_R FILLER_202_779 ();
 DECAPx10_ASAP7_75t_R FILLER_202_801 ();
 DECAPx10_ASAP7_75t_R FILLER_202_823 ();
 DECAPx10_ASAP7_75t_R FILLER_202_845 ();
 DECAPx6_ASAP7_75t_R FILLER_202_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_881 ();
 DECAPx2_ASAP7_75t_R FILLER_202_892 ();
 FILLER_ASAP7_75t_R FILLER_202_898 ();
 DECAPx10_ASAP7_75t_R FILLER_202_906 ();
 DECAPx6_ASAP7_75t_R FILLER_202_928 ();
 DECAPx1_ASAP7_75t_R FILLER_202_942 ();
 DECAPx10_ASAP7_75t_R FILLER_202_964 ();
 DECAPx2_ASAP7_75t_R FILLER_202_994 ();
 FILLER_ASAP7_75t_R FILLER_202_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1008 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1040 ();
 FILLER_ASAP7_75t_R FILLER_202_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1098 ();
 FILLER_ASAP7_75t_R FILLER_202_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1164 ();
 FILLER_ASAP7_75t_R FILLER_202_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1186 ();
 FILLER_ASAP7_75t_R FILLER_202_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_203_172 ();
 FILLER_ASAP7_75t_R FILLER_203_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_188 ();
 DECAPx1_ASAP7_75t_R FILLER_203_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_203 ();
 DECAPx10_ASAP7_75t_R FILLER_203_220 ();
 DECAPx2_ASAP7_75t_R FILLER_203_242 ();
 FILLER_ASAP7_75t_R FILLER_203_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_250 ();
 DECAPx4_ASAP7_75t_R FILLER_203_266 ();
 FILLER_ASAP7_75t_R FILLER_203_276 ();
 DECAPx4_ASAP7_75t_R FILLER_203_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_297 ();
 DECAPx10_ASAP7_75t_R FILLER_203_301 ();
 FILLER_ASAP7_75t_R FILLER_203_323 ();
 FILLER_ASAP7_75t_R FILLER_203_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_333 ();
 DECAPx10_ASAP7_75t_R FILLER_203_350 ();
 DECAPx10_ASAP7_75t_R FILLER_203_372 ();
 FILLER_ASAP7_75t_R FILLER_203_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_396 ();
 DECAPx6_ASAP7_75t_R FILLER_203_407 ();
 DECAPx2_ASAP7_75t_R FILLER_203_421 ();
 DECAPx6_ASAP7_75t_R FILLER_203_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_449 ();
 DECAPx2_ASAP7_75t_R FILLER_203_490 ();
 DECAPx1_ASAP7_75t_R FILLER_203_513 ();
 DECAPx4_ASAP7_75t_R FILLER_203_523 ();
 FILLER_ASAP7_75t_R FILLER_203_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_535 ();
 DECAPx2_ASAP7_75t_R FILLER_203_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_563 ();
 DECAPx6_ASAP7_75t_R FILLER_203_570 ();
 FILLER_ASAP7_75t_R FILLER_203_584 ();
 DECAPx10_ASAP7_75t_R FILLER_203_607 ();
 DECAPx2_ASAP7_75t_R FILLER_203_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_635 ();
 DECAPx2_ASAP7_75t_R FILLER_203_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_650 ();
 DECAPx10_ASAP7_75t_R FILLER_203_661 ();
 DECAPx10_ASAP7_75t_R FILLER_203_683 ();
 DECAPx1_ASAP7_75t_R FILLER_203_705 ();
 DECAPx1_ASAP7_75t_R FILLER_203_719 ();
 DECAPx10_ASAP7_75t_R FILLER_203_739 ();
 DECAPx10_ASAP7_75t_R FILLER_203_761 ();
 DECAPx6_ASAP7_75t_R FILLER_203_783 ();
 DECAPx2_ASAP7_75t_R FILLER_203_797 ();
 DECAPx10_ASAP7_75t_R FILLER_203_813 ();
 DECAPx10_ASAP7_75t_R FILLER_203_835 ();
 DECAPx10_ASAP7_75t_R FILLER_203_857 ();
 DECAPx4_ASAP7_75t_R FILLER_203_879 ();
 DECAPx6_ASAP7_75t_R FILLER_203_916 ();
 FILLER_ASAP7_75t_R FILLER_203_930 ();
 DECAPx10_ASAP7_75t_R FILLER_203_938 ();
 DECAPx4_ASAP7_75t_R FILLER_203_960 ();
 FILLER_ASAP7_75t_R FILLER_203_970 ();
 DECAPx6_ASAP7_75t_R FILLER_203_982 ();
 DECAPx1_ASAP7_75t_R FILLER_203_996 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1029 ();
 FILLER_ASAP7_75t_R FILLER_203_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1080 ();
 FILLER_ASAP7_75t_R FILLER_203_1086 ();
 FILLER_ASAP7_75t_R FILLER_203_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1168 ();
 FILLER_ASAP7_75t_R FILLER_203_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1269 ();
 FILLER_ASAP7_75t_R FILLER_203_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_204_172 ();
 DECAPx1_ASAP7_75t_R FILLER_204_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_190 ();
 DECAPx2_ASAP7_75t_R FILLER_204_194 ();
 DECAPx2_ASAP7_75t_R FILLER_204_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_227 ();
 DECAPx10_ASAP7_75t_R FILLER_204_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_258 ();
 DECAPx6_ASAP7_75t_R FILLER_204_271 ();
 DECAPx1_ASAP7_75t_R FILLER_204_285 ();
 DECAPx6_ASAP7_75t_R FILLER_204_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_317 ();
 DECAPx1_ASAP7_75t_R FILLER_204_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_331 ();
 DECAPx10_ASAP7_75t_R FILLER_204_347 ();
 DECAPx2_ASAP7_75t_R FILLER_204_369 ();
 FILLER_ASAP7_75t_R FILLER_204_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_377 ();
 DECAPx2_ASAP7_75t_R FILLER_204_390 ();
 DECAPx10_ASAP7_75t_R FILLER_204_408 ();
 DECAPx2_ASAP7_75t_R FILLER_204_430 ();
 FILLER_ASAP7_75t_R FILLER_204_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_438 ();
 DECAPx1_ASAP7_75t_R FILLER_204_444 ();
 DECAPx4_ASAP7_75t_R FILLER_204_453 ();
 FILLER_ASAP7_75t_R FILLER_204_473 ();
 DECAPx10_ASAP7_75t_R FILLER_204_483 ();
 DECAPx10_ASAP7_75t_R FILLER_204_505 ();
 DECAPx4_ASAP7_75t_R FILLER_204_527 ();
 DECAPx2_ASAP7_75t_R FILLER_204_543 ();
 FILLER_ASAP7_75t_R FILLER_204_549 ();
 DECAPx10_ASAP7_75t_R FILLER_204_559 ();
 DECAPx2_ASAP7_75t_R FILLER_204_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_587 ();
 DECAPx10_ASAP7_75t_R FILLER_204_595 ();
 DECAPx6_ASAP7_75t_R FILLER_204_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_631 ();
 FILLER_ASAP7_75t_R FILLER_204_634 ();
 DECAPx10_ASAP7_75t_R FILLER_204_660 ();
 DECAPx4_ASAP7_75t_R FILLER_204_692 ();
 FILLER_ASAP7_75t_R FILLER_204_702 ();
 DECAPx6_ASAP7_75t_R FILLER_204_710 ();
 DECAPx1_ASAP7_75t_R FILLER_204_724 ();
 DECAPx10_ASAP7_75t_R FILLER_204_734 ();
 DECAPx10_ASAP7_75t_R FILLER_204_756 ();
 DECAPx6_ASAP7_75t_R FILLER_204_778 ();
 DECAPx1_ASAP7_75t_R FILLER_204_792 ();
 DECAPx10_ASAP7_75t_R FILLER_204_805 ();
 DECAPx6_ASAP7_75t_R FILLER_204_827 ();
 DECAPx1_ASAP7_75t_R FILLER_204_841 ();
 DECAPx10_ASAP7_75t_R FILLER_204_865 ();
 DECAPx10_ASAP7_75t_R FILLER_204_887 ();
 DECAPx1_ASAP7_75t_R FILLER_204_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_913 ();
 DECAPx1_ASAP7_75t_R FILLER_204_920 ();
 DECAPx10_ASAP7_75t_R FILLER_204_930 ();
 DECAPx6_ASAP7_75t_R FILLER_204_952 ();
 FILLER_ASAP7_75t_R FILLER_204_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_968 ();
 DECAPx6_ASAP7_75t_R FILLER_204_975 ();
 FILLER_ASAP7_75t_R FILLER_204_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_991 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1104 ();
 FILLER_ASAP7_75t_R FILLER_204_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_205_172 ();
 FILLER_ASAP7_75t_R FILLER_205_186 ();
 FILLER_ASAP7_75t_R FILLER_205_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_204 ();
 DECAPx2_ASAP7_75t_R FILLER_205_214 ();
 FILLER_ASAP7_75t_R FILLER_205_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_228 ();
 DECAPx10_ASAP7_75t_R FILLER_205_248 ();
 DECAPx10_ASAP7_75t_R FILLER_205_270 ();
 FILLER_ASAP7_75t_R FILLER_205_292 ();
 DECAPx6_ASAP7_75t_R FILLER_205_303 ();
 FILLER_ASAP7_75t_R FILLER_205_317 ();
 DECAPx4_ASAP7_75t_R FILLER_205_326 ();
 DECAPx6_ASAP7_75t_R FILLER_205_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_377 ();
 DECAPx6_ASAP7_75t_R FILLER_205_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_404 ();
 DECAPx6_ASAP7_75t_R FILLER_205_411 ();
 DECAPx1_ASAP7_75t_R FILLER_205_425 ();
 DECAPx2_ASAP7_75t_R FILLER_205_443 ();
 DECAPx4_ASAP7_75t_R FILLER_205_463 ();
 DECAPx10_ASAP7_75t_R FILLER_205_483 ();
 FILLER_ASAP7_75t_R FILLER_205_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_507 ();
 DECAPx2_ASAP7_75t_R FILLER_205_532 ();
 FILLER_ASAP7_75t_R FILLER_205_538 ();
 DECAPx4_ASAP7_75t_R FILLER_205_546 ();
 FILLER_ASAP7_75t_R FILLER_205_556 ();
 DECAPx1_ASAP7_75t_R FILLER_205_566 ();
 FILLER_ASAP7_75t_R FILLER_205_578 ();
 DECAPx4_ASAP7_75t_R FILLER_205_592 ();
 FILLER_ASAP7_75t_R FILLER_205_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_604 ();
 DECAPx6_ASAP7_75t_R FILLER_205_613 ();
 DECAPx2_ASAP7_75t_R FILLER_205_636 ();
 FILLER_ASAP7_75t_R FILLER_205_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_644 ();
 DECAPx6_ASAP7_75t_R FILLER_205_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_669 ();
 DECAPx10_ASAP7_75t_R FILLER_205_680 ();
 DECAPx10_ASAP7_75t_R FILLER_205_702 ();
 DECAPx10_ASAP7_75t_R FILLER_205_724 ();
 DECAPx10_ASAP7_75t_R FILLER_205_746 ();
 DECAPx10_ASAP7_75t_R FILLER_205_768 ();
 DECAPx6_ASAP7_75t_R FILLER_205_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_804 ();
 DECAPx6_ASAP7_75t_R FILLER_205_811 ();
 DECAPx2_ASAP7_75t_R FILLER_205_825 ();
 DECAPx10_ASAP7_75t_R FILLER_205_838 ();
 DECAPx4_ASAP7_75t_R FILLER_205_860 ();
 FILLER_ASAP7_75t_R FILLER_205_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_872 ();
 DECAPx10_ASAP7_75t_R FILLER_205_885 ();
 DECAPx10_ASAP7_75t_R FILLER_205_917 ();
 DECAPx2_ASAP7_75t_R FILLER_205_945 ();
 FILLER_ASAP7_75t_R FILLER_205_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_953 ();
 DECAPx4_ASAP7_75t_R FILLER_205_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_971 ();
 DECAPx1_ASAP7_75t_R FILLER_205_978 ();
 FILLER_ASAP7_75t_R FILLER_205_992 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1002 ();
 FILLER_ASAP7_75t_R FILLER_205_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1096 ();
 FILLER_ASAP7_75t_R FILLER_205_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1126 ();
 FILLER_ASAP7_75t_R FILLER_205_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1174 ();
 FILLER_ASAP7_75t_R FILLER_205_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1186 ();
 FILLER_ASAP7_75t_R FILLER_205_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1285 ();
 FILLER_ASAP7_75t_R FILLER_205_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_206_172 ();
 FILLER_ASAP7_75t_R FILLER_206_186 ();
 DECAPx2_ASAP7_75t_R FILLER_206_214 ();
 FILLER_ASAP7_75t_R FILLER_206_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_222 ();
 DECAPx10_ASAP7_75t_R FILLER_206_241 ();
 DECAPx2_ASAP7_75t_R FILLER_206_263 ();
 DECAPx2_ASAP7_75t_R FILLER_206_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_316 ();
 DECAPx6_ASAP7_75t_R FILLER_206_325 ();
 DECAPx1_ASAP7_75t_R FILLER_206_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_343 ();
 DECAPx10_ASAP7_75t_R FILLER_206_351 ();
 DECAPx1_ASAP7_75t_R FILLER_206_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_377 ();
 DECAPx2_ASAP7_75t_R FILLER_206_386 ();
 FILLER_ASAP7_75t_R FILLER_206_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_394 ();
 DECAPx1_ASAP7_75t_R FILLER_206_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_404 ();
 DECAPx10_ASAP7_75t_R FILLER_206_421 ();
 DECAPx2_ASAP7_75t_R FILLER_206_443 ();
 FILLER_ASAP7_75t_R FILLER_206_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_451 ();
 DECAPx1_ASAP7_75t_R FILLER_206_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_466 ();
 DECAPx10_ASAP7_75t_R FILLER_206_479 ();
 DECAPx6_ASAP7_75t_R FILLER_206_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_515 ();
 DECAPx6_ASAP7_75t_R FILLER_206_524 ();
 DECAPx1_ASAP7_75t_R FILLER_206_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_542 ();
 DECAPx4_ASAP7_75t_R FILLER_206_554 ();
 DECAPx4_ASAP7_75t_R FILLER_206_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_598 ();
 DECAPx4_ASAP7_75t_R FILLER_206_620 ();
 FILLER_ASAP7_75t_R FILLER_206_630 ();
 DECAPx6_ASAP7_75t_R FILLER_206_634 ();
 FILLER_ASAP7_75t_R FILLER_206_648 ();
 DECAPx10_ASAP7_75t_R FILLER_206_656 ();
 DECAPx4_ASAP7_75t_R FILLER_206_678 ();
 DECAPx2_ASAP7_75t_R FILLER_206_694 ();
 FILLER_ASAP7_75t_R FILLER_206_700 ();
 DECAPx6_ASAP7_75t_R FILLER_206_708 ();
 DECAPx2_ASAP7_75t_R FILLER_206_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_728 ();
 DECAPx4_ASAP7_75t_R FILLER_206_735 ();
 FILLER_ASAP7_75t_R FILLER_206_745 ();
 DECAPx10_ASAP7_75t_R FILLER_206_759 ();
 DECAPx6_ASAP7_75t_R FILLER_206_781 ();
 DECAPx2_ASAP7_75t_R FILLER_206_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_801 ();
 DECAPx6_ASAP7_75t_R FILLER_206_808 ();
 FILLER_ASAP7_75t_R FILLER_206_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_824 ();
 DECAPx10_ASAP7_75t_R FILLER_206_835 ();
 DECAPx6_ASAP7_75t_R FILLER_206_857 ();
 DECAPx1_ASAP7_75t_R FILLER_206_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_875 ();
 DECAPx10_ASAP7_75t_R FILLER_206_882 ();
 DECAPx6_ASAP7_75t_R FILLER_206_920 ();
 FILLER_ASAP7_75t_R FILLER_206_934 ();
 FILLER_ASAP7_75t_R FILLER_206_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_950 ();
 DECAPx10_ASAP7_75t_R FILLER_206_966 ();
 DECAPx10_ASAP7_75t_R FILLER_206_988 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1054 ();
 FILLER_ASAP7_75t_R FILLER_206_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1066 ();
 FILLER_ASAP7_75t_R FILLER_206_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1111 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1122 ();
 FILLER_ASAP7_75t_R FILLER_206_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1140 ();
 FILLER_ASAP7_75t_R FILLER_206_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1194 ();
 FILLER_ASAP7_75t_R FILLER_206_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_207_172 ();
 DECAPx4_ASAP7_75t_R FILLER_207_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_204 ();
 FILLER_ASAP7_75t_R FILLER_207_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_233 ();
 DECAPx1_ASAP7_75t_R FILLER_207_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_259 ();
 DECAPx2_ASAP7_75t_R FILLER_207_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_281 ();
 DECAPx4_ASAP7_75t_R FILLER_207_291 ();
 FILLER_ASAP7_75t_R FILLER_207_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_316 ();
 DECAPx1_ASAP7_75t_R FILLER_207_331 ();
 DECAPx10_ASAP7_75t_R FILLER_207_345 ();
 DECAPx10_ASAP7_75t_R FILLER_207_367 ();
 DECAPx2_ASAP7_75t_R FILLER_207_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_395 ();
 DECAPx4_ASAP7_75t_R FILLER_207_408 ();
 FILLER_ASAP7_75t_R FILLER_207_418 ();
 DECAPx10_ASAP7_75t_R FILLER_207_428 ();
 DECAPx2_ASAP7_75t_R FILLER_207_450 ();
 FILLER_ASAP7_75t_R FILLER_207_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_458 ();
 DECAPx2_ASAP7_75t_R FILLER_207_467 ();
 DECAPx4_ASAP7_75t_R FILLER_207_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_491 ();
 DECAPx4_ASAP7_75t_R FILLER_207_504 ();
 DECAPx6_ASAP7_75t_R FILLER_207_520 ();
 DECAPx1_ASAP7_75t_R FILLER_207_534 ();
 DECAPx2_ASAP7_75t_R FILLER_207_559 ();
 FILLER_ASAP7_75t_R FILLER_207_565 ();
 DECAPx6_ASAP7_75t_R FILLER_207_573 ();
 DECAPx2_ASAP7_75t_R FILLER_207_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_593 ();
 DECAPx1_ASAP7_75t_R FILLER_207_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_631 ();
 DECAPx2_ASAP7_75t_R FILLER_207_638 ();
 DECAPx6_ASAP7_75t_R FILLER_207_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_670 ();
 DECAPx10_ASAP7_75t_R FILLER_207_683 ();
 DECAPx2_ASAP7_75t_R FILLER_207_705 ();
 DECAPx2_ASAP7_75t_R FILLER_207_717 ();
 FILLER_ASAP7_75t_R FILLER_207_723 ();
 DECAPx10_ASAP7_75t_R FILLER_207_731 ();
 DECAPx10_ASAP7_75t_R FILLER_207_753 ();
 DECAPx4_ASAP7_75t_R FILLER_207_775 ();
 FILLER_ASAP7_75t_R FILLER_207_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_787 ();
 DECAPx2_ASAP7_75t_R FILLER_207_794 ();
 DECAPx10_ASAP7_75t_R FILLER_207_822 ();
 DECAPx10_ASAP7_75t_R FILLER_207_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_875 ();
 DECAPx4_ASAP7_75t_R FILLER_207_892 ();
 DECAPx10_ASAP7_75t_R FILLER_207_914 ();
 DECAPx2_ASAP7_75t_R FILLER_207_936 ();
 DECAPx2_ASAP7_75t_R FILLER_207_952 ();
 FILLER_ASAP7_75t_R FILLER_207_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_960 ();
 DECAPx2_ASAP7_75t_R FILLER_207_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_973 ();
 DECAPx1_ASAP7_75t_R FILLER_207_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_984 ();
 DECAPx4_ASAP7_75t_R FILLER_207_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1042 ();
 DECAPx4_ASAP7_75t_R FILLER_207_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1187 ();
 FILLER_ASAP7_75t_R FILLER_207_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_208_172 ();
 DECAPx2_ASAP7_75t_R FILLER_208_194 ();
 FILLER_ASAP7_75t_R FILLER_208_200 ();
 DECAPx1_ASAP7_75t_R FILLER_208_220 ();
 DECAPx6_ASAP7_75t_R FILLER_208_233 ();
 DECAPx1_ASAP7_75t_R FILLER_208_247 ();
 DECAPx2_ASAP7_75t_R FILLER_208_258 ();
 DECAPx10_ASAP7_75t_R FILLER_208_278 ();
 DECAPx2_ASAP7_75t_R FILLER_208_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_306 ();
 FILLER_ASAP7_75t_R FILLER_208_313 ();
 DECAPx2_ASAP7_75t_R FILLER_208_322 ();
 FILLER_ASAP7_75t_R FILLER_208_340 ();
 DECAPx10_ASAP7_75t_R FILLER_208_348 ();
 DECAPx1_ASAP7_75t_R FILLER_208_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_374 ();
 DECAPx4_ASAP7_75t_R FILLER_208_381 ();
 FILLER_ASAP7_75t_R FILLER_208_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_393 ();
 DECAPx2_ASAP7_75t_R FILLER_208_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_406 ();
 DECAPx2_ASAP7_75t_R FILLER_208_429 ();
 FILLER_ASAP7_75t_R FILLER_208_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_437 ();
 DECAPx10_ASAP7_75t_R FILLER_208_448 ();
 DECAPx1_ASAP7_75t_R FILLER_208_490 ();
 DECAPx4_ASAP7_75t_R FILLER_208_510 ();
 FILLER_ASAP7_75t_R FILLER_208_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_522 ();
 DECAPx10_ASAP7_75t_R FILLER_208_535 ();
 FILLER_ASAP7_75t_R FILLER_208_557 ();
 DECAPx2_ASAP7_75t_R FILLER_208_580 ();
 FILLER_ASAP7_75t_R FILLER_208_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_588 ();
 DECAPx10_ASAP7_75t_R FILLER_208_592 ();
 DECAPx6_ASAP7_75t_R FILLER_208_614 ();
 DECAPx1_ASAP7_75t_R FILLER_208_628 ();
 DECAPx10_ASAP7_75t_R FILLER_208_634 ();
 DECAPx4_ASAP7_75t_R FILLER_208_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_666 ();
 DECAPx10_ASAP7_75t_R FILLER_208_677 ();
 DECAPx6_ASAP7_75t_R FILLER_208_699 ();
 FILLER_ASAP7_75t_R FILLER_208_713 ();
 DECAPx10_ASAP7_75t_R FILLER_208_737 ();
 DECAPx10_ASAP7_75t_R FILLER_208_759 ();
 DECAPx2_ASAP7_75t_R FILLER_208_781 ();
 FILLER_ASAP7_75t_R FILLER_208_787 ();
 DECAPx10_ASAP7_75t_R FILLER_208_811 ();
 DECAPx6_ASAP7_75t_R FILLER_208_833 ();
 DECAPx1_ASAP7_75t_R FILLER_208_847 ();
 DECAPx2_ASAP7_75t_R FILLER_208_859 ();
 FILLER_ASAP7_75t_R FILLER_208_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_867 ();
 DECAPx10_ASAP7_75t_R FILLER_208_878 ();
 DECAPx10_ASAP7_75t_R FILLER_208_900 ();
 DECAPx6_ASAP7_75t_R FILLER_208_922 ();
 FILLER_ASAP7_75t_R FILLER_208_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_938 ();
 DECAPx6_ASAP7_75t_R FILLER_208_947 ();
 FILLER_ASAP7_75t_R FILLER_208_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_963 ();
 DECAPx10_ASAP7_75t_R FILLER_208_976 ();
 DECAPx4_ASAP7_75t_R FILLER_208_998 ();
 FILLER_ASAP7_75t_R FILLER_208_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1079 ();
 FILLER_ASAP7_75t_R FILLER_208_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1184 ();
 FILLER_ASAP7_75t_R FILLER_208_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1277 ();
 FILLER_ASAP7_75t_R FILLER_208_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_209_172 ();
 DECAPx2_ASAP7_75t_R FILLER_209_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_200 ();
 DECAPx10_ASAP7_75t_R FILLER_209_216 ();
 DECAPx10_ASAP7_75t_R FILLER_209_238 ();
 DECAPx10_ASAP7_75t_R FILLER_209_260 ();
 DECAPx2_ASAP7_75t_R FILLER_209_282 ();
 FILLER_ASAP7_75t_R FILLER_209_288 ();
 DECAPx6_ASAP7_75t_R FILLER_209_297 ();
 DECAPx2_ASAP7_75t_R FILLER_209_311 ();
 DECAPx6_ASAP7_75t_R FILLER_209_324 ();
 FILLER_ASAP7_75t_R FILLER_209_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_340 ();
 DECAPx4_ASAP7_75t_R FILLER_209_350 ();
 FILLER_ASAP7_75t_R FILLER_209_360 ();
 DECAPx2_ASAP7_75t_R FILLER_209_374 ();
 FILLER_ASAP7_75t_R FILLER_209_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_390 ();
 DECAPx6_ASAP7_75t_R FILLER_209_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_415 ();
 DECAPx2_ASAP7_75t_R FILLER_209_448 ();
 DECAPx10_ASAP7_75t_R FILLER_209_474 ();
 DECAPx6_ASAP7_75t_R FILLER_209_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_510 ();
 DECAPx1_ASAP7_75t_R FILLER_209_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_523 ();
 DECAPx6_ASAP7_75t_R FILLER_209_532 ();
 DECAPx2_ASAP7_75t_R FILLER_209_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_552 ();
 DECAPx2_ASAP7_75t_R FILLER_209_567 ();
 FILLER_ASAP7_75t_R FILLER_209_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_575 ();
 DECAPx10_ASAP7_75t_R FILLER_209_593 ();
 DECAPx10_ASAP7_75t_R FILLER_209_615 ();
 DECAPx4_ASAP7_75t_R FILLER_209_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_647 ();
 DECAPx1_ASAP7_75t_R FILLER_209_657 ();
 DECAPx10_ASAP7_75t_R FILLER_209_668 ();
 DECAPx6_ASAP7_75t_R FILLER_209_690 ();
 FILLER_ASAP7_75t_R FILLER_209_704 ();
 DECAPx2_ASAP7_75t_R FILLER_209_712 ();
 FILLER_ASAP7_75t_R FILLER_209_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_720 ();
 DECAPx10_ASAP7_75t_R FILLER_209_727 ();
 DECAPx10_ASAP7_75t_R FILLER_209_749 ();
 DECAPx10_ASAP7_75t_R FILLER_209_780 ();
 DECAPx10_ASAP7_75t_R FILLER_209_802 ();
 DECAPx10_ASAP7_75t_R FILLER_209_824 ();
 FILLER_ASAP7_75t_R FILLER_209_846 ();
 DECAPx10_ASAP7_75t_R FILLER_209_860 ();
 DECAPx10_ASAP7_75t_R FILLER_209_882 ();
 DECAPx4_ASAP7_75t_R FILLER_209_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_914 ();
 DECAPx2_ASAP7_75t_R FILLER_209_927 ();
 FILLER_ASAP7_75t_R FILLER_209_933 ();
 DECAPx6_ASAP7_75t_R FILLER_209_971 ();
 DECAPx2_ASAP7_75t_R FILLER_209_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_991 ();
 FILLER_ASAP7_75t_R FILLER_209_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_210_172 ();
 FILLER_ASAP7_75t_R FILLER_210_186 ();
 DECAPx2_ASAP7_75t_R FILLER_210_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_200 ();
 FILLER_ASAP7_75t_R FILLER_210_208 ();
 FILLER_ASAP7_75t_R FILLER_210_219 ();
 DECAPx10_ASAP7_75t_R FILLER_210_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_246 ();
 FILLER_ASAP7_75t_R FILLER_210_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_256 ();
 DECAPx10_ASAP7_75t_R FILLER_210_261 ();
 DECAPx4_ASAP7_75t_R FILLER_210_283 ();
 FILLER_ASAP7_75t_R FILLER_210_293 ();
 DECAPx1_ASAP7_75t_R FILLER_210_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_319 ();
 DECAPx2_ASAP7_75t_R FILLER_210_327 ();
 FILLER_ASAP7_75t_R FILLER_210_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_335 ();
 DECAPx1_ASAP7_75t_R FILLER_210_356 ();
 DECAPx6_ASAP7_75t_R FILLER_210_369 ();
 FILLER_ASAP7_75t_R FILLER_210_383 ();
 FILLER_ASAP7_75t_R FILLER_210_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_393 ();
 DECAPx10_ASAP7_75t_R FILLER_210_404 ();
 DECAPx6_ASAP7_75t_R FILLER_210_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_440 ();
 DECAPx4_ASAP7_75t_R FILLER_210_455 ();
 FILLER_ASAP7_75t_R FILLER_210_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_467 ();
 FILLER_ASAP7_75t_R FILLER_210_496 ();
 DECAPx1_ASAP7_75t_R FILLER_210_512 ();
 DECAPx2_ASAP7_75t_R FILLER_210_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_546 ();
 DECAPx6_ASAP7_75t_R FILLER_210_558 ();
 DECAPx2_ASAP7_75t_R FILLER_210_572 ();
 DECAPx10_ASAP7_75t_R FILLER_210_599 ();
 DECAPx4_ASAP7_75t_R FILLER_210_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_631 ();
 FILLER_ASAP7_75t_R FILLER_210_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_636 ();
 DECAPx6_ASAP7_75t_R FILLER_210_647 ();
 FILLER_ASAP7_75t_R FILLER_210_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_663 ();
 DECAPx10_ASAP7_75t_R FILLER_210_670 ();
 DECAPx6_ASAP7_75t_R FILLER_210_692 ();
 FILLER_ASAP7_75t_R FILLER_210_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_708 ();
 DECAPx2_ASAP7_75t_R FILLER_210_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_725 ();
 DECAPx6_ASAP7_75t_R FILLER_210_732 ();
 DECAPx2_ASAP7_75t_R FILLER_210_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_752 ();
 DECAPx4_ASAP7_75t_R FILLER_210_759 ();
 FILLER_ASAP7_75t_R FILLER_210_775 ();
 DECAPx10_ASAP7_75t_R FILLER_210_783 ();
 DECAPx10_ASAP7_75t_R FILLER_210_805 ();
 FILLER_ASAP7_75t_R FILLER_210_827 ();
 FILLER_ASAP7_75t_R FILLER_210_839 ();
 FILLER_ASAP7_75t_R FILLER_210_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_883 ();
 DECAPx1_ASAP7_75t_R FILLER_210_900 ();
 DECAPx4_ASAP7_75t_R FILLER_210_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_921 ();
 FILLER_ASAP7_75t_R FILLER_210_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_934 ();
 DECAPx2_ASAP7_75t_R FILLER_210_983 ();
 FILLER_ASAP7_75t_R FILLER_210_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_991 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1022 ();
 FILLER_ASAP7_75t_R FILLER_210_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1096 ();
 FILLER_ASAP7_75t_R FILLER_210_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1124 ();
 FILLER_ASAP7_75t_R FILLER_210_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_210_1162 ();
 FILLER_ASAP7_75t_R FILLER_210_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1193 ();
 FILLER_ASAP7_75t_R FILLER_210_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_210_1280 ();
 FILLER_ASAP7_75t_R FILLER_210_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_211_172 ();
 FILLER_ASAP7_75t_R FILLER_211_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_184 ();
 FILLER_ASAP7_75t_R FILLER_211_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_201 ();
 FILLER_ASAP7_75t_R FILLER_211_209 ();
 DECAPx6_ASAP7_75t_R FILLER_211_219 ();
 FILLER_ASAP7_75t_R FILLER_211_233 ();
 DECAPx2_ASAP7_75t_R FILLER_211_242 ();
 FILLER_ASAP7_75t_R FILLER_211_248 ();
 DECAPx2_ASAP7_75t_R FILLER_211_257 ();
 DECAPx4_ASAP7_75t_R FILLER_211_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_288 ();
 DECAPx2_ASAP7_75t_R FILLER_211_301 ();
 FILLER_ASAP7_75t_R FILLER_211_307 ();
 DECAPx1_ASAP7_75t_R FILLER_211_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_319 ();
 DECAPx2_ASAP7_75t_R FILLER_211_326 ();
 FILLER_ASAP7_75t_R FILLER_211_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_334 ();
 DECAPx1_ASAP7_75t_R FILLER_211_342 ();
 FILLER_ASAP7_75t_R FILLER_211_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_355 ();
 DECAPx4_ASAP7_75t_R FILLER_211_362 ();
 FILLER_ASAP7_75t_R FILLER_211_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_374 ();
 DECAPx2_ASAP7_75t_R FILLER_211_388 ();
 FILLER_ASAP7_75t_R FILLER_211_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_396 ();
 DECAPx2_ASAP7_75t_R FILLER_211_409 ();
 FILLER_ASAP7_75t_R FILLER_211_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_417 ();
 DECAPx6_ASAP7_75t_R FILLER_211_424 ();
 DECAPx1_ASAP7_75t_R FILLER_211_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_442 ();
 DECAPx2_ASAP7_75t_R FILLER_211_451 ();
 FILLER_ASAP7_75t_R FILLER_211_457 ();
 DECAPx10_ASAP7_75t_R FILLER_211_478 ();
 DECAPx6_ASAP7_75t_R FILLER_211_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_514 ();
 DECAPx6_ASAP7_75t_R FILLER_211_523 ();
 FILLER_ASAP7_75t_R FILLER_211_537 ();
 DECAPx10_ASAP7_75t_R FILLER_211_560 ();
 DECAPx10_ASAP7_75t_R FILLER_211_582 ();
 DECAPx10_ASAP7_75t_R FILLER_211_604 ();
 DECAPx2_ASAP7_75t_R FILLER_211_626 ();
 FILLER_ASAP7_75t_R FILLER_211_632 ();
 DECAPx10_ASAP7_75t_R FILLER_211_646 ();
 DECAPx10_ASAP7_75t_R FILLER_211_668 ();
 DECAPx4_ASAP7_75t_R FILLER_211_690 ();
 DECAPx6_ASAP7_75t_R FILLER_211_710 ();
 DECAPx1_ASAP7_75t_R FILLER_211_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_728 ();
 DECAPx6_ASAP7_75t_R FILLER_211_736 ();
 FILLER_ASAP7_75t_R FILLER_211_750 ();
 DECAPx10_ASAP7_75t_R FILLER_211_758 ();
 DECAPx10_ASAP7_75t_R FILLER_211_780 ();
 DECAPx2_ASAP7_75t_R FILLER_211_802 ();
 DECAPx10_ASAP7_75t_R FILLER_211_818 ();
 DECAPx2_ASAP7_75t_R FILLER_211_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_846 ();
 DECAPx1_ASAP7_75t_R FILLER_211_877 ();
 DECAPx1_ASAP7_75t_R FILLER_211_887 ();
 DECAPx4_ASAP7_75t_R FILLER_211_901 ();
 FILLER_ASAP7_75t_R FILLER_211_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_913 ();
 DECAPx4_ASAP7_75t_R FILLER_211_920 ();
 FILLER_ASAP7_75t_R FILLER_211_930 ();
 DECAPx1_ASAP7_75t_R FILLER_211_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_949 ();
 DECAPx10_ASAP7_75t_R FILLER_211_956 ();
 DECAPx4_ASAP7_75t_R FILLER_211_978 ();
 FILLER_ASAP7_75t_R FILLER_211_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_990 ();
 FILLER_ASAP7_75t_R FILLER_211_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1028 ();
 FILLER_ASAP7_75t_R FILLER_211_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1050 ();
 FILLER_ASAP7_75t_R FILLER_211_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1070 ();
 FILLER_ASAP7_75t_R FILLER_211_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_211_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_211_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_212_172 ();
 DECAPx2_ASAP7_75t_R FILLER_212_201 ();
 FILLER_ASAP7_75t_R FILLER_212_207 ();
 DECAPx1_ASAP7_75t_R FILLER_212_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_219 ();
 DECAPx2_ASAP7_75t_R FILLER_212_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_235 ();
 FILLER_ASAP7_75t_R FILLER_212_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_267 ();
 DECAPx4_ASAP7_75t_R FILLER_212_297 ();
 FILLER_ASAP7_75t_R FILLER_212_307 ();
 FILLER_ASAP7_75t_R FILLER_212_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_317 ();
 DECAPx10_ASAP7_75t_R FILLER_212_341 ();
 DECAPx10_ASAP7_75t_R FILLER_212_363 ();
 DECAPx2_ASAP7_75t_R FILLER_212_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_391 ();
 FILLER_ASAP7_75t_R FILLER_212_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_400 ();
 DECAPx4_ASAP7_75t_R FILLER_212_409 ();
 FILLER_ASAP7_75t_R FILLER_212_419 ();
 DECAPx10_ASAP7_75t_R FILLER_212_429 ();
 DECAPx10_ASAP7_75t_R FILLER_212_451 ();
 DECAPx6_ASAP7_75t_R FILLER_212_473 ();
 FILLER_ASAP7_75t_R FILLER_212_487 ();
 DECAPx10_ASAP7_75t_R FILLER_212_499 ();
 DECAPx1_ASAP7_75t_R FILLER_212_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_525 ();
 DECAPx10_ASAP7_75t_R FILLER_212_532 ();
 DECAPx10_ASAP7_75t_R FILLER_212_554 ();
 DECAPx4_ASAP7_75t_R FILLER_212_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_586 ();
 FILLER_ASAP7_75t_R FILLER_212_595 ();
 FILLER_ASAP7_75t_R FILLER_212_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_613 ();
 DECAPx4_ASAP7_75t_R FILLER_212_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_634 ();
 DECAPx2_ASAP7_75t_R FILLER_212_656 ();
 DECAPx10_ASAP7_75t_R FILLER_212_672 ();
 DECAPx6_ASAP7_75t_R FILLER_212_694 ();
 FILLER_ASAP7_75t_R FILLER_212_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_710 ();
 FILLER_ASAP7_75t_R FILLER_212_717 ();
 DECAPx10_ASAP7_75t_R FILLER_212_725 ();
 DECAPx4_ASAP7_75t_R FILLER_212_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_757 ();
 DECAPx6_ASAP7_75t_R FILLER_212_761 ();
 DECAPx1_ASAP7_75t_R FILLER_212_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_789 ();
 DECAPx6_ASAP7_75t_R FILLER_212_798 ();
 DECAPx1_ASAP7_75t_R FILLER_212_812 ();
 DECAPx6_ASAP7_75t_R FILLER_212_824 ();
 DECAPx1_ASAP7_75t_R FILLER_212_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_842 ();
 DECAPx6_ASAP7_75t_R FILLER_212_849 ();
 DECAPx6_ASAP7_75t_R FILLER_212_871 ();
 DECAPx1_ASAP7_75t_R FILLER_212_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_889 ();
 DECAPx10_ASAP7_75t_R FILLER_212_896 ();
 DECAPx6_ASAP7_75t_R FILLER_212_918 ();
 DECAPx1_ASAP7_75t_R FILLER_212_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_936 ();
 DECAPx6_ASAP7_75t_R FILLER_212_943 ();
 DECAPx1_ASAP7_75t_R FILLER_212_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_961 ();
 DECAPx10_ASAP7_75t_R FILLER_212_971 ();
 DECAPx6_ASAP7_75t_R FILLER_212_993 ();
 FILLER_ASAP7_75t_R FILLER_212_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1040 ();
 FILLER_ASAP7_75t_R FILLER_212_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1063 ();
 FILLER_ASAP7_75t_R FILLER_212_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1082 ();
 FILLER_ASAP7_75t_R FILLER_212_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1148 ();
 FILLER_ASAP7_75t_R FILLER_212_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1277 ();
 FILLER_ASAP7_75t_R FILLER_212_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_213_172 ();
 FILLER_ASAP7_75t_R FILLER_213_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_191 ();
 DECAPx1_ASAP7_75t_R FILLER_213_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_215 ();
 DECAPx1_ASAP7_75t_R FILLER_213_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_233 ();
 DECAPx10_ASAP7_75t_R FILLER_213_242 ();
 DECAPx4_ASAP7_75t_R FILLER_213_264 ();
 FILLER_ASAP7_75t_R FILLER_213_280 ();
 FILLER_ASAP7_75t_R FILLER_213_294 ();
 DECAPx10_ASAP7_75t_R FILLER_213_308 ();
 DECAPx1_ASAP7_75t_R FILLER_213_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_334 ();
 DECAPx1_ASAP7_75t_R FILLER_213_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_352 ();
 DECAPx4_ASAP7_75t_R FILLER_213_362 ();
 FILLER_ASAP7_75t_R FILLER_213_372 ();
 DECAPx10_ASAP7_75t_R FILLER_213_388 ();
 DECAPx1_ASAP7_75t_R FILLER_213_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_414 ();
 DECAPx4_ASAP7_75t_R FILLER_213_425 ();
 FILLER_ASAP7_75t_R FILLER_213_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_437 ();
 DECAPx10_ASAP7_75t_R FILLER_213_458 ();
 DECAPx1_ASAP7_75t_R FILLER_213_480 ();
 DECAPx10_ASAP7_75t_R FILLER_213_492 ();
 DECAPx4_ASAP7_75t_R FILLER_213_514 ();
 FILLER_ASAP7_75t_R FILLER_213_524 ();
 FILLER_ASAP7_75t_R FILLER_213_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_536 ();
 DECAPx2_ASAP7_75t_R FILLER_213_540 ();
 FILLER_ASAP7_75t_R FILLER_213_554 ();
 DECAPx2_ASAP7_75t_R FILLER_213_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_565 ();
 DECAPx1_ASAP7_75t_R FILLER_213_580 ();
 DECAPx1_ASAP7_75t_R FILLER_213_587 ();
 DECAPx6_ASAP7_75t_R FILLER_213_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_611 ();
 DECAPx10_ASAP7_75t_R FILLER_213_615 ();
 DECAPx6_ASAP7_75t_R FILLER_213_637 ();
 FILLER_ASAP7_75t_R FILLER_213_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_653 ();
 DECAPx10_ASAP7_75t_R FILLER_213_672 ();
 DECAPx10_ASAP7_75t_R FILLER_213_694 ();
 DECAPx10_ASAP7_75t_R FILLER_213_722 ();
 DECAPx10_ASAP7_75t_R FILLER_213_744 ();
 DECAPx6_ASAP7_75t_R FILLER_213_766 ();
 DECAPx2_ASAP7_75t_R FILLER_213_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_786 ();
 DECAPx10_ASAP7_75t_R FILLER_213_797 ();
 DECAPx2_ASAP7_75t_R FILLER_213_819 ();
 DECAPx6_ASAP7_75t_R FILLER_213_831 ();
 FILLER_ASAP7_75t_R FILLER_213_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_847 ();
 DECAPx4_ASAP7_75t_R FILLER_213_856 ();
 FILLER_ASAP7_75t_R FILLER_213_866 ();
 DECAPx4_ASAP7_75t_R FILLER_213_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_888 ();
 DECAPx10_ASAP7_75t_R FILLER_213_895 ();
 DECAPx6_ASAP7_75t_R FILLER_213_917 ();
 DECAPx1_ASAP7_75t_R FILLER_213_931 ();
 DECAPx10_ASAP7_75t_R FILLER_213_941 ();
 DECAPx10_ASAP7_75t_R FILLER_213_963 ();
 DECAPx6_ASAP7_75t_R FILLER_213_985 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1031 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1118 ();
 FILLER_ASAP7_75t_R FILLER_213_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_214_172 ();
 DECAPx6_ASAP7_75t_R FILLER_214_194 ();
 DECAPx1_ASAP7_75t_R FILLER_214_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_212 ();
 DECAPx4_ASAP7_75t_R FILLER_214_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_235 ();
 DECAPx10_ASAP7_75t_R FILLER_214_242 ();
 DECAPx1_ASAP7_75t_R FILLER_214_264 ();
 DECAPx2_ASAP7_75t_R FILLER_214_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_277 ();
 DECAPx6_ASAP7_75t_R FILLER_214_284 ();
 FILLER_ASAP7_75t_R FILLER_214_298 ();
 FILLER_ASAP7_75t_R FILLER_214_306 ();
 DECAPx2_ASAP7_75t_R FILLER_214_317 ();
 FILLER_ASAP7_75t_R FILLER_214_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_325 ();
 DECAPx1_ASAP7_75t_R FILLER_214_334 ();
 DECAPx4_ASAP7_75t_R FILLER_214_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_355 ();
 DECAPx4_ASAP7_75t_R FILLER_214_368 ();
 DECAPx2_ASAP7_75t_R FILLER_214_384 ();
 DECAPx2_ASAP7_75t_R FILLER_214_440 ();
 FILLER_ASAP7_75t_R FILLER_214_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_448 ();
 DECAPx1_ASAP7_75t_R FILLER_214_457 ();
 DECAPx10_ASAP7_75t_R FILLER_214_479 ();
 DECAPx2_ASAP7_75t_R FILLER_214_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_507 ();
 FILLER_ASAP7_75t_R FILLER_214_516 ();
 DECAPx1_ASAP7_75t_R FILLER_214_539 ();
 DECAPx1_ASAP7_75t_R FILLER_214_564 ();
 DECAPx1_ASAP7_75t_R FILLER_214_589 ();
 DECAPx6_ASAP7_75t_R FILLER_214_614 ();
 DECAPx1_ASAP7_75t_R FILLER_214_628 ();
 DECAPx10_ASAP7_75t_R FILLER_214_644 ();
 DECAPx6_ASAP7_75t_R FILLER_214_666 ();
 DECAPx6_ASAP7_75t_R FILLER_214_690 ();
 FILLER_ASAP7_75t_R FILLER_214_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_706 ();
 DECAPx6_ASAP7_75t_R FILLER_214_713 ();
 DECAPx1_ASAP7_75t_R FILLER_214_727 ();
 DECAPx10_ASAP7_75t_R FILLER_214_739 ();
 DECAPx10_ASAP7_75t_R FILLER_214_761 ();
 DECAPx2_ASAP7_75t_R FILLER_214_783 ();
 FILLER_ASAP7_75t_R FILLER_214_789 ();
 DECAPx2_ASAP7_75t_R FILLER_214_797 ();
 FILLER_ASAP7_75t_R FILLER_214_803 ();
 DECAPx10_ASAP7_75t_R FILLER_214_811 ();
 DECAPx6_ASAP7_75t_R FILLER_214_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_847 ();
 DECAPx10_ASAP7_75t_R FILLER_214_856 ();
 DECAPx10_ASAP7_75t_R FILLER_214_878 ();
 DECAPx1_ASAP7_75t_R FILLER_214_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_904 ();
 DECAPx1_ASAP7_75t_R FILLER_214_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_923 ();
 DECAPx1_ASAP7_75t_R FILLER_214_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_934 ();
 DECAPx6_ASAP7_75t_R FILLER_214_944 ();
 FILLER_ASAP7_75t_R FILLER_214_958 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1117 ();
 FILLER_ASAP7_75t_R FILLER_214_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1177 ();
 FILLER_ASAP7_75t_R FILLER_214_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1280 ();
 FILLER_ASAP7_75t_R FILLER_214_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_215_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_194 ();
 FILLER_ASAP7_75t_R FILLER_215_203 ();
 DECAPx10_ASAP7_75t_R FILLER_215_212 ();
 FILLER_ASAP7_75t_R FILLER_215_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_236 ();
 DECAPx4_ASAP7_75t_R FILLER_215_251 ();
 FILLER_ASAP7_75t_R FILLER_215_267 ();
 DECAPx1_ASAP7_75t_R FILLER_215_287 ();
 DECAPx10_ASAP7_75t_R FILLER_215_297 ();
 DECAPx10_ASAP7_75t_R FILLER_215_319 ();
 DECAPx6_ASAP7_75t_R FILLER_215_341 ();
 FILLER_ASAP7_75t_R FILLER_215_355 ();
 DECAPx2_ASAP7_75t_R FILLER_215_367 ();
 FILLER_ASAP7_75t_R FILLER_215_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_382 ();
 DECAPx10_ASAP7_75t_R FILLER_215_393 ();
 DECAPx10_ASAP7_75t_R FILLER_215_415 ();
 DECAPx6_ASAP7_75t_R FILLER_215_437 ();
 FILLER_ASAP7_75t_R FILLER_215_482 ();
 FILLER_ASAP7_75t_R FILLER_215_490 ();
 DECAPx10_ASAP7_75t_R FILLER_215_512 ();
 DECAPx4_ASAP7_75t_R FILLER_215_534 ();
 DECAPx10_ASAP7_75t_R FILLER_215_550 ();
 DECAPx6_ASAP7_75t_R FILLER_215_572 ();
 FILLER_ASAP7_75t_R FILLER_215_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_588 ();
 DECAPx10_ASAP7_75t_R FILLER_215_597 ();
 DECAPx10_ASAP7_75t_R FILLER_215_619 ();
 DECAPx6_ASAP7_75t_R FILLER_215_641 ();
 DECAPx1_ASAP7_75t_R FILLER_215_655 ();
 DECAPx4_ASAP7_75t_R FILLER_215_662 ();
 DECAPx10_ASAP7_75t_R FILLER_215_682 ();
 FILLER_ASAP7_75t_R FILLER_215_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_706 ();
 DECAPx10_ASAP7_75t_R FILLER_215_729 ();
 DECAPx6_ASAP7_75t_R FILLER_215_751 ();
 DECAPx1_ASAP7_75t_R FILLER_215_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_769 ();
 DECAPx6_ASAP7_75t_R FILLER_215_776 ();
 FILLER_ASAP7_75t_R FILLER_215_790 ();
 DECAPx2_ASAP7_75t_R FILLER_215_798 ();
 DECAPx4_ASAP7_75t_R FILLER_215_810 ();
 FILLER_ASAP7_75t_R FILLER_215_820 ();
 DECAPx10_ASAP7_75t_R FILLER_215_828 ();
 DECAPx10_ASAP7_75t_R FILLER_215_850 ();
 DECAPx2_ASAP7_75t_R FILLER_215_872 ();
 FILLER_ASAP7_75t_R FILLER_215_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_880 ();
 DECAPx4_ASAP7_75t_R FILLER_215_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_908 ();
 DECAPx4_ASAP7_75t_R FILLER_215_915 ();
 FILLER_ASAP7_75t_R FILLER_215_925 ();
 DECAPx1_ASAP7_75t_R FILLER_215_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_937 ();
 DECAPx1_ASAP7_75t_R FILLER_215_950 ();
 FILLER_ASAP7_75t_R FILLER_215_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_968 ();
 DECAPx6_ASAP7_75t_R FILLER_215_977 ();
 FILLER_ASAP7_75t_R FILLER_215_991 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1019 ();
 FILLER_ASAP7_75t_R FILLER_215_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1036 ();
 FILLER_ASAP7_75t_R FILLER_215_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1056 ();
 FILLER_ASAP7_75t_R FILLER_215_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1152 ();
 FILLER_ASAP7_75t_R FILLER_215_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_215_1182 ();
 FILLER_ASAP7_75t_R FILLER_215_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_216_172 ();
 FILLER_ASAP7_75t_R FILLER_216_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_184 ();
 DECAPx4_ASAP7_75t_R FILLER_216_194 ();
 FILLER_ASAP7_75t_R FILLER_216_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_206 ();
 DECAPx1_ASAP7_75t_R FILLER_216_219 ();
 DECAPx6_ASAP7_75t_R FILLER_216_263 ();
 DECAPx2_ASAP7_75t_R FILLER_216_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_283 ();
 DECAPx1_ASAP7_75t_R FILLER_216_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_294 ();
 FILLER_ASAP7_75t_R FILLER_216_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_303 ();
 DECAPx1_ASAP7_75t_R FILLER_216_312 ();
 DECAPx4_ASAP7_75t_R FILLER_216_326 ();
 FILLER_ASAP7_75t_R FILLER_216_336 ();
 DECAPx10_ASAP7_75t_R FILLER_216_346 ();
 DECAPx1_ASAP7_75t_R FILLER_216_368 ();
 DECAPx6_ASAP7_75t_R FILLER_216_380 ();
 DECAPx2_ASAP7_75t_R FILLER_216_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_410 ();
 DECAPx4_ASAP7_75t_R FILLER_216_417 ();
 DECAPx10_ASAP7_75t_R FILLER_216_442 ();
 DECAPx2_ASAP7_75t_R FILLER_216_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_481 ();
 DECAPx10_ASAP7_75t_R FILLER_216_500 ();
 DECAPx2_ASAP7_75t_R FILLER_216_522 ();
 DECAPx6_ASAP7_75t_R FILLER_216_534 ();
 FILLER_ASAP7_75t_R FILLER_216_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_550 ();
 DECAPx1_ASAP7_75t_R FILLER_216_570 ();
 DECAPx2_ASAP7_75t_R FILLER_216_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_614 ();
 DECAPx2_ASAP7_75t_R FILLER_216_623 ();
 FILLER_ASAP7_75t_R FILLER_216_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_631 ();
 DECAPx4_ASAP7_75t_R FILLER_216_634 ();
 FILLER_ASAP7_75t_R FILLER_216_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_646 ();
 DECAPx4_ASAP7_75t_R FILLER_216_665 ();
 DECAPx10_ASAP7_75t_R FILLER_216_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_703 ();
 DECAPx10_ASAP7_75t_R FILLER_216_712 ();
 DECAPx10_ASAP7_75t_R FILLER_216_734 ();
 DECAPx10_ASAP7_75t_R FILLER_216_756 ();
 DECAPx10_ASAP7_75t_R FILLER_216_778 ();
 DECAPx1_ASAP7_75t_R FILLER_216_800 ();
 DECAPx10_ASAP7_75t_R FILLER_216_822 ();
 DECAPx6_ASAP7_75t_R FILLER_216_852 ();
 DECAPx1_ASAP7_75t_R FILLER_216_866 ();
 DECAPx2_ASAP7_75t_R FILLER_216_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_905 ();
 DECAPx6_ASAP7_75t_R FILLER_216_918 ();
 DECAPx2_ASAP7_75t_R FILLER_216_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_938 ();
 DECAPx10_ASAP7_75t_R FILLER_216_945 ();
 FILLER_ASAP7_75t_R FILLER_216_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_969 ();
 DECAPx10_ASAP7_75t_R FILLER_216_979 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1001 ();
 FILLER_ASAP7_75t_R FILLER_216_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1043 ();
 FILLER_ASAP7_75t_R FILLER_216_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1091 ();
 FILLER_ASAP7_75t_R FILLER_216_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_217_172 ();
 FILLER_ASAP7_75t_R FILLER_217_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_193 ();
 DECAPx2_ASAP7_75t_R FILLER_217_197 ();
 FILLER_ASAP7_75t_R FILLER_217_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_205 ();
 DECAPx4_ASAP7_75t_R FILLER_217_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_224 ();
 DECAPx10_ASAP7_75t_R FILLER_217_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_263 ();
 DECAPx10_ASAP7_75t_R FILLER_217_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_301 ();
 FILLER_ASAP7_75t_R FILLER_217_322 ();
 DECAPx2_ASAP7_75t_R FILLER_217_331 ();
 DECAPx4_ASAP7_75t_R FILLER_217_351 ();
 FILLER_ASAP7_75t_R FILLER_217_361 ();
 DECAPx6_ASAP7_75t_R FILLER_217_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_390 ();
 DECAPx6_ASAP7_75t_R FILLER_217_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_411 ();
 DECAPx2_ASAP7_75t_R FILLER_217_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_428 ();
 DECAPx4_ASAP7_75t_R FILLER_217_440 ();
 FILLER_ASAP7_75t_R FILLER_217_450 ();
 DECAPx10_ASAP7_75t_R FILLER_217_458 ();
 DECAPx4_ASAP7_75t_R FILLER_217_480 ();
 FILLER_ASAP7_75t_R FILLER_217_490 ();
 FILLER_ASAP7_75t_R FILLER_217_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_502 ();
 FILLER_ASAP7_75t_R FILLER_217_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_529 ();
 FILLER_ASAP7_75t_R FILLER_217_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_592 ();
 DECAPx10_ASAP7_75t_R FILLER_217_599 ();
 DECAPx4_ASAP7_75t_R FILLER_217_621 ();
 FILLER_ASAP7_75t_R FILLER_217_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_633 ();
 DECAPx10_ASAP7_75t_R FILLER_217_655 ();
 DECAPx10_ASAP7_75t_R FILLER_217_677 ();
 DECAPx10_ASAP7_75t_R FILLER_217_699 ();
 DECAPx10_ASAP7_75t_R FILLER_217_721 ();
 DECAPx10_ASAP7_75t_R FILLER_217_743 ();
 DECAPx4_ASAP7_75t_R FILLER_217_765 ();
 DECAPx4_ASAP7_75t_R FILLER_217_787 ();
 DECAPx10_ASAP7_75t_R FILLER_217_803 ();
 DECAPx10_ASAP7_75t_R FILLER_217_825 ();
 DECAPx10_ASAP7_75t_R FILLER_217_847 ();
 DECAPx2_ASAP7_75t_R FILLER_217_869 ();
 FILLER_ASAP7_75t_R FILLER_217_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_877 ();
 DECAPx10_ASAP7_75t_R FILLER_217_884 ();
 DECAPx6_ASAP7_75t_R FILLER_217_906 ();
 DECAPx1_ASAP7_75t_R FILLER_217_920 ();
 DECAPx6_ASAP7_75t_R FILLER_217_930 ();
 DECAPx1_ASAP7_75t_R FILLER_217_944 ();
 DECAPx10_ASAP7_75t_R FILLER_217_954 ();
 DECAPx10_ASAP7_75t_R FILLER_217_976 ();
 DECAPx10_ASAP7_75t_R FILLER_217_998 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1036 ();
 FILLER_ASAP7_75t_R FILLER_217_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1070 ();
 FILLER_ASAP7_75t_R FILLER_217_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_217_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1170 ();
 DECAPx4_ASAP7_75t_R FILLER_217_1179 ();
 FILLER_ASAP7_75t_R FILLER_217_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_218_172 ();
 FILLER_ASAP7_75t_R FILLER_218_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_180 ();
 DECAPx10_ASAP7_75t_R FILLER_218_210 ();
 DECAPx10_ASAP7_75t_R FILLER_218_232 ();
 DECAPx6_ASAP7_75t_R FILLER_218_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_268 ();
 DECAPx10_ASAP7_75t_R FILLER_218_272 ();
 DECAPx6_ASAP7_75t_R FILLER_218_294 ();
 FILLER_ASAP7_75t_R FILLER_218_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_310 ();
 FILLER_ASAP7_75t_R FILLER_218_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_329 ();
 DECAPx4_ASAP7_75t_R FILLER_218_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_359 ();
 FILLER_ASAP7_75t_R FILLER_218_368 ();
 FILLER_ASAP7_75t_R FILLER_218_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_378 ();
 FILLER_ASAP7_75t_R FILLER_218_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_388 ();
 FILLER_ASAP7_75t_R FILLER_218_396 ();
 DECAPx10_ASAP7_75t_R FILLER_218_405 ();
 DECAPx1_ASAP7_75t_R FILLER_218_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_431 ();
 DECAPx1_ASAP7_75t_R FILLER_218_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_449 ();
 DECAPx1_ASAP7_75t_R FILLER_218_460 ();
 DECAPx6_ASAP7_75t_R FILLER_218_474 ();
 DECAPx1_ASAP7_75t_R FILLER_218_488 ();
 DECAPx10_ASAP7_75t_R FILLER_218_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_524 ();
 DECAPx6_ASAP7_75t_R FILLER_218_576 ();
 FILLER_ASAP7_75t_R FILLER_218_590 ();
 DECAPx6_ASAP7_75t_R FILLER_218_613 ();
 DECAPx1_ASAP7_75t_R FILLER_218_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_631 ();
 DECAPx10_ASAP7_75t_R FILLER_218_634 ();
 DECAPx10_ASAP7_75t_R FILLER_218_656 ();
 DECAPx10_ASAP7_75t_R FILLER_218_678 ();
 DECAPx10_ASAP7_75t_R FILLER_218_700 ();
 DECAPx10_ASAP7_75t_R FILLER_218_722 ();
 DECAPx10_ASAP7_75t_R FILLER_218_744 ();
 DECAPx4_ASAP7_75t_R FILLER_218_766 ();
 DECAPx10_ASAP7_75t_R FILLER_218_786 ();
 DECAPx10_ASAP7_75t_R FILLER_218_808 ();
 DECAPx6_ASAP7_75t_R FILLER_218_830 ();
 DECAPx10_ASAP7_75t_R FILLER_218_880 ();
 DECAPx6_ASAP7_75t_R FILLER_218_902 ();
 DECAPx1_ASAP7_75t_R FILLER_218_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_920 ();
 DECAPx10_ASAP7_75t_R FILLER_218_933 ();
 DECAPx4_ASAP7_75t_R FILLER_218_955 ();
 FILLER_ASAP7_75t_R FILLER_218_965 ();
 DECAPx1_ASAP7_75t_R FILLER_218_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_982 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_218_1029 ();
 FILLER_ASAP7_75t_R FILLER_218_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1142 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1186 ();
 FILLER_ASAP7_75t_R FILLER_218_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1276 ();
 FILLER_ASAP7_75t_R FILLER_218_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_219_172 ();
 DECAPx2_ASAP7_75t_R FILLER_219_194 ();
 FILLER_ASAP7_75t_R FILLER_219_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_202 ();
 DECAPx6_ASAP7_75t_R FILLER_219_215 ();
 DECAPx2_ASAP7_75t_R FILLER_219_237 ();
 FILLER_ASAP7_75t_R FILLER_219_243 ();
 DECAPx10_ASAP7_75t_R FILLER_219_274 ();
 DECAPx10_ASAP7_75t_R FILLER_219_296 ();
 DECAPx2_ASAP7_75t_R FILLER_219_318 ();
 FILLER_ASAP7_75t_R FILLER_219_324 ();
 DECAPx10_ASAP7_75t_R FILLER_219_334 ();
 DECAPx1_ASAP7_75t_R FILLER_219_356 ();
 DECAPx2_ASAP7_75t_R FILLER_219_366 ();
 FILLER_ASAP7_75t_R FILLER_219_372 ();
 DECAPx10_ASAP7_75t_R FILLER_219_386 ();
 FILLER_ASAP7_75t_R FILLER_219_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_424 ();
 DECAPx2_ASAP7_75t_R FILLER_219_435 ();
 DECAPx2_ASAP7_75t_R FILLER_219_447 ();
 DECAPx1_ASAP7_75t_R FILLER_219_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_465 ();
 DECAPx6_ASAP7_75t_R FILLER_219_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_487 ();
 DECAPx10_ASAP7_75t_R FILLER_219_495 ();
 DECAPx6_ASAP7_75t_R FILLER_219_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_531 ();
 DECAPx1_ASAP7_75t_R FILLER_219_542 ();
 DECAPx10_ASAP7_75t_R FILLER_219_576 ();
 DECAPx10_ASAP7_75t_R FILLER_219_598 ();
 DECAPx10_ASAP7_75t_R FILLER_219_620 ();
 DECAPx1_ASAP7_75t_R FILLER_219_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_646 ();
 DECAPx1_ASAP7_75t_R FILLER_219_655 ();
 DECAPx10_ASAP7_75t_R FILLER_219_665 ();
 DECAPx10_ASAP7_75t_R FILLER_219_687 ();
 DECAPx6_ASAP7_75t_R FILLER_219_709 ();
 FILLER_ASAP7_75t_R FILLER_219_723 ();
 DECAPx4_ASAP7_75t_R FILLER_219_740 ();
 FILLER_ASAP7_75t_R FILLER_219_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_752 ();
 DECAPx10_ASAP7_75t_R FILLER_219_765 ();
 DECAPx10_ASAP7_75t_R FILLER_219_787 ();
 DECAPx10_ASAP7_75t_R FILLER_219_809 ();
 FILLER_ASAP7_75t_R FILLER_219_831 ();
 DECAPx2_ASAP7_75t_R FILLER_219_844 ();
 FILLER_ASAP7_75t_R FILLER_219_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_852 ();
 DECAPx2_ASAP7_75t_R FILLER_219_863 ();
 DECAPx10_ASAP7_75t_R FILLER_219_876 ();
 FILLER_ASAP7_75t_R FILLER_219_898 ();
 DECAPx10_ASAP7_75t_R FILLER_219_903 ();
 DECAPx10_ASAP7_75t_R FILLER_219_925 ();
 DECAPx4_ASAP7_75t_R FILLER_219_947 ();
 DECAPx2_ASAP7_75t_R FILLER_219_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_984 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_219_1047 ();
 FILLER_ASAP7_75t_R FILLER_219_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_219_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_219_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_219_1170 ();
 FILLER_ASAP7_75t_R FILLER_219_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_219_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_220_172 ();
 DECAPx2_ASAP7_75t_R FILLER_220_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_200 ();
 DECAPx10_ASAP7_75t_R FILLER_220_209 ();
 DECAPx6_ASAP7_75t_R FILLER_220_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_245 ();
 FILLER_ASAP7_75t_R FILLER_220_252 ();
 DECAPx2_ASAP7_75t_R FILLER_220_260 ();
 FILLER_ASAP7_75t_R FILLER_220_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_268 ();
 DECAPx2_ASAP7_75t_R FILLER_220_277 ();
 FILLER_ASAP7_75t_R FILLER_220_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_285 ();
 DECAPx6_ASAP7_75t_R FILLER_220_294 ();
 DECAPx2_ASAP7_75t_R FILLER_220_308 ();
 DECAPx4_ASAP7_75t_R FILLER_220_332 ();
 FILLER_ASAP7_75t_R FILLER_220_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_344 ();
 DECAPx2_ASAP7_75t_R FILLER_220_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_359 ();
 DECAPx2_ASAP7_75t_R FILLER_220_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_373 ();
 DECAPx10_ASAP7_75t_R FILLER_220_380 ();
 DECAPx1_ASAP7_75t_R FILLER_220_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_406 ();
 DECAPx6_ASAP7_75t_R FILLER_220_417 ();
 FILLER_ASAP7_75t_R FILLER_220_431 ();
 DECAPx6_ASAP7_75t_R FILLER_220_449 ();
 FILLER_ASAP7_75t_R FILLER_220_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_465 ();
 FILLER_ASAP7_75t_R FILLER_220_472 ();
 DECAPx6_ASAP7_75t_R FILLER_220_498 ();
 DECAPx1_ASAP7_75t_R FILLER_220_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_516 ();
 DECAPx10_ASAP7_75t_R FILLER_220_525 ();
 DECAPx1_ASAP7_75t_R FILLER_220_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_551 ();
 DECAPx10_ASAP7_75t_R FILLER_220_560 ();
 DECAPx6_ASAP7_75t_R FILLER_220_582 ();
 DECAPx6_ASAP7_75t_R FILLER_220_610 ();
 DECAPx2_ASAP7_75t_R FILLER_220_634 ();
 DECAPx6_ASAP7_75t_R FILLER_220_670 ();
 DECAPx1_ASAP7_75t_R FILLER_220_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_701 ();
 DECAPx6_ASAP7_75t_R FILLER_220_712 ();
 DECAPx2_ASAP7_75t_R FILLER_220_729 ();
 DECAPx6_ASAP7_75t_R FILLER_220_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_755 ();
 DECAPx10_ASAP7_75t_R FILLER_220_768 ();
 FILLER_ASAP7_75t_R FILLER_220_790 ();
 FILLER_ASAP7_75t_R FILLER_220_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_807 ();
 DECAPx4_ASAP7_75t_R FILLER_220_814 ();
 FILLER_ASAP7_75t_R FILLER_220_824 ();
 DECAPx10_ASAP7_75t_R FILLER_220_847 ();
 FILLER_ASAP7_75t_R FILLER_220_869 ();
 FILLER_ASAP7_75t_R FILLER_220_910 ();
 DECAPx6_ASAP7_75t_R FILLER_220_919 ();
 FILLER_ASAP7_75t_R FILLER_220_933 ();
 DECAPx6_ASAP7_75t_R FILLER_220_946 ();
 FILLER_ASAP7_75t_R FILLER_220_960 ();
 DECAPx10_ASAP7_75t_R FILLER_220_969 ();
 DECAPx2_ASAP7_75t_R FILLER_220_998 ();
 FILLER_ASAP7_75t_R FILLER_220_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1079 ();
 FILLER_ASAP7_75t_R FILLER_220_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1111 ();
 FILLER_ASAP7_75t_R FILLER_220_1117 ();
 FILLER_ASAP7_75t_R FILLER_220_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_221_172 ();
 DECAPx2_ASAP7_75t_R FILLER_221_194 ();
 FILLER_ASAP7_75t_R FILLER_221_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_239 ();
 FILLER_ASAP7_75t_R FILLER_221_246 ();
 DECAPx6_ASAP7_75t_R FILLER_221_257 ();
 DECAPx2_ASAP7_75t_R FILLER_221_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_277 ();
 DECAPx6_ASAP7_75t_R FILLER_221_288 ();
 DECAPx1_ASAP7_75t_R FILLER_221_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_318 ();
 DECAPx10_ASAP7_75t_R FILLER_221_331 ();
 DECAPx2_ASAP7_75t_R FILLER_221_353 ();
 FILLER_ASAP7_75t_R FILLER_221_359 ();
 DECAPx1_ASAP7_75t_R FILLER_221_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_371 ();
 DECAPx6_ASAP7_75t_R FILLER_221_382 ();
 DECAPx2_ASAP7_75t_R FILLER_221_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_402 ();
 DECAPx2_ASAP7_75t_R FILLER_221_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_415 ();
 DECAPx2_ASAP7_75t_R FILLER_221_423 ();
 FILLER_ASAP7_75t_R FILLER_221_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_431 ();
 DECAPx10_ASAP7_75t_R FILLER_221_438 ();
 DECAPx4_ASAP7_75t_R FILLER_221_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_487 ();
 DECAPx6_ASAP7_75t_R FILLER_221_498 ();
 DECAPx1_ASAP7_75t_R FILLER_221_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_516 ();
 FILLER_ASAP7_75t_R FILLER_221_525 ();
 DECAPx2_ASAP7_75t_R FILLER_221_535 ();
 FILLER_ASAP7_75t_R FILLER_221_541 ();
 DECAPx2_ASAP7_75t_R FILLER_221_568 ();
 FILLER_ASAP7_75t_R FILLER_221_574 ();
 FILLER_ASAP7_75t_R FILLER_221_582 ();
 DECAPx1_ASAP7_75t_R FILLER_221_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_596 ();
 DECAPx4_ASAP7_75t_R FILLER_221_618 ();
 FILLER_ASAP7_75t_R FILLER_221_628 ();
 DECAPx4_ASAP7_75t_R FILLER_221_638 ();
 DECAPx4_ASAP7_75t_R FILLER_221_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_666 ();
 DECAPx4_ASAP7_75t_R FILLER_221_673 ();
 FILLER_ASAP7_75t_R FILLER_221_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_685 ();
 DECAPx2_ASAP7_75t_R FILLER_221_692 ();
 DECAPx6_ASAP7_75t_R FILLER_221_710 ();
 FILLER_ASAP7_75t_R FILLER_221_724 ();
 DECAPx10_ASAP7_75t_R FILLER_221_736 ();
 DECAPx10_ASAP7_75t_R FILLER_221_758 ();
 DECAPx6_ASAP7_75t_R FILLER_221_780 ();
 DECAPx10_ASAP7_75t_R FILLER_221_817 ();
 DECAPx10_ASAP7_75t_R FILLER_221_839 ();
 DECAPx4_ASAP7_75t_R FILLER_221_861 ();
 FILLER_ASAP7_75t_R FILLER_221_871 ();
 DECAPx10_ASAP7_75t_R FILLER_221_893 ();
 DECAPx4_ASAP7_75t_R FILLER_221_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_925 ();
 DECAPx10_ASAP7_75t_R FILLER_221_947 ();
 FILLER_ASAP7_75t_R FILLER_221_969 ();
 DECAPx10_ASAP7_75t_R FILLER_221_978 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1000 ();
 FILLER_ASAP7_75t_R FILLER_221_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1034 ();
 FILLER_ASAP7_75t_R FILLER_221_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1118 ();
 FILLER_ASAP7_75t_R FILLER_221_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1129 ();
 FILLER_ASAP7_75t_R FILLER_221_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1279 ();
 DECAPx6_ASAP7_75t_R FILLER_222_172 ();
 DECAPx2_ASAP7_75t_R FILLER_222_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_229 ();
 DECAPx10_ASAP7_75t_R FILLER_222_238 ();
 DECAPx10_ASAP7_75t_R FILLER_222_260 ();
 FILLER_ASAP7_75t_R FILLER_222_282 ();
 DECAPx6_ASAP7_75t_R FILLER_222_304 ();
 FILLER_ASAP7_75t_R FILLER_222_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_320 ();
 DECAPx2_ASAP7_75t_R FILLER_222_340 ();
 DECAPx2_ASAP7_75t_R FILLER_222_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_370 ();
 DECAPx1_ASAP7_75t_R FILLER_222_400 ();
 DECAPx2_ASAP7_75t_R FILLER_222_425 ();
 FILLER_ASAP7_75t_R FILLER_222_437 ();
 DECAPx2_ASAP7_75t_R FILLER_222_447 ();
 DECAPx4_ASAP7_75t_R FILLER_222_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_469 ();
 DECAPx1_ASAP7_75t_R FILLER_222_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_480 ();
 DECAPx2_ASAP7_75t_R FILLER_222_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_494 ();
 DECAPx6_ASAP7_75t_R FILLER_222_505 ();
 DECAPx2_ASAP7_75t_R FILLER_222_519 ();
 DECAPx6_ASAP7_75t_R FILLER_222_533 ();
 DECAPx1_ASAP7_75t_R FILLER_222_547 ();
 DECAPx4_ASAP7_75t_R FILLER_222_572 ();
 DECAPx4_ASAP7_75t_R FILLER_222_603 ();
 DECAPx2_ASAP7_75t_R FILLER_222_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_631 ();
 DECAPx10_ASAP7_75t_R FILLER_222_634 ();
 DECAPx10_ASAP7_75t_R FILLER_222_656 ();
 DECAPx10_ASAP7_75t_R FILLER_222_678 ();
 DECAPx6_ASAP7_75t_R FILLER_222_700 ();
 DECAPx2_ASAP7_75t_R FILLER_222_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_720 ();
 DECAPx10_ASAP7_75t_R FILLER_222_729 ();
 DECAPx2_ASAP7_75t_R FILLER_222_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_757 ();
 DECAPx10_ASAP7_75t_R FILLER_222_764 ();
 DECAPx10_ASAP7_75t_R FILLER_222_786 ();
 DECAPx10_ASAP7_75t_R FILLER_222_808 ();
 DECAPx2_ASAP7_75t_R FILLER_222_830 ();
 FILLER_ASAP7_75t_R FILLER_222_836 ();
 DECAPx2_ASAP7_75t_R FILLER_222_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_855 ();
 DECAPx10_ASAP7_75t_R FILLER_222_867 ();
 DECAPx10_ASAP7_75t_R FILLER_222_889 ();
 FILLER_ASAP7_75t_R FILLER_222_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_913 ();
 DECAPx2_ASAP7_75t_R FILLER_222_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_930 ();
 DECAPx1_ASAP7_75t_R FILLER_222_938 ();
 DECAPx6_ASAP7_75t_R FILLER_222_957 ();
 DECAPx1_ASAP7_75t_R FILLER_222_971 ();
 DECAPx1_ASAP7_75t_R FILLER_222_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_998 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_222_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1167 ();
 FILLER_ASAP7_75t_R FILLER_222_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_223_172 ();
 FILLER_ASAP7_75t_R FILLER_223_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_218 ();
 DECAPx10_ASAP7_75t_R FILLER_223_231 ();
 DECAPx10_ASAP7_75t_R FILLER_223_253 ();
 DECAPx2_ASAP7_75t_R FILLER_223_275 ();
 FILLER_ASAP7_75t_R FILLER_223_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_283 ();
 DECAPx4_ASAP7_75t_R FILLER_223_290 ();
 FILLER_ASAP7_75t_R FILLER_223_300 ();
 DECAPx6_ASAP7_75t_R FILLER_223_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_373 ();
 DECAPx10_ASAP7_75t_R FILLER_223_380 ();
 DECAPx4_ASAP7_75t_R FILLER_223_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_419 ();
 FILLER_ASAP7_75t_R FILLER_223_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_429 ();
 FILLER_ASAP7_75t_R FILLER_223_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_440 ();
 DECAPx4_ASAP7_75t_R FILLER_223_447 ();
 DECAPx2_ASAP7_75t_R FILLER_223_475 ();
 DECAPx10_ASAP7_75t_R FILLER_223_489 ();
 DECAPx10_ASAP7_75t_R FILLER_223_511 ();
 DECAPx10_ASAP7_75t_R FILLER_223_533 ();
 FILLER_ASAP7_75t_R FILLER_223_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_557 ();
 DECAPx10_ASAP7_75t_R FILLER_223_572 ();
 DECAPx10_ASAP7_75t_R FILLER_223_594 ();
 DECAPx10_ASAP7_75t_R FILLER_223_616 ();
 DECAPx2_ASAP7_75t_R FILLER_223_638 ();
 FILLER_ASAP7_75t_R FILLER_223_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_652 ();
 DECAPx1_ASAP7_75t_R FILLER_223_659 ();
 FILLER_ASAP7_75t_R FILLER_223_669 ();
 DECAPx10_ASAP7_75t_R FILLER_223_687 ();
 DECAPx10_ASAP7_75t_R FILLER_223_709 ();
 DECAPx10_ASAP7_75t_R FILLER_223_731 ();
 DECAPx10_ASAP7_75t_R FILLER_223_753 ();
 DECAPx1_ASAP7_75t_R FILLER_223_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_779 ();
 DECAPx10_ASAP7_75t_R FILLER_223_786 ();
 DECAPx10_ASAP7_75t_R FILLER_223_808 ();
 FILLER_ASAP7_75t_R FILLER_223_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_832 ();
 DECAPx10_ASAP7_75t_R FILLER_223_875 ();
 DECAPx6_ASAP7_75t_R FILLER_223_897 ();
 DECAPx1_ASAP7_75t_R FILLER_223_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_915 ();
 DECAPx6_ASAP7_75t_R FILLER_223_924 ();
 DECAPx1_ASAP7_75t_R FILLER_223_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_942 ();
 DECAPx4_ASAP7_75t_R FILLER_223_985 ();
 FILLER_ASAP7_75t_R FILLER_223_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_223_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1166 ();
 FILLER_ASAP7_75t_R FILLER_223_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_223_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_224_172 ();
 DECAPx2_ASAP7_75t_R FILLER_224_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_192 ();
 DECAPx6_ASAP7_75t_R FILLER_224_213 ();
 FILLER_ASAP7_75t_R FILLER_224_241 ();
 DECAPx6_ASAP7_75t_R FILLER_224_269 ();
 DECAPx1_ASAP7_75t_R FILLER_224_283 ();
 DECAPx6_ASAP7_75t_R FILLER_224_298 ();
 FILLER_ASAP7_75t_R FILLER_224_312 ();
 DECAPx10_ASAP7_75t_R FILLER_224_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_342 ();
 DECAPx2_ASAP7_75t_R FILLER_224_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_355 ();
 DECAPx1_ASAP7_75t_R FILLER_224_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_368 ();
 DECAPx10_ASAP7_75t_R FILLER_224_375 ();
 DECAPx10_ASAP7_75t_R FILLER_224_397 ();
 DECAPx6_ASAP7_75t_R FILLER_224_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_433 ();
 DECAPx6_ASAP7_75t_R FILLER_224_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_456 ();
 DECAPx10_ASAP7_75t_R FILLER_224_469 ();
 DECAPx6_ASAP7_75t_R FILLER_224_491 ();
 FILLER_ASAP7_75t_R FILLER_224_505 ();
 DECAPx10_ASAP7_75t_R FILLER_224_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_539 ();
 DECAPx2_ASAP7_75t_R FILLER_224_546 ();
 FILLER_ASAP7_75t_R FILLER_224_552 ();
 DECAPx10_ASAP7_75t_R FILLER_224_562 ();
 DECAPx10_ASAP7_75t_R FILLER_224_584 ();
 DECAPx2_ASAP7_75t_R FILLER_224_606 ();
 FILLER_ASAP7_75t_R FILLER_224_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_614 ();
 DECAPx2_ASAP7_75t_R FILLER_224_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_651 ();
 DECAPx10_ASAP7_75t_R FILLER_224_668 ();
 DECAPx2_ASAP7_75t_R FILLER_224_690 ();
 FILLER_ASAP7_75t_R FILLER_224_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_698 ();
 DECAPx6_ASAP7_75t_R FILLER_224_709 ();
 DECAPx2_ASAP7_75t_R FILLER_224_723 ();
 DECAPx10_ASAP7_75t_R FILLER_224_735 ();
 DECAPx10_ASAP7_75t_R FILLER_224_757 ();
 DECAPx10_ASAP7_75t_R FILLER_224_779 ();
 DECAPx4_ASAP7_75t_R FILLER_224_801 ();
 FILLER_ASAP7_75t_R FILLER_224_811 ();
 DECAPx2_ASAP7_75t_R FILLER_224_825 ();
 FILLER_ASAP7_75t_R FILLER_224_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_833 ();
 DECAPx10_ASAP7_75t_R FILLER_224_840 ();
 DECAPx10_ASAP7_75t_R FILLER_224_862 ();
 DECAPx2_ASAP7_75t_R FILLER_224_898 ();
 FILLER_ASAP7_75t_R FILLER_224_904 ();
 DECAPx10_ASAP7_75t_R FILLER_224_930 ();
 FILLER_ASAP7_75t_R FILLER_224_952 ();
 DECAPx10_ASAP7_75t_R FILLER_224_957 ();
 DECAPx2_ASAP7_75t_R FILLER_224_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1014 ();
 FILLER_ASAP7_75t_R FILLER_224_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1037 ();
 FILLER_ASAP7_75t_R FILLER_224_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_224_1105 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1112 ();
 FILLER_ASAP7_75t_R FILLER_224_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1168 ();
 FILLER_ASAP7_75t_R FILLER_224_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1284 ();
 FILLER_ASAP7_75t_R FILLER_224_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_225_172 ();
 FILLER_ASAP7_75t_R FILLER_225_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_196 ();
 DECAPx1_ASAP7_75t_R FILLER_225_214 ();
 DECAPx4_ASAP7_75t_R FILLER_225_230 ();
 FILLER_ASAP7_75t_R FILLER_225_240 ();
 DECAPx2_ASAP7_75t_R FILLER_225_248 ();
 DECAPx10_ASAP7_75t_R FILLER_225_261 ();
 DECAPx2_ASAP7_75t_R FILLER_225_283 ();
 FILLER_ASAP7_75t_R FILLER_225_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_291 ();
 DECAPx6_ASAP7_75t_R FILLER_225_302 ();
 FILLER_ASAP7_75t_R FILLER_225_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_318 ();
 DECAPx1_ASAP7_75t_R FILLER_225_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_333 ();
 DECAPx1_ASAP7_75t_R FILLER_225_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_344 ();
 DECAPx10_ASAP7_75t_R FILLER_225_354 ();
 DECAPx2_ASAP7_75t_R FILLER_225_376 ();
 DECAPx6_ASAP7_75t_R FILLER_225_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_402 ();
 DECAPx6_ASAP7_75t_R FILLER_225_409 ();
 FILLER_ASAP7_75t_R FILLER_225_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_425 ();
 DECAPx10_ASAP7_75t_R FILLER_225_434 ();
 DECAPx2_ASAP7_75t_R FILLER_225_456 ();
 FILLER_ASAP7_75t_R FILLER_225_462 ();
 DECAPx2_ASAP7_75t_R FILLER_225_482 ();
 FILLER_ASAP7_75t_R FILLER_225_488 ();
 DECAPx10_ASAP7_75t_R FILLER_225_497 ();
 DECAPx10_ASAP7_75t_R FILLER_225_519 ();
 FILLER_ASAP7_75t_R FILLER_225_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_551 ();
 DECAPx2_ASAP7_75t_R FILLER_225_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_561 ();
 DECAPx10_ASAP7_75t_R FILLER_225_573 ();
 DECAPx2_ASAP7_75t_R FILLER_225_603 ();
 DECAPx10_ASAP7_75t_R FILLER_225_639 ();
 DECAPx10_ASAP7_75t_R FILLER_225_661 ();
 DECAPx4_ASAP7_75t_R FILLER_225_683 ();
 FILLER_ASAP7_75t_R FILLER_225_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_695 ();
 FILLER_ASAP7_75t_R FILLER_225_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_708 ();
 DECAPx6_ASAP7_75t_R FILLER_225_733 ();
 FILLER_ASAP7_75t_R FILLER_225_747 ();
 DECAPx4_ASAP7_75t_R FILLER_225_755 ();
 FILLER_ASAP7_75t_R FILLER_225_765 ();
 DECAPx1_ASAP7_75t_R FILLER_225_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_777 ();
 DECAPx10_ASAP7_75t_R FILLER_225_784 ();
 DECAPx10_ASAP7_75t_R FILLER_225_806 ();
 FILLER_ASAP7_75t_R FILLER_225_828 ();
 DECAPx10_ASAP7_75t_R FILLER_225_836 ();
 DECAPx6_ASAP7_75t_R FILLER_225_858 ();
 FILLER_ASAP7_75t_R FILLER_225_872 ();
 FILLER_ASAP7_75t_R FILLER_225_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_888 ();
 DECAPx10_ASAP7_75t_R FILLER_225_910 ();
 DECAPx10_ASAP7_75t_R FILLER_225_932 ();
 DECAPx6_ASAP7_75t_R FILLER_225_954 ();
 DECAPx1_ASAP7_75t_R FILLER_225_968 ();
 DECAPx10_ASAP7_75t_R FILLER_225_975 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1051 ();
 FILLER_ASAP7_75t_R FILLER_225_1061 ();
 FILLER_ASAP7_75t_R FILLER_225_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1098 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1120 ();
 FILLER_ASAP7_75t_R FILLER_225_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_225_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_226_172 ();
 DECAPx2_ASAP7_75t_R FILLER_226_194 ();
 DECAPx4_ASAP7_75t_R FILLER_226_230 ();
 FILLER_ASAP7_75t_R FILLER_226_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_242 ();
 DECAPx4_ASAP7_75t_R FILLER_226_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_263 ();
 DECAPx2_ASAP7_75t_R FILLER_226_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_280 ();
 DECAPx2_ASAP7_75t_R FILLER_226_297 ();
 FILLER_ASAP7_75t_R FILLER_226_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_305 ();
 DECAPx10_ASAP7_75t_R FILLER_226_318 ();
 DECAPx10_ASAP7_75t_R FILLER_226_340 ();
 DECAPx10_ASAP7_75t_R FILLER_226_362 ();
 DECAPx6_ASAP7_75t_R FILLER_226_384 ();
 DECAPx2_ASAP7_75t_R FILLER_226_398 ();
 DECAPx1_ASAP7_75t_R FILLER_226_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_414 ();
 DECAPx10_ASAP7_75t_R FILLER_226_429 ();
 DECAPx1_ASAP7_75t_R FILLER_226_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_455 ();
 FILLER_ASAP7_75t_R FILLER_226_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_464 ();
 DECAPx4_ASAP7_75t_R FILLER_226_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_504 ();
 DECAPx6_ASAP7_75t_R FILLER_226_516 ();
 DECAPx2_ASAP7_75t_R FILLER_226_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_536 ();
 DECAPx4_ASAP7_75t_R FILLER_226_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_631 ();
 DECAPx4_ASAP7_75t_R FILLER_226_634 ();
 FILLER_ASAP7_75t_R FILLER_226_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_646 ();
 DECAPx10_ASAP7_75t_R FILLER_226_657 ();
 DECAPx2_ASAP7_75t_R FILLER_226_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_685 ();
 DECAPx10_ASAP7_75t_R FILLER_226_704 ();
 DECAPx10_ASAP7_75t_R FILLER_226_726 ();
 DECAPx1_ASAP7_75t_R FILLER_226_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_752 ();
 DECAPx2_ASAP7_75t_R FILLER_226_763 ();
 DECAPx1_ASAP7_75t_R FILLER_226_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_789 ();
 FILLER_ASAP7_75t_R FILLER_226_800 ();
 DECAPx10_ASAP7_75t_R FILLER_226_810 ();
 DECAPx10_ASAP7_75t_R FILLER_226_832 ();
 DECAPx10_ASAP7_75t_R FILLER_226_854 ();
 DECAPx10_ASAP7_75t_R FILLER_226_876 ();
 DECAPx6_ASAP7_75t_R FILLER_226_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_912 ();
 DECAPx1_ASAP7_75t_R FILLER_226_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_941 ();
 DECAPx2_ASAP7_75t_R FILLER_226_950 ();
 FILLER_ASAP7_75t_R FILLER_226_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_958 ();
 FILLER_ASAP7_75t_R FILLER_226_980 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1077 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1081 ();
 FILLER_ASAP7_75t_R FILLER_226_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_226_1123 ();
 FILLER_ASAP7_75t_R FILLER_226_1129 ();
 FILLER_ASAP7_75t_R FILLER_226_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1160 ();
 FILLER_ASAP7_75t_R FILLER_226_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1276 ();
 FILLER_ASAP7_75t_R FILLER_226_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_227_172 ();
 FILLER_ASAP7_75t_R FILLER_227_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_196 ();
 DECAPx2_ASAP7_75t_R FILLER_227_218 ();
 FILLER_ASAP7_75t_R FILLER_227_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_226 ();
 DECAPx1_ASAP7_75t_R FILLER_227_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_238 ();
 FILLER_ASAP7_75t_R FILLER_227_248 ();
 DECAPx10_ASAP7_75t_R FILLER_227_256 ();
 DECAPx4_ASAP7_75t_R FILLER_227_278 ();
 FILLER_ASAP7_75t_R FILLER_227_288 ();
 FILLER_ASAP7_75t_R FILLER_227_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_307 ();
 DECAPx1_ASAP7_75t_R FILLER_227_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_318 ();
 FILLER_ASAP7_75t_R FILLER_227_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_327 ();
 DECAPx1_ASAP7_75t_R FILLER_227_334 ();
 DECAPx10_ASAP7_75t_R FILLER_227_344 ();
 DECAPx1_ASAP7_75t_R FILLER_227_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_384 ();
 DECAPx1_ASAP7_75t_R FILLER_227_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_397 ();
 DECAPx10_ASAP7_75t_R FILLER_227_438 ();
 DECAPx4_ASAP7_75t_R FILLER_227_460 ();
 FILLER_ASAP7_75t_R FILLER_227_470 ();
 FILLER_ASAP7_75t_R FILLER_227_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_480 ();
 DECAPx10_ASAP7_75t_R FILLER_227_489 ();
 DECAPx6_ASAP7_75t_R FILLER_227_511 ();
 DECAPx2_ASAP7_75t_R FILLER_227_533 ();
 FILLER_ASAP7_75t_R FILLER_227_539 ();
 FILLER_ASAP7_75t_R FILLER_227_549 ();
 DECAPx10_ASAP7_75t_R FILLER_227_565 ();
 DECAPx1_ASAP7_75t_R FILLER_227_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_591 ();
 DECAPx4_ASAP7_75t_R FILLER_227_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_608 ();
 DECAPx4_ASAP7_75t_R FILLER_227_639 ();
 FILLER_ASAP7_75t_R FILLER_227_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_651 ();
 FILLER_ASAP7_75t_R FILLER_227_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_662 ();
 DECAPx1_ASAP7_75t_R FILLER_227_671 ();
 DECAPx10_ASAP7_75t_R FILLER_227_685 ();
 DECAPx10_ASAP7_75t_R FILLER_227_707 ();
 DECAPx10_ASAP7_75t_R FILLER_227_729 ();
 DECAPx10_ASAP7_75t_R FILLER_227_751 ();
 DECAPx2_ASAP7_75t_R FILLER_227_773 ();
 DECAPx10_ASAP7_75t_R FILLER_227_785 ();
 DECAPx10_ASAP7_75t_R FILLER_227_807 ();
 DECAPx6_ASAP7_75t_R FILLER_227_829 ();
 FILLER_ASAP7_75t_R FILLER_227_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_845 ();
 FILLER_ASAP7_75t_R FILLER_227_866 ();
 DECAPx1_ASAP7_75t_R FILLER_227_874 ();
 DECAPx6_ASAP7_75t_R FILLER_227_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_898 ();
 DECAPx6_ASAP7_75t_R FILLER_227_913 ();
 FILLER_ASAP7_75t_R FILLER_227_927 ();
 FILLER_ASAP7_75t_R FILLER_227_958 ();
 DECAPx2_ASAP7_75t_R FILLER_227_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1016 ();
 FILLER_ASAP7_75t_R FILLER_227_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1079 ();
 FILLER_ASAP7_75t_R FILLER_227_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1118 ();
 FILLER_ASAP7_75t_R FILLER_227_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_227_1283 ();
 DECAPx6_ASAP7_75t_R FILLER_228_172 ();
 DECAPx1_ASAP7_75t_R FILLER_228_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_198 ();
 FILLER_ASAP7_75t_R FILLER_228_215 ();
 DECAPx4_ASAP7_75t_R FILLER_228_225 ();
 FILLER_ASAP7_75t_R FILLER_228_235 ();
 DECAPx6_ASAP7_75t_R FILLER_228_249 ();
 FILLER_ASAP7_75t_R FILLER_228_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_265 ();
 DECAPx6_ASAP7_75t_R FILLER_228_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_286 ();
 DECAPx4_ASAP7_75t_R FILLER_228_293 ();
 FILLER_ASAP7_75t_R FILLER_228_303 ();
 DECAPx4_ASAP7_75t_R FILLER_228_311 ();
 FILLER_ASAP7_75t_R FILLER_228_321 ();
 DECAPx4_ASAP7_75t_R FILLER_228_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_359 ();
 FILLER_ASAP7_75t_R FILLER_228_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_369 ();
 DECAPx2_ASAP7_75t_R FILLER_228_378 ();
 DECAPx10_ASAP7_75t_R FILLER_228_390 ();
 DECAPx4_ASAP7_75t_R FILLER_228_412 ();
 FILLER_ASAP7_75t_R FILLER_228_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_424 ();
 FILLER_ASAP7_75t_R FILLER_228_431 ();
 DECAPx4_ASAP7_75t_R FILLER_228_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_450 ();
 DECAPx4_ASAP7_75t_R FILLER_228_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_497 ();
 FILLER_ASAP7_75t_R FILLER_228_504 ();
 DECAPx10_ASAP7_75t_R FILLER_228_514 ();
 DECAPx10_ASAP7_75t_R FILLER_228_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_558 ();
 DECAPx2_ASAP7_75t_R FILLER_228_565 ();
 FILLER_ASAP7_75t_R FILLER_228_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_587 ();
 DECAPx6_ASAP7_75t_R FILLER_228_594 ();
 DECAPx1_ASAP7_75t_R FILLER_228_608 ();
 DECAPx2_ASAP7_75t_R FILLER_228_620 ();
 FILLER_ASAP7_75t_R FILLER_228_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_631 ();
 DECAPx2_ASAP7_75t_R FILLER_228_634 ();
 DECAPx2_ASAP7_75t_R FILLER_228_656 ();
 FILLER_ASAP7_75t_R FILLER_228_662 ();
 DECAPx10_ASAP7_75t_R FILLER_228_680 ();
 DECAPx10_ASAP7_75t_R FILLER_228_702 ();
 DECAPx10_ASAP7_75t_R FILLER_228_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_746 ();
 DECAPx4_ASAP7_75t_R FILLER_228_753 ();
 FILLER_ASAP7_75t_R FILLER_228_763 ();
 DECAPx4_ASAP7_75t_R FILLER_228_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_781 ();
 DECAPx10_ASAP7_75t_R FILLER_228_788 ();
 DECAPx10_ASAP7_75t_R FILLER_228_810 ();
 DECAPx4_ASAP7_75t_R FILLER_228_832 ();
 FILLER_ASAP7_75t_R FILLER_228_842 ();
 DECAPx2_ASAP7_75t_R FILLER_228_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_887 ();
 DECAPx6_ASAP7_75t_R FILLER_228_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_926 ();
 FILLER_ASAP7_75t_R FILLER_228_930 ();
 DECAPx1_ASAP7_75t_R FILLER_228_938 ();
 DECAPx4_ASAP7_75t_R FILLER_228_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_961 ();
 FILLER_ASAP7_75t_R FILLER_228_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_992 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1057 ();
 FILLER_ASAP7_75t_R FILLER_228_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_228_1084 ();
 FILLER_ASAP7_75t_R FILLER_228_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1099 ();
 FILLER_ASAP7_75t_R FILLER_228_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_228_1149 ();
 FILLER_ASAP7_75t_R FILLER_228_1159 ();
 FILLER_ASAP7_75t_R FILLER_228_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_229_172 ();
 DECAPx2_ASAP7_75t_R FILLER_229_194 ();
 FILLER_ASAP7_75t_R FILLER_229_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_202 ();
 DECAPx2_ASAP7_75t_R FILLER_229_212 ();
 DECAPx4_ASAP7_75t_R FILLER_229_230 ();
 FILLER_ASAP7_75t_R FILLER_229_240 ();
 DECAPx4_ASAP7_75t_R FILLER_229_251 ();
 FILLER_ASAP7_75t_R FILLER_229_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_263 ();
 DECAPx1_ASAP7_75t_R FILLER_229_274 ();
 DECAPx2_ASAP7_75t_R FILLER_229_291 ();
 FILLER_ASAP7_75t_R FILLER_229_297 ();
 DECAPx1_ASAP7_75t_R FILLER_229_311 ();
 DECAPx6_ASAP7_75t_R FILLER_229_322 ();
 DECAPx2_ASAP7_75t_R FILLER_229_336 ();
 DECAPx6_ASAP7_75t_R FILLER_229_348 ();
 FILLER_ASAP7_75t_R FILLER_229_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_374 ();
 DECAPx10_ASAP7_75t_R FILLER_229_383 ();
 DECAPx10_ASAP7_75t_R FILLER_229_405 ();
 DECAPx2_ASAP7_75t_R FILLER_229_427 ();
 FILLER_ASAP7_75t_R FILLER_229_433 ();
 DECAPx4_ASAP7_75t_R FILLER_229_451 ();
 FILLER_ASAP7_75t_R FILLER_229_461 ();
 FILLER_ASAP7_75t_R FILLER_229_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_472 ();
 DECAPx1_ASAP7_75t_R FILLER_229_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_493 ();
 DECAPx10_ASAP7_75t_R FILLER_229_502 ();
 DECAPx2_ASAP7_75t_R FILLER_229_524 ();
 FILLER_ASAP7_75t_R FILLER_229_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_532 ();
 DECAPx6_ASAP7_75t_R FILLER_229_539 ();
 FILLER_ASAP7_75t_R FILLER_229_553 ();
 DECAPx6_ASAP7_75t_R FILLER_229_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_583 ();
 DECAPx2_ASAP7_75t_R FILLER_229_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_598 ();
 FILLER_ASAP7_75t_R FILLER_229_602 ();
 DECAPx6_ASAP7_75t_R FILLER_229_625 ();
 DECAPx1_ASAP7_75t_R FILLER_229_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_643 ();
 DECAPx2_ASAP7_75t_R FILLER_229_660 ();
 FILLER_ASAP7_75t_R FILLER_229_666 ();
 DECAPx2_ASAP7_75t_R FILLER_229_674 ();
 FILLER_ASAP7_75t_R FILLER_229_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_682 ();
 DECAPx10_ASAP7_75t_R FILLER_229_690 ();
 DECAPx1_ASAP7_75t_R FILLER_229_712 ();
 DECAPx2_ASAP7_75t_R FILLER_229_728 ();
 DECAPx1_ASAP7_75t_R FILLER_229_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_744 ();
 DECAPx6_ASAP7_75t_R FILLER_229_751 ();
 DECAPx1_ASAP7_75t_R FILLER_229_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_769 ();
 DECAPx2_ASAP7_75t_R FILLER_229_776 ();
 DECAPx4_ASAP7_75t_R FILLER_229_792 ();
 FILLER_ASAP7_75t_R FILLER_229_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_804 ();
 DECAPx6_ASAP7_75t_R FILLER_229_815 ();
 FILLER_ASAP7_75t_R FILLER_229_829 ();
 DECAPx6_ASAP7_75t_R FILLER_229_848 ();
 DECAPx2_ASAP7_75t_R FILLER_229_862 ();
 DECAPx1_ASAP7_75t_R FILLER_229_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_878 ();
 DECAPx10_ASAP7_75t_R FILLER_229_885 ();
 FILLER_ASAP7_75t_R FILLER_229_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_909 ();
 DECAPx6_ASAP7_75t_R FILLER_229_939 ();
 FILLER_ASAP7_75t_R FILLER_229_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_955 ();
 DECAPx6_ASAP7_75t_R FILLER_229_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_973 ();
 DECAPx10_ASAP7_75t_R FILLER_229_982 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1096 ();
 FILLER_ASAP7_75t_R FILLER_229_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1129 ();
 FILLER_ASAP7_75t_R FILLER_229_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_230_172 ();
 DECAPx2_ASAP7_75t_R FILLER_230_194 ();
 FILLER_ASAP7_75t_R FILLER_230_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_214 ();
 DECAPx10_ASAP7_75t_R FILLER_230_224 ();
 DECAPx10_ASAP7_75t_R FILLER_230_246 ();
 DECAPx1_ASAP7_75t_R FILLER_230_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_278 ();
 FILLER_ASAP7_75t_R FILLER_230_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_287 ();
 DECAPx10_ASAP7_75t_R FILLER_230_294 ();
 DECAPx10_ASAP7_75t_R FILLER_230_316 ();
 DECAPx10_ASAP7_75t_R FILLER_230_338 ();
 DECAPx6_ASAP7_75t_R FILLER_230_360 ();
 DECAPx6_ASAP7_75t_R FILLER_230_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_391 ();
 DECAPx6_ASAP7_75t_R FILLER_230_416 ();
 DECAPx1_ASAP7_75t_R FILLER_230_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_442 ();
 DECAPx10_ASAP7_75t_R FILLER_230_449 ();
 DECAPx2_ASAP7_75t_R FILLER_230_471 ();
 DECAPx10_ASAP7_75t_R FILLER_230_493 ();
 DECAPx4_ASAP7_75t_R FILLER_230_515 ();
 FILLER_ASAP7_75t_R FILLER_230_525 ();
 FILLER_ASAP7_75t_R FILLER_230_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_547 ();
 DECAPx2_ASAP7_75t_R FILLER_230_551 ();
 FILLER_ASAP7_75t_R FILLER_230_557 ();
 DECAPx2_ASAP7_75t_R FILLER_230_570 ();
 FILLER_ASAP7_75t_R FILLER_230_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_578 ();
 DECAPx10_ASAP7_75t_R FILLER_230_600 ();
 DECAPx1_ASAP7_75t_R FILLER_230_622 ();
 FILLER_ASAP7_75t_R FILLER_230_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_631 ();
 DECAPx2_ASAP7_75t_R FILLER_230_634 ();
 FILLER_ASAP7_75t_R FILLER_230_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_642 ();
 DECAPx10_ASAP7_75t_R FILLER_230_649 ();
 DECAPx1_ASAP7_75t_R FILLER_230_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_675 ();
 DECAPx1_ASAP7_75t_R FILLER_230_688 ();
 DECAPx10_ASAP7_75t_R FILLER_230_704 ();
 DECAPx10_ASAP7_75t_R FILLER_230_726 ();
 DECAPx10_ASAP7_75t_R FILLER_230_748 ();
 DECAPx10_ASAP7_75t_R FILLER_230_770 ();
 DECAPx10_ASAP7_75t_R FILLER_230_792 ();
 DECAPx10_ASAP7_75t_R FILLER_230_814 ();
 DECAPx10_ASAP7_75t_R FILLER_230_836 ();
 DECAPx10_ASAP7_75t_R FILLER_230_858 ();
 DECAPx10_ASAP7_75t_R FILLER_230_880 ();
 DECAPx6_ASAP7_75t_R FILLER_230_902 ();
 DECAPx2_ASAP7_75t_R FILLER_230_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_922 ();
 DECAPx6_ASAP7_75t_R FILLER_230_929 ();
 DECAPx1_ASAP7_75t_R FILLER_230_943 ();
 FILLER_ASAP7_75t_R FILLER_230_961 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1069 ();
 DECAPx4_ASAP7_75t_R FILLER_230_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_230_1121 ();
 FILLER_ASAP7_75t_R FILLER_230_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1150 ();
 FILLER_ASAP7_75t_R FILLER_230_1156 ();
 FILLER_ASAP7_75t_R FILLER_230_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1268 ();
 FILLER_ASAP7_75t_R FILLER_230_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_231_172 ();
 DECAPx4_ASAP7_75t_R FILLER_231_194 ();
 FILLER_ASAP7_75t_R FILLER_231_204 ();
 DECAPx2_ASAP7_75t_R FILLER_231_226 ();
 FILLER_ASAP7_75t_R FILLER_231_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_234 ();
 FILLER_ASAP7_75t_R FILLER_231_247 ();
 DECAPx10_ASAP7_75t_R FILLER_231_252 ();
 DECAPx10_ASAP7_75t_R FILLER_231_274 ();
 DECAPx2_ASAP7_75t_R FILLER_231_296 ();
 FILLER_ASAP7_75t_R FILLER_231_302 ();
 DECAPx1_ASAP7_75t_R FILLER_231_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_316 ();
 DECAPx1_ASAP7_75t_R FILLER_231_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_327 ();
 DECAPx10_ASAP7_75t_R FILLER_231_335 ();
 DECAPx6_ASAP7_75t_R FILLER_231_357 ();
 DECAPx1_ASAP7_75t_R FILLER_231_371 ();
 DECAPx6_ASAP7_75t_R FILLER_231_389 ();
 DECAPx1_ASAP7_75t_R FILLER_231_403 ();
 FILLER_ASAP7_75t_R FILLER_231_410 ();
 DECAPx2_ASAP7_75t_R FILLER_231_420 ();
 FILLER_ASAP7_75t_R FILLER_231_426 ();
 DECAPx1_ASAP7_75t_R FILLER_231_440 ();
 DECAPx2_ASAP7_75t_R FILLER_231_453 ();
 DECAPx2_ASAP7_75t_R FILLER_231_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_481 ();
 DECAPx10_ASAP7_75t_R FILLER_231_489 ();
 DECAPx6_ASAP7_75t_R FILLER_231_511 ();
 DECAPx2_ASAP7_75t_R FILLER_231_525 ();
 DECAPx1_ASAP7_75t_R FILLER_231_552 ();
 DECAPx6_ASAP7_75t_R FILLER_231_577 ();
 DECAPx1_ASAP7_75t_R FILLER_231_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_595 ();
 FILLER_ASAP7_75t_R FILLER_231_606 ();
 DECAPx4_ASAP7_75t_R FILLER_231_616 ();
 DECAPx6_ASAP7_75t_R FILLER_231_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_675 ();
 DECAPx4_ASAP7_75t_R FILLER_231_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_692 ();
 DECAPx10_ASAP7_75t_R FILLER_231_699 ();
 DECAPx10_ASAP7_75t_R FILLER_231_721 ();
 DECAPx10_ASAP7_75t_R FILLER_231_743 ();
 DECAPx10_ASAP7_75t_R FILLER_231_765 ();
 DECAPx10_ASAP7_75t_R FILLER_231_787 ();
 DECAPx10_ASAP7_75t_R FILLER_231_809 ();
 DECAPx6_ASAP7_75t_R FILLER_231_831 ();
 FILLER_ASAP7_75t_R FILLER_231_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_847 ();
 DECAPx10_ASAP7_75t_R FILLER_231_865 ();
 DECAPx4_ASAP7_75t_R FILLER_231_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_897 ();
 DECAPx10_ASAP7_75t_R FILLER_231_907 ();
 DECAPx4_ASAP7_75t_R FILLER_231_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_939 ();
 DECAPx1_ASAP7_75t_R FILLER_231_943 ();
 DECAPx6_ASAP7_75t_R FILLER_231_968 ();
 DECAPx2_ASAP7_75t_R FILLER_231_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_988 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_231_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1031 ();
 FILLER_ASAP7_75t_R FILLER_231_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1086 ();
 FILLER_ASAP7_75t_R FILLER_231_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_231_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_232_172 ();
 DECAPx6_ASAP7_75t_R FILLER_232_194 ();
 DECAPx2_ASAP7_75t_R FILLER_232_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_214 ();
 DECAPx1_ASAP7_75t_R FILLER_232_221 ();
 DECAPx1_ASAP7_75t_R FILLER_232_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_245 ();
 DECAPx10_ASAP7_75t_R FILLER_232_255 ();
 FILLER_ASAP7_75t_R FILLER_232_277 ();
 DECAPx4_ASAP7_75t_R FILLER_232_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_302 ();
 FILLER_ASAP7_75t_R FILLER_232_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_323 ();
 DECAPx2_ASAP7_75t_R FILLER_232_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_347 ();
 FILLER_ASAP7_75t_R FILLER_232_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_377 ();
 DECAPx10_ASAP7_75t_R FILLER_232_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_408 ();
 DECAPx2_ASAP7_75t_R FILLER_232_423 ();
 FILLER_ASAP7_75t_R FILLER_232_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_431 ();
 DECAPx2_ASAP7_75t_R FILLER_232_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_446 ();
 DECAPx4_ASAP7_75t_R FILLER_232_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_463 ();
 DECAPx10_ASAP7_75t_R FILLER_232_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_492 ();
 DECAPx10_ASAP7_75t_R FILLER_232_501 ();
 DECAPx1_ASAP7_75t_R FILLER_232_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_527 ();
 DECAPx10_ASAP7_75t_R FILLER_232_538 ();
 DECAPx10_ASAP7_75t_R FILLER_232_560 ();
 DECAPx10_ASAP7_75t_R FILLER_232_582 ();
 DECAPx6_ASAP7_75t_R FILLER_232_604 ();
 DECAPx2_ASAP7_75t_R FILLER_232_618 ();
 DECAPx10_ASAP7_75t_R FILLER_232_634 ();
 DECAPx1_ASAP7_75t_R FILLER_232_656 ();
 DECAPx2_ASAP7_75t_R FILLER_232_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_672 ();
 DECAPx4_ASAP7_75t_R FILLER_232_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_705 ();
 DECAPx10_ASAP7_75t_R FILLER_232_717 ();
 DECAPx10_ASAP7_75t_R FILLER_232_739 ();
 DECAPx1_ASAP7_75t_R FILLER_232_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_765 ();
 DECAPx10_ASAP7_75t_R FILLER_232_772 ();
 DECAPx10_ASAP7_75t_R FILLER_232_794 ();
 DECAPx4_ASAP7_75t_R FILLER_232_816 ();
 FILLER_ASAP7_75t_R FILLER_232_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_828 ();
 DECAPx2_ASAP7_75t_R FILLER_232_843 ();
 FILLER_ASAP7_75t_R FILLER_232_849 ();
 DECAPx2_ASAP7_75t_R FILLER_232_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_886 ();
 DECAPx4_ASAP7_75t_R FILLER_232_890 ();
 DECAPx6_ASAP7_75t_R FILLER_232_908 ();
 DECAPx1_ASAP7_75t_R FILLER_232_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_926 ();
 DECAPx2_ASAP7_75t_R FILLER_232_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_936 ();
 DECAPx10_ASAP7_75t_R FILLER_232_945 ();
 DECAPx4_ASAP7_75t_R FILLER_232_967 ();
 FILLER_ASAP7_75t_R FILLER_232_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_979 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1026 ();
 FILLER_ASAP7_75t_R FILLER_232_1036 ();
 FILLER_ASAP7_75t_R FILLER_232_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1097 ();
 FILLER_ASAP7_75t_R FILLER_232_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1280 ();
 FILLER_ASAP7_75t_R FILLER_232_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_233_172 ();
 DECAPx10_ASAP7_75t_R FILLER_233_194 ();
 DECAPx10_ASAP7_75t_R FILLER_233_216 ();
 FILLER_ASAP7_75t_R FILLER_233_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_240 ();
 DECAPx1_ASAP7_75t_R FILLER_233_279 ();
 DECAPx2_ASAP7_75t_R FILLER_233_307 ();
 FILLER_ASAP7_75t_R FILLER_233_313 ();
 DECAPx1_ASAP7_75t_R FILLER_233_322 ();
 DECAPx4_ASAP7_75t_R FILLER_233_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_342 ();
 DECAPx2_ASAP7_75t_R FILLER_233_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_363 ();
 DECAPx10_ASAP7_75t_R FILLER_233_370 ();
 FILLER_ASAP7_75t_R FILLER_233_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_394 ();
 DECAPx10_ASAP7_75t_R FILLER_233_398 ();
 DECAPx2_ASAP7_75t_R FILLER_233_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_426 ();
 DECAPx10_ASAP7_75t_R FILLER_233_433 ();
 DECAPx10_ASAP7_75t_R FILLER_233_455 ();
 DECAPx2_ASAP7_75t_R FILLER_233_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_499 ();
 DECAPx10_ASAP7_75t_R FILLER_233_510 ();
 DECAPx10_ASAP7_75t_R FILLER_233_532 ();
 DECAPx10_ASAP7_75t_R FILLER_233_568 ();
 DECAPx10_ASAP7_75t_R FILLER_233_590 ();
 DECAPx10_ASAP7_75t_R FILLER_233_615 ();
 DECAPx10_ASAP7_75t_R FILLER_233_637 ();
 DECAPx6_ASAP7_75t_R FILLER_233_665 ();
 FILLER_ASAP7_75t_R FILLER_233_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_681 ();
 DECAPx1_ASAP7_75t_R FILLER_233_700 ();
 DECAPx10_ASAP7_75t_R FILLER_233_714 ();
 DECAPx4_ASAP7_75t_R FILLER_233_736 ();
 FILLER_ASAP7_75t_R FILLER_233_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_748 ();
 DECAPx1_ASAP7_75t_R FILLER_233_759 ();
 DECAPx4_ASAP7_75t_R FILLER_233_769 ();
 FILLER_ASAP7_75t_R FILLER_233_779 ();
 DECAPx10_ASAP7_75t_R FILLER_233_793 ();
 DECAPx2_ASAP7_75t_R FILLER_233_815 ();
 FILLER_ASAP7_75t_R FILLER_233_821 ();
 DECAPx10_ASAP7_75t_R FILLER_233_828 ();
 DECAPx6_ASAP7_75t_R FILLER_233_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_864 ();
 FILLER_ASAP7_75t_R FILLER_233_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_930 ();
 DECAPx10_ASAP7_75t_R FILLER_233_958 ();
 DECAPx10_ASAP7_75t_R FILLER_233_980 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1002 ();
 FILLER_ASAP7_75t_R FILLER_233_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1064 ();
 FILLER_ASAP7_75t_R FILLER_233_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1108 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_234_172 ();
 DECAPx10_ASAP7_75t_R FILLER_234_194 ();
 DECAPx10_ASAP7_75t_R FILLER_234_216 ();
 DECAPx10_ASAP7_75t_R FILLER_234_238 ();
 DECAPx6_ASAP7_75t_R FILLER_234_260 ();
 FILLER_ASAP7_75t_R FILLER_234_274 ();
 DECAPx6_ASAP7_75t_R FILLER_234_282 ();
 DECAPx10_ASAP7_75t_R FILLER_234_302 ();
 DECAPx10_ASAP7_75t_R FILLER_234_324 ();
 FILLER_ASAP7_75t_R FILLER_234_346 ();
 DECAPx2_ASAP7_75t_R FILLER_234_356 ();
 DECAPx2_ASAP7_75t_R FILLER_234_368 ();
 FILLER_ASAP7_75t_R FILLER_234_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_382 ();
 DECAPx2_ASAP7_75t_R FILLER_234_399 ();
 FILLER_ASAP7_75t_R FILLER_234_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_407 ();
 FILLER_ASAP7_75t_R FILLER_234_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_422 ();
 FILLER_ASAP7_75t_R FILLER_234_431 ();
 DECAPx6_ASAP7_75t_R FILLER_234_439 ();
 DECAPx1_ASAP7_75t_R FILLER_234_453 ();
 FILLER_ASAP7_75t_R FILLER_234_469 ();
 DECAPx1_ASAP7_75t_R FILLER_234_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_498 ();
 DECAPx6_ASAP7_75t_R FILLER_234_515 ();
 DECAPx2_ASAP7_75t_R FILLER_234_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_535 ();
 DECAPx4_ASAP7_75t_R FILLER_234_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_564 ();
 DECAPx2_ASAP7_75t_R FILLER_234_568 ();
 DECAPx2_ASAP7_75t_R FILLER_234_582 ();
 DECAPx6_ASAP7_75t_R FILLER_234_591 ();
 DECAPx2_ASAP7_75t_R FILLER_234_626 ();
 DECAPx1_ASAP7_75t_R FILLER_234_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_638 ();
 DECAPx6_ASAP7_75t_R FILLER_234_660 ();
 DECAPx2_ASAP7_75t_R FILLER_234_674 ();
 DECAPx4_ASAP7_75t_R FILLER_234_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_696 ();
 DECAPx10_ASAP7_75t_R FILLER_234_703 ();
 DECAPx4_ASAP7_75t_R FILLER_234_725 ();
 FILLER_ASAP7_75t_R FILLER_234_735 ();
 DECAPx4_ASAP7_75t_R FILLER_234_751 ();
 FILLER_ASAP7_75t_R FILLER_234_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_763 ();
 DECAPx6_ASAP7_75t_R FILLER_234_772 ();
 FILLER_ASAP7_75t_R FILLER_234_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_788 ();
 DECAPx4_ASAP7_75t_R FILLER_234_799 ();
 DECAPx4_ASAP7_75t_R FILLER_234_815 ();
 FILLER_ASAP7_75t_R FILLER_234_825 ();
 DECAPx2_ASAP7_75t_R FILLER_234_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_841 ();
 FILLER_ASAP7_75t_R FILLER_234_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_852 ();
 DECAPx6_ASAP7_75t_R FILLER_234_859 ();
 FILLER_ASAP7_75t_R FILLER_234_873 ();
 DECAPx10_ASAP7_75t_R FILLER_234_881 ();
 DECAPx4_ASAP7_75t_R FILLER_234_903 ();
 FILLER_ASAP7_75t_R FILLER_234_913 ();
 DECAPx10_ASAP7_75t_R FILLER_234_936 ();
 FILLER_ASAP7_75t_R FILLER_234_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_960 ();
 DECAPx1_ASAP7_75t_R FILLER_234_990 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1036 ();
 FILLER_ASAP7_75t_R FILLER_234_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1082 ();
 FILLER_ASAP7_75t_R FILLER_234_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1122 ();
 FILLER_ASAP7_75t_R FILLER_234_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_234_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_235_172 ();
 DECAPx10_ASAP7_75t_R FILLER_235_194 ();
 DECAPx4_ASAP7_75t_R FILLER_235_216 ();
 FILLER_ASAP7_75t_R FILLER_235_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_228 ();
 DECAPx10_ASAP7_75t_R FILLER_235_237 ();
 DECAPx10_ASAP7_75t_R FILLER_235_259 ();
 DECAPx10_ASAP7_75t_R FILLER_235_295 ();
 DECAPx10_ASAP7_75t_R FILLER_235_317 ();
 DECAPx6_ASAP7_75t_R FILLER_235_339 ();
 DECAPx2_ASAP7_75t_R FILLER_235_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_359 ();
 DECAPx1_ASAP7_75t_R FILLER_235_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_370 ();
 DECAPx2_ASAP7_75t_R FILLER_235_377 ();
 FILLER_ASAP7_75t_R FILLER_235_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_385 ();
 DECAPx10_ASAP7_75t_R FILLER_235_404 ();
 DECAPx4_ASAP7_75t_R FILLER_235_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_436 ();
 DECAPx6_ASAP7_75t_R FILLER_235_445 ();
 DECAPx4_ASAP7_75t_R FILLER_235_467 ();
 DECAPx2_ASAP7_75t_R FILLER_235_485 ();
 FILLER_ASAP7_75t_R FILLER_235_491 ();
 DECAPx6_ASAP7_75t_R FILLER_235_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_535 ();
 DECAPx1_ASAP7_75t_R FILLER_235_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_548 ();
 DECAPx4_ASAP7_75t_R FILLER_235_591 ();
 FILLER_ASAP7_75t_R FILLER_235_601 ();
 DECAPx10_ASAP7_75t_R FILLER_235_611 ();
 FILLER_ASAP7_75t_R FILLER_235_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_635 ();
 DECAPx10_ASAP7_75t_R FILLER_235_652 ();
 DECAPx10_ASAP7_75t_R FILLER_235_674 ();
 DECAPx10_ASAP7_75t_R FILLER_235_702 ();
 FILLER_ASAP7_75t_R FILLER_235_724 ();
 DECAPx10_ASAP7_75t_R FILLER_235_750 ();
 DECAPx10_ASAP7_75t_R FILLER_235_772 ();
 DECAPx6_ASAP7_75t_R FILLER_235_794 ();
 DECAPx2_ASAP7_75t_R FILLER_235_829 ();
 FILLER_ASAP7_75t_R FILLER_235_835 ();
 DECAPx2_ASAP7_75t_R FILLER_235_845 ();
 FILLER_ASAP7_75t_R FILLER_235_851 ();
 DECAPx2_ASAP7_75t_R FILLER_235_861 ();
 DECAPx4_ASAP7_75t_R FILLER_235_870 ();
 FILLER_ASAP7_75t_R FILLER_235_880 ();
 DECAPx10_ASAP7_75t_R FILLER_235_890 ();
 DECAPx6_ASAP7_75t_R FILLER_235_912 ();
 FILLER_ASAP7_75t_R FILLER_235_926 ();
 DECAPx1_ASAP7_75t_R FILLER_235_936 ();
 DECAPx10_ASAP7_75t_R FILLER_235_943 ();
 FILLER_ASAP7_75t_R FILLER_235_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_967 ();
 DECAPx6_ASAP7_75t_R FILLER_235_979 ();
 DECAPx2_ASAP7_75t_R FILLER_235_993 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1007 ();
 FILLER_ASAP7_75t_R FILLER_235_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1028 ();
 FILLER_ASAP7_75t_R FILLER_235_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1085 ();
 FILLER_ASAP7_75t_R FILLER_235_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1093 ();
 FILLER_ASAP7_75t_R FILLER_235_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1102 ();
 FILLER_ASAP7_75t_R FILLER_235_1108 ();
 FILLER_ASAP7_75t_R FILLER_235_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_235_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_236_172 ();
 DECAPx10_ASAP7_75t_R FILLER_236_194 ();
 DECAPx10_ASAP7_75t_R FILLER_236_216 ();
 DECAPx1_ASAP7_75t_R FILLER_236_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_242 ();
 DECAPx6_ASAP7_75t_R FILLER_236_257 ();
 FILLER_ASAP7_75t_R FILLER_236_271 ();
 DECAPx6_ASAP7_75t_R FILLER_236_280 ();
 DECAPx1_ASAP7_75t_R FILLER_236_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_298 ();
 DECAPx4_ASAP7_75t_R FILLER_236_305 ();
 FILLER_ASAP7_75t_R FILLER_236_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_317 ();
 DECAPx2_ASAP7_75t_R FILLER_236_324 ();
 FILLER_ASAP7_75t_R FILLER_236_330 ();
 FILLER_ASAP7_75t_R FILLER_236_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_340 ();
 DECAPx4_ASAP7_75t_R FILLER_236_355 ();
 FILLER_ASAP7_75t_R FILLER_236_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_367 ();
 DECAPx2_ASAP7_75t_R FILLER_236_383 ();
 DECAPx4_ASAP7_75t_R FILLER_236_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_405 ();
 DECAPx4_ASAP7_75t_R FILLER_236_412 ();
 DECAPx1_ASAP7_75t_R FILLER_236_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_434 ();
 FILLER_ASAP7_75t_R FILLER_236_443 ();
 DECAPx4_ASAP7_75t_R FILLER_236_451 ();
 DECAPx6_ASAP7_75t_R FILLER_236_469 ();
 FILLER_ASAP7_75t_R FILLER_236_483 ();
 DECAPx4_ASAP7_75t_R FILLER_236_495 ();
 FILLER_ASAP7_75t_R FILLER_236_505 ();
 DECAPx10_ASAP7_75t_R FILLER_236_513 ();
 DECAPx2_ASAP7_75t_R FILLER_236_535 ();
 FILLER_ASAP7_75t_R FILLER_236_541 ();
 DECAPx10_ASAP7_75t_R FILLER_236_553 ();
 DECAPx2_ASAP7_75t_R FILLER_236_575 ();
 FILLER_ASAP7_75t_R FILLER_236_595 ();
 DECAPx6_ASAP7_75t_R FILLER_236_611 ();
 DECAPx2_ASAP7_75t_R FILLER_236_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_631 ();
 DECAPx10_ASAP7_75t_R FILLER_236_634 ();
 DECAPx1_ASAP7_75t_R FILLER_236_656 ();
 FILLER_ASAP7_75t_R FILLER_236_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_668 ();
 FILLER_ASAP7_75t_R FILLER_236_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_679 ();
 DECAPx4_ASAP7_75t_R FILLER_236_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_693 ();
 DECAPx10_ASAP7_75t_R FILLER_236_710 ();
 DECAPx10_ASAP7_75t_R FILLER_236_732 ();
 DECAPx10_ASAP7_75t_R FILLER_236_754 ();
 DECAPx6_ASAP7_75t_R FILLER_236_776 ();
 DECAPx10_ASAP7_75t_R FILLER_236_797 ();
 DECAPx10_ASAP7_75t_R FILLER_236_819 ();
 FILLER_ASAP7_75t_R FILLER_236_841 ();
 FILLER_ASAP7_75t_R FILLER_236_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_881 ();
 DECAPx10_ASAP7_75t_R FILLER_236_891 ();
 DECAPx2_ASAP7_75t_R FILLER_236_913 ();
 DECAPx1_ASAP7_75t_R FILLER_236_927 ();
 FILLER_ASAP7_75t_R FILLER_236_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_954 ();
 DECAPx1_ASAP7_75t_R FILLER_236_966 ();
 DECAPx6_ASAP7_75t_R FILLER_236_976 ();
 DECAPx1_ASAP7_75t_R FILLER_236_990 ();
 DECAPx2_ASAP7_75t_R FILLER_236_1008 ();
 FILLER_ASAP7_75t_R FILLER_236_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1112 ();
 FILLER_ASAP7_75t_R FILLER_236_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_236_1151 ();
 FILLER_ASAP7_75t_R FILLER_236_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_236_1173 ();
 FILLER_ASAP7_75t_R FILLER_236_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_236_1281 ();
 FILLER_ASAP7_75t_R FILLER_236_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_237_172 ();
 DECAPx10_ASAP7_75t_R FILLER_237_194 ();
 DECAPx10_ASAP7_75t_R FILLER_237_216 ();
 DECAPx4_ASAP7_75t_R FILLER_237_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_248 ();
 FILLER_ASAP7_75t_R FILLER_237_252 ();
 DECAPx2_ASAP7_75t_R FILLER_237_267 ();
 FILLER_ASAP7_75t_R FILLER_237_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_275 ();
 DECAPx10_ASAP7_75t_R FILLER_237_282 ();
 DECAPx4_ASAP7_75t_R FILLER_237_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_321 ();
 FILLER_ASAP7_75t_R FILLER_237_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_332 ();
 DECAPx2_ASAP7_75t_R FILLER_237_339 ();
 FILLER_ASAP7_75t_R FILLER_237_345 ();
 DECAPx2_ASAP7_75t_R FILLER_237_353 ();
 DECAPx10_ASAP7_75t_R FILLER_237_377 ();
 DECAPx2_ASAP7_75t_R FILLER_237_399 ();
 FILLER_ASAP7_75t_R FILLER_237_405 ();
 FILLER_ASAP7_75t_R FILLER_237_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_421 ();
 FILLER_ASAP7_75t_R FILLER_237_442 ();
 DECAPx6_ASAP7_75t_R FILLER_237_450 ();
 FILLER_ASAP7_75t_R FILLER_237_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_474 ();
 DECAPx10_ASAP7_75t_R FILLER_237_497 ();
 DECAPx10_ASAP7_75t_R FILLER_237_519 ();
 DECAPx10_ASAP7_75t_R FILLER_237_541 ();
 DECAPx6_ASAP7_75t_R FILLER_237_563 ();
 DECAPx2_ASAP7_75t_R FILLER_237_577 ();
 DECAPx10_ASAP7_75t_R FILLER_237_618 ();
 DECAPx6_ASAP7_75t_R FILLER_237_640 ();
 FILLER_ASAP7_75t_R FILLER_237_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_656 ();
 DECAPx10_ASAP7_75t_R FILLER_237_686 ();
 DECAPx10_ASAP7_75t_R FILLER_237_708 ();
 DECAPx1_ASAP7_75t_R FILLER_237_730 ();
 DECAPx6_ASAP7_75t_R FILLER_237_744 ();
 DECAPx2_ASAP7_75t_R FILLER_237_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_764 ();
 DECAPx4_ASAP7_75t_R FILLER_237_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_785 ();
 DECAPx10_ASAP7_75t_R FILLER_237_793 ();
 DECAPx10_ASAP7_75t_R FILLER_237_815 ();
 DECAPx6_ASAP7_75t_R FILLER_237_837 ();
 DECAPx2_ASAP7_75t_R FILLER_237_857 ();
 FILLER_ASAP7_75t_R FILLER_237_863 ();
 FILLER_ASAP7_75t_R FILLER_237_886 ();
 DECAPx6_ASAP7_75t_R FILLER_237_899 ();
 DECAPx1_ASAP7_75t_R FILLER_237_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_924 ();
 DECAPx1_ASAP7_75t_R FILLER_237_928 ();
 DECAPx10_ASAP7_75t_R FILLER_237_974 ();
 DECAPx6_ASAP7_75t_R FILLER_237_996 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1051 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1073 ();
 FILLER_ASAP7_75t_R FILLER_237_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1085 ();
 FILLER_ASAP7_75t_R FILLER_237_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1129 ();
 FILLER_ASAP7_75t_R FILLER_237_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1169 ();
 FILLER_ASAP7_75t_R FILLER_237_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_238_172 ();
 DECAPx10_ASAP7_75t_R FILLER_238_194 ();
 DECAPx10_ASAP7_75t_R FILLER_238_216 ();
 DECAPx4_ASAP7_75t_R FILLER_238_238 ();
 FILLER_ASAP7_75t_R FILLER_238_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_250 ();
 DECAPx2_ASAP7_75t_R FILLER_238_269 ();
 DECAPx2_ASAP7_75t_R FILLER_238_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_314 ();
 DECAPx10_ASAP7_75t_R FILLER_238_325 ();
 DECAPx6_ASAP7_75t_R FILLER_238_347 ();
 DECAPx10_ASAP7_75t_R FILLER_238_368 ();
 DECAPx6_ASAP7_75t_R FILLER_238_390 ();
 FILLER_ASAP7_75t_R FILLER_238_404 ();
 DECAPx10_ASAP7_75t_R FILLER_238_417 ();
 DECAPx10_ASAP7_75t_R FILLER_238_439 ();
 DECAPx2_ASAP7_75t_R FILLER_238_461 ();
 FILLER_ASAP7_75t_R FILLER_238_467 ();
 DECAPx10_ASAP7_75t_R FILLER_238_481 ();
 DECAPx10_ASAP7_75t_R FILLER_238_503 ();
 DECAPx10_ASAP7_75t_R FILLER_238_525 ();
 DECAPx10_ASAP7_75t_R FILLER_238_547 ();
 DECAPx10_ASAP7_75t_R FILLER_238_569 ();
 DECAPx2_ASAP7_75t_R FILLER_238_591 ();
 FILLER_ASAP7_75t_R FILLER_238_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_599 ();
 DECAPx4_ASAP7_75t_R FILLER_238_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_631 ();
 DECAPx10_ASAP7_75t_R FILLER_238_634 ();
 DECAPx10_ASAP7_75t_R FILLER_238_656 ();
 DECAPx10_ASAP7_75t_R FILLER_238_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_700 ();
 FILLER_ASAP7_75t_R FILLER_238_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_711 ();
 DECAPx2_ASAP7_75t_R FILLER_238_715 ();
 DECAPx2_ASAP7_75t_R FILLER_238_729 ();
 FILLER_ASAP7_75t_R FILLER_238_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_737 ();
 DECAPx6_ASAP7_75t_R FILLER_238_756 ();
 FILLER_ASAP7_75t_R FILLER_238_770 ();
 DECAPx10_ASAP7_75t_R FILLER_238_788 ();
 DECAPx1_ASAP7_75t_R FILLER_238_810 ();
 DECAPx10_ASAP7_75t_R FILLER_238_834 ();
 DECAPx10_ASAP7_75t_R FILLER_238_856 ();
 DECAPx1_ASAP7_75t_R FILLER_238_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_882 ();
 DECAPx2_ASAP7_75t_R FILLER_238_904 ();
 DECAPx10_ASAP7_75t_R FILLER_238_931 ();
 DECAPx6_ASAP7_75t_R FILLER_238_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_974 ();
 FILLER_ASAP7_75t_R FILLER_238_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_980 ();
 DECAPx2_ASAP7_75t_R FILLER_238_998 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1127 ();
 FILLER_ASAP7_75t_R FILLER_238_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_239_172 ();
 DECAPx10_ASAP7_75t_R FILLER_239_194 ();
 DECAPx10_ASAP7_75t_R FILLER_239_216 ();
 DECAPx4_ASAP7_75t_R FILLER_239_238 ();
 FILLER_ASAP7_75t_R FILLER_239_248 ();
 DECAPx10_ASAP7_75t_R FILLER_239_256 ();
 DECAPx4_ASAP7_75t_R FILLER_239_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_294 ();
 DECAPx10_ASAP7_75t_R FILLER_239_306 ();
 FILLER_ASAP7_75t_R FILLER_239_328 ();
 DECAPx6_ASAP7_75t_R FILLER_239_345 ();
 DECAPx1_ASAP7_75t_R FILLER_239_359 ();
 DECAPx6_ASAP7_75t_R FILLER_239_369 ();
 DECAPx1_ASAP7_75t_R FILLER_239_383 ();
 DECAPx10_ASAP7_75t_R FILLER_239_395 ();
 DECAPx6_ASAP7_75t_R FILLER_239_417 ();
 FILLER_ASAP7_75t_R FILLER_239_431 ();
 DECAPx1_ASAP7_75t_R FILLER_239_439 ();
 DECAPx6_ASAP7_75t_R FILLER_239_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_467 ();
 DECAPx2_ASAP7_75t_R FILLER_239_476 ();
 DECAPx10_ASAP7_75t_R FILLER_239_490 ();
 DECAPx10_ASAP7_75t_R FILLER_239_512 ();
 DECAPx10_ASAP7_75t_R FILLER_239_534 ();
 DECAPx10_ASAP7_75t_R FILLER_239_556 ();
 DECAPx2_ASAP7_75t_R FILLER_239_578 ();
 FILLER_ASAP7_75t_R FILLER_239_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_609 ();
 DECAPx6_ASAP7_75t_R FILLER_239_616 ();
 FILLER_ASAP7_75t_R FILLER_239_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_632 ();
 DECAPx10_ASAP7_75t_R FILLER_239_639 ();
 DECAPx6_ASAP7_75t_R FILLER_239_661 ();
 DECAPx1_ASAP7_75t_R FILLER_239_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_679 ();
 DECAPx2_ASAP7_75t_R FILLER_239_686 ();
 FILLER_ASAP7_75t_R FILLER_239_692 ();
 DECAPx10_ASAP7_75t_R FILLER_239_715 ();
 DECAPx2_ASAP7_75t_R FILLER_239_737 ();
 FILLER_ASAP7_75t_R FILLER_239_743 ();
 DECAPx10_ASAP7_75t_R FILLER_239_757 ();
 DECAPx2_ASAP7_75t_R FILLER_239_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_785 ();
 DECAPx10_ASAP7_75t_R FILLER_239_792 ();
 DECAPx10_ASAP7_75t_R FILLER_239_814 ();
 DECAPx4_ASAP7_75t_R FILLER_239_836 ();
 FILLER_ASAP7_75t_R FILLER_239_846 ();
 DECAPx2_ASAP7_75t_R FILLER_239_854 ();
 DECAPx4_ASAP7_75t_R FILLER_239_866 ();
 FILLER_ASAP7_75t_R FILLER_239_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_878 ();
 DECAPx4_ASAP7_75t_R FILLER_239_887 ();
 FILLER_ASAP7_75t_R FILLER_239_897 ();
 DECAPx10_ASAP7_75t_R FILLER_239_905 ();
 DECAPx10_ASAP7_75t_R FILLER_239_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_978 ();
 FILLER_ASAP7_75t_R FILLER_239_1000 ();
 FILLER_ASAP7_75t_R FILLER_239_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_239_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_240_172 ();
 DECAPx10_ASAP7_75t_R FILLER_240_194 ();
 DECAPx10_ASAP7_75t_R FILLER_240_216 ();
 DECAPx1_ASAP7_75t_R FILLER_240_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_242 ();
 DECAPx4_ASAP7_75t_R FILLER_240_246 ();
 DECAPx6_ASAP7_75t_R FILLER_240_266 ();
 DECAPx2_ASAP7_75t_R FILLER_240_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_286 ();
 DECAPx6_ASAP7_75t_R FILLER_240_302 ();
 DECAPx2_ASAP7_75t_R FILLER_240_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_322 ();
 DECAPx2_ASAP7_75t_R FILLER_240_329 ();
 DECAPx2_ASAP7_75t_R FILLER_240_346 ();
 FILLER_ASAP7_75t_R FILLER_240_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_354 ();
 DECAPx4_ASAP7_75t_R FILLER_240_361 ();
 FILLER_ASAP7_75t_R FILLER_240_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_404 ();
 DECAPx1_ASAP7_75t_R FILLER_240_417 ();
 DECAPx1_ASAP7_75t_R FILLER_240_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_431 ();
 DECAPx2_ASAP7_75t_R FILLER_240_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_444 ();
 DECAPx2_ASAP7_75t_R FILLER_240_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_472 ();
 DECAPx6_ASAP7_75t_R FILLER_240_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_495 ();
 DECAPx10_ASAP7_75t_R FILLER_240_502 ();
 DECAPx10_ASAP7_75t_R FILLER_240_524 ();
 DECAPx10_ASAP7_75t_R FILLER_240_546 ();
 DECAPx10_ASAP7_75t_R FILLER_240_568 ();
 DECAPx2_ASAP7_75t_R FILLER_240_590 ();
 FILLER_ASAP7_75t_R FILLER_240_596 ();
 DECAPx2_ASAP7_75t_R FILLER_240_606 ();
 FILLER_ASAP7_75t_R FILLER_240_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_631 ();
 FILLER_ASAP7_75t_R FILLER_240_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_636 ();
 DECAPx6_ASAP7_75t_R FILLER_240_648 ();
 DECAPx2_ASAP7_75t_R FILLER_240_662 ();
 DECAPx2_ASAP7_75t_R FILLER_240_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_682 ();
 DECAPx2_ASAP7_75t_R FILLER_240_689 ();
 FILLER_ASAP7_75t_R FILLER_240_695 ();
 DECAPx10_ASAP7_75t_R FILLER_240_705 ();
 DECAPx10_ASAP7_75t_R FILLER_240_727 ();
 DECAPx10_ASAP7_75t_R FILLER_240_749 ();
 DECAPx10_ASAP7_75t_R FILLER_240_771 ();
 DECAPx6_ASAP7_75t_R FILLER_240_793 ();
 DECAPx2_ASAP7_75t_R FILLER_240_807 ();
 DECAPx10_ASAP7_75t_R FILLER_240_820 ();
 DECAPx2_ASAP7_75t_R FILLER_240_842 ();
 FILLER_ASAP7_75t_R FILLER_240_848 ();
 DECAPx6_ASAP7_75t_R FILLER_240_856 ();
 DECAPx1_ASAP7_75t_R FILLER_240_870 ();
 DECAPx2_ASAP7_75t_R FILLER_240_912 ();
 FILLER_ASAP7_75t_R FILLER_240_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_920 ();
 DECAPx2_ASAP7_75t_R FILLER_240_942 ();
 FILLER_ASAP7_75t_R FILLER_240_948 ();
 DECAPx10_ASAP7_75t_R FILLER_240_971 ();
 DECAPx10_ASAP7_75t_R FILLER_240_993 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_240_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_240_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1281 ();
 FILLER_ASAP7_75t_R FILLER_240_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_241_172 ();
 DECAPx10_ASAP7_75t_R FILLER_241_194 ();
 DECAPx10_ASAP7_75t_R FILLER_241_216 ();
 DECAPx10_ASAP7_75t_R FILLER_241_238 ();
 DECAPx2_ASAP7_75t_R FILLER_241_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_266 ();
 DECAPx1_ASAP7_75t_R FILLER_241_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_277 ();
 DECAPx4_ASAP7_75t_R FILLER_241_292 ();
 DECAPx4_ASAP7_75t_R FILLER_241_310 ();
 FILLER_ASAP7_75t_R FILLER_241_320 ();
 DECAPx2_ASAP7_75t_R FILLER_241_344 ();
 FILLER_ASAP7_75t_R FILLER_241_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_352 ();
 DECAPx2_ASAP7_75t_R FILLER_241_361 ();
 FILLER_ASAP7_75t_R FILLER_241_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_369 ();
 DECAPx4_ASAP7_75t_R FILLER_241_378 ();
 FILLER_ASAP7_75t_R FILLER_241_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_398 ();
 DECAPx2_ASAP7_75t_R FILLER_241_405 ();
 DECAPx4_ASAP7_75t_R FILLER_241_433 ();
 FILLER_ASAP7_75t_R FILLER_241_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_445 ();
 DECAPx4_ASAP7_75t_R FILLER_241_456 ();
 FILLER_ASAP7_75t_R FILLER_241_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_468 ();
 DECAPx1_ASAP7_75t_R FILLER_241_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_481 ();
 DECAPx1_ASAP7_75t_R FILLER_241_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_492 ();
 FILLER_ASAP7_75t_R FILLER_241_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_501 ();
 DECAPx10_ASAP7_75t_R FILLER_241_510 ();
 DECAPx10_ASAP7_75t_R FILLER_241_532 ();
 DECAPx10_ASAP7_75t_R FILLER_241_554 ();
 DECAPx10_ASAP7_75t_R FILLER_241_576 ();
 DECAPx4_ASAP7_75t_R FILLER_241_598 ();
 FILLER_ASAP7_75t_R FILLER_241_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_631 ();
 DECAPx4_ASAP7_75t_R FILLER_241_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_663 ();
 DECAPx10_ASAP7_75t_R FILLER_241_667 ();
 DECAPx10_ASAP7_75t_R FILLER_241_689 ();
 DECAPx10_ASAP7_75t_R FILLER_241_711 ();
 DECAPx10_ASAP7_75t_R FILLER_241_733 ();
 DECAPx10_ASAP7_75t_R FILLER_241_755 ();
 DECAPx6_ASAP7_75t_R FILLER_241_777 ();
 DECAPx2_ASAP7_75t_R FILLER_241_791 ();
 DECAPx10_ASAP7_75t_R FILLER_241_801 ();
 DECAPx10_ASAP7_75t_R FILLER_241_823 ();
 DECAPx10_ASAP7_75t_R FILLER_241_845 ();
 DECAPx10_ASAP7_75t_R FILLER_241_867 ();
 DECAPx6_ASAP7_75t_R FILLER_241_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_903 ();
 DECAPx2_ASAP7_75t_R FILLER_241_918 ();
 FILLER_ASAP7_75t_R FILLER_241_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_935 ();
 DECAPx4_ASAP7_75t_R FILLER_241_939 ();
 FILLER_ASAP7_75t_R FILLER_241_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_965 ();
 DECAPx10_ASAP7_75t_R FILLER_241_969 ();
 DECAPx6_ASAP7_75t_R FILLER_241_991 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_241_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1120 ();
 FILLER_ASAP7_75t_R FILLER_241_1134 ();
 FILLER_ASAP7_75t_R FILLER_241_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1269 ();
 FILLER_ASAP7_75t_R FILLER_241_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_242_172 ();
 DECAPx10_ASAP7_75t_R FILLER_242_194 ();
 DECAPx10_ASAP7_75t_R FILLER_242_216 ();
 DECAPx10_ASAP7_75t_R FILLER_242_238 ();
 DECAPx1_ASAP7_75t_R FILLER_242_260 ();
 DECAPx4_ASAP7_75t_R FILLER_242_278 ();
 FILLER_ASAP7_75t_R FILLER_242_288 ();
 FILLER_ASAP7_75t_R FILLER_242_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_300 ();
 DECAPx2_ASAP7_75t_R FILLER_242_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_315 ();
 DECAPx10_ASAP7_75t_R FILLER_242_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_352 ();
 DECAPx2_ASAP7_75t_R FILLER_242_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_383 ();
 DECAPx2_ASAP7_75t_R FILLER_242_390 ();
 FILLER_ASAP7_75t_R FILLER_242_396 ();
 DECAPx1_ASAP7_75t_R FILLER_242_406 ();
 DECAPx10_ASAP7_75t_R FILLER_242_416 ();
 DECAPx2_ASAP7_75t_R FILLER_242_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_444 ();
 DECAPx6_ASAP7_75t_R FILLER_242_452 ();
 DECAPx2_ASAP7_75t_R FILLER_242_466 ();
 DECAPx1_ASAP7_75t_R FILLER_242_485 ();
 DECAPx1_ASAP7_75t_R FILLER_242_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_499 ();
 DECAPx10_ASAP7_75t_R FILLER_242_516 ();
 DECAPx10_ASAP7_75t_R FILLER_242_538 ();
 DECAPx6_ASAP7_75t_R FILLER_242_560 ();
 FILLER_ASAP7_75t_R FILLER_242_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_576 ();
 DECAPx10_ASAP7_75t_R FILLER_242_587 ();
 DECAPx6_ASAP7_75t_R FILLER_242_609 ();
 DECAPx6_ASAP7_75t_R FILLER_242_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_648 ();
 DECAPx10_ASAP7_75t_R FILLER_242_670 ();
 DECAPx1_ASAP7_75t_R FILLER_242_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_696 ();
 DECAPx2_ASAP7_75t_R FILLER_242_705 ();
 FILLER_ASAP7_75t_R FILLER_242_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_737 ();
 DECAPx2_ASAP7_75t_R FILLER_242_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_755 ();
 DECAPx6_ASAP7_75t_R FILLER_242_777 ();
 DECAPx4_ASAP7_75t_R FILLER_242_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_817 ();
 FILLER_ASAP7_75t_R FILLER_242_832 ();
 DECAPx2_ASAP7_75t_R FILLER_242_837 ();
 FILLER_ASAP7_75t_R FILLER_242_843 ();
 DECAPx10_ASAP7_75t_R FILLER_242_851 ();
 FILLER_ASAP7_75t_R FILLER_242_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_875 ();
 DECAPx4_ASAP7_75t_R FILLER_242_884 ();
 DECAPx10_ASAP7_75t_R FILLER_242_945 ();
 DECAPx10_ASAP7_75t_R FILLER_242_967 ();
 DECAPx6_ASAP7_75t_R FILLER_242_989 ();
 FILLER_ASAP7_75t_R FILLER_242_1003 ();
 FILLER_ASAP7_75t_R FILLER_242_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_242_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_242_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_242_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_243_172 ();
 DECAPx10_ASAP7_75t_R FILLER_243_194 ();
 DECAPx10_ASAP7_75t_R FILLER_243_216 ();
 DECAPx10_ASAP7_75t_R FILLER_243_238 ();
 DECAPx4_ASAP7_75t_R FILLER_243_260 ();
 FILLER_ASAP7_75t_R FILLER_243_270 ();
 DECAPx1_ASAP7_75t_R FILLER_243_278 ();
 DECAPx10_ASAP7_75t_R FILLER_243_304 ();
 DECAPx6_ASAP7_75t_R FILLER_243_326 ();
 FILLER_ASAP7_75t_R FILLER_243_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_342 ();
 DECAPx6_ASAP7_75t_R FILLER_243_363 ();
 FILLER_ASAP7_75t_R FILLER_243_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_379 ();
 DECAPx6_ASAP7_75t_R FILLER_243_395 ();
 DECAPx1_ASAP7_75t_R FILLER_243_409 ();
 DECAPx10_ASAP7_75t_R FILLER_243_419 ();
 DECAPx1_ASAP7_75t_R FILLER_243_441 ();
 FILLER_ASAP7_75t_R FILLER_243_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_483 ();
 DECAPx1_ASAP7_75t_R FILLER_243_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_494 ();
 DECAPx10_ASAP7_75t_R FILLER_243_501 ();
 DECAPx10_ASAP7_75t_R FILLER_243_523 ();
 DECAPx10_ASAP7_75t_R FILLER_243_545 ();
 DECAPx10_ASAP7_75t_R FILLER_243_567 ();
 DECAPx6_ASAP7_75t_R FILLER_243_589 ();
 DECAPx1_ASAP7_75t_R FILLER_243_603 ();
 DECAPx10_ASAP7_75t_R FILLER_243_615 ();
 DECAPx6_ASAP7_75t_R FILLER_243_637 ();
 FILLER_ASAP7_75t_R FILLER_243_651 ();
 DECAPx2_ASAP7_75t_R FILLER_243_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_673 ();
 DECAPx1_ASAP7_75t_R FILLER_243_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_694 ();
 DECAPx2_ASAP7_75t_R FILLER_243_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_715 ();
 DECAPx2_ASAP7_75t_R FILLER_243_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_730 ();
 DECAPx2_ASAP7_75t_R FILLER_243_772 ();
 FILLER_ASAP7_75t_R FILLER_243_778 ();
 FILLER_ASAP7_75t_R FILLER_243_783 ();
 DECAPx2_ASAP7_75t_R FILLER_243_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_849 ();
 DECAPx6_ASAP7_75t_R FILLER_243_858 ();
 FILLER_ASAP7_75t_R FILLER_243_872 ();
 DECAPx10_ASAP7_75t_R FILLER_243_882 ();
 DECAPx6_ASAP7_75t_R FILLER_243_904 ();
 DECAPx2_ASAP7_75t_R FILLER_243_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_924 ();
 DECAPx1_ASAP7_75t_R FILLER_243_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_941 ();
 DECAPx10_ASAP7_75t_R FILLER_243_951 ();
 DECAPx1_ASAP7_75t_R FILLER_243_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_977 ();
 DECAPx2_ASAP7_75t_R FILLER_243_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_992 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_243_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_243_1086 ();
 FILLER_ASAP7_75t_R FILLER_243_1092 ();
 DECAPx4_ASAP7_75t_R FILLER_243_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_243_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_243_1148 ();
 FILLER_ASAP7_75t_R FILLER_243_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_243_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_244_172 ();
 DECAPx10_ASAP7_75t_R FILLER_244_194 ();
 DECAPx10_ASAP7_75t_R FILLER_244_216 ();
 DECAPx10_ASAP7_75t_R FILLER_244_238 ();
 DECAPx6_ASAP7_75t_R FILLER_244_260 ();
 DECAPx2_ASAP7_75t_R FILLER_244_274 ();
 DECAPx10_ASAP7_75t_R FILLER_244_298 ();
 DECAPx10_ASAP7_75t_R FILLER_244_320 ();
 DECAPx2_ASAP7_75t_R FILLER_244_342 ();
 FILLER_ASAP7_75t_R FILLER_244_348 ();
 DECAPx2_ASAP7_75t_R FILLER_244_358 ();
 FILLER_ASAP7_75t_R FILLER_244_364 ();
 DECAPx2_ASAP7_75t_R FILLER_244_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_382 ();
 DECAPx6_ASAP7_75t_R FILLER_244_390 ();
 DECAPx2_ASAP7_75t_R FILLER_244_404 ();
 DECAPx2_ASAP7_75t_R FILLER_244_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_428 ();
 FILLER_ASAP7_75t_R FILLER_244_442 ();
 DECAPx2_ASAP7_75t_R FILLER_244_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_468 ();
 FILLER_ASAP7_75t_R FILLER_244_476 ();
 DECAPx10_ASAP7_75t_R FILLER_244_496 ();
 DECAPx10_ASAP7_75t_R FILLER_244_518 ();
 DECAPx4_ASAP7_75t_R FILLER_244_540 ();
 DECAPx10_ASAP7_75t_R FILLER_244_568 ();
 DECAPx10_ASAP7_75t_R FILLER_244_590 ();
 DECAPx2_ASAP7_75t_R FILLER_244_612 ();
 FILLER_ASAP7_75t_R FILLER_244_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_631 ();
 DECAPx10_ASAP7_75t_R FILLER_244_634 ();
 DECAPx2_ASAP7_75t_R FILLER_244_656 ();
 FILLER_ASAP7_75t_R FILLER_244_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_664 ();
 DECAPx6_ASAP7_75t_R FILLER_244_673 ();
 FILLER_ASAP7_75t_R FILLER_244_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_689 ();
 DECAPx4_ASAP7_75t_R FILLER_244_704 ();
 FILLER_ASAP7_75t_R FILLER_244_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_716 ();
 DECAPx2_ASAP7_75t_R FILLER_244_725 ();
 FILLER_ASAP7_75t_R FILLER_244_731 ();
 DECAPx10_ASAP7_75t_R FILLER_244_757 ();
 DECAPx4_ASAP7_75t_R FILLER_244_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_789 ();
 DECAPx4_ASAP7_75t_R FILLER_244_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_806 ();
 DECAPx10_ASAP7_75t_R FILLER_244_818 ();
 DECAPx4_ASAP7_75t_R FILLER_244_840 ();
 FILLER_ASAP7_75t_R FILLER_244_856 ();
 DECAPx10_ASAP7_75t_R FILLER_244_882 ();
 DECAPx6_ASAP7_75t_R FILLER_244_904 ();
 DECAPx1_ASAP7_75t_R FILLER_244_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_922 ();
 DECAPx4_ASAP7_75t_R FILLER_244_934 ();
 DECAPx2_ASAP7_75t_R FILLER_244_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_958 ();
 DECAPx1_ASAP7_75t_R FILLER_244_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_971 ();
 DECAPx4_ASAP7_75t_R FILLER_244_993 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1098 ();
 FILLER_ASAP7_75t_R FILLER_244_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1125 ();
 FILLER_ASAP7_75t_R FILLER_244_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_245_172 ();
 DECAPx10_ASAP7_75t_R FILLER_245_194 ();
 DECAPx10_ASAP7_75t_R FILLER_245_216 ();
 DECAPx10_ASAP7_75t_R FILLER_245_238 ();
 DECAPx10_ASAP7_75t_R FILLER_245_260 ();
 FILLER_ASAP7_75t_R FILLER_245_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_284 ();
 DECAPx2_ASAP7_75t_R FILLER_245_305 ();
 FILLER_ASAP7_75t_R FILLER_245_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_327 ();
 DECAPx1_ASAP7_75t_R FILLER_245_342 ();
 FILLER_ASAP7_75t_R FILLER_245_354 ();
 DECAPx2_ASAP7_75t_R FILLER_245_364 ();
 FILLER_ASAP7_75t_R FILLER_245_370 ();
 FILLER_ASAP7_75t_R FILLER_245_382 ();
 DECAPx6_ASAP7_75t_R FILLER_245_390 ();
 DECAPx1_ASAP7_75t_R FILLER_245_404 ();
 DECAPx1_ASAP7_75t_R FILLER_245_420 ();
 FILLER_ASAP7_75t_R FILLER_245_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_441 ();
 DECAPx10_ASAP7_75t_R FILLER_245_464 ();
 DECAPx2_ASAP7_75t_R FILLER_245_486 ();
 DECAPx10_ASAP7_75t_R FILLER_245_512 ();
 DECAPx10_ASAP7_75t_R FILLER_245_534 ();
 DECAPx10_ASAP7_75t_R FILLER_245_556 ();
 DECAPx10_ASAP7_75t_R FILLER_245_578 ();
 DECAPx2_ASAP7_75t_R FILLER_245_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_606 ();
 DECAPx1_ASAP7_75t_R FILLER_245_628 ();
 DECAPx10_ASAP7_75t_R FILLER_245_656 ();
 DECAPx4_ASAP7_75t_R FILLER_245_678 ();
 FILLER_ASAP7_75t_R FILLER_245_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_690 ();
 DECAPx2_ASAP7_75t_R FILLER_245_699 ();
 FILLER_ASAP7_75t_R FILLER_245_705 ();
 DECAPx10_ASAP7_75t_R FILLER_245_710 ();
 DECAPx10_ASAP7_75t_R FILLER_245_732 ();
 DECAPx10_ASAP7_75t_R FILLER_245_762 ();
 FILLER_ASAP7_75t_R FILLER_245_784 ();
 DECAPx2_ASAP7_75t_R FILLER_245_792 ();
 FILLER_ASAP7_75t_R FILLER_245_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_822 ();
 DECAPx10_ASAP7_75t_R FILLER_245_831 ();
 FILLER_ASAP7_75t_R FILLER_245_853 ();
 DECAPx6_ASAP7_75t_R FILLER_245_886 ();
 FILLER_ASAP7_75t_R FILLER_245_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_962 ();
 DECAPx4_ASAP7_75t_R FILLER_245_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_976 ();
 DECAPx2_ASAP7_75t_R FILLER_245_986 ();
 FILLER_ASAP7_75t_R FILLER_245_992 ();
 DECAPx2_ASAP7_75t_R FILLER_245_997 ();
 FILLER_ASAP7_75t_R FILLER_245_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1033 ();
 FILLER_ASAP7_75t_R FILLER_245_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1057 ();
 FILLER_ASAP7_75t_R FILLER_245_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1083 ();
 FILLER_ASAP7_75t_R FILLER_245_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1096 ();
 FILLER_ASAP7_75t_R FILLER_245_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1120 ();
 FILLER_ASAP7_75t_R FILLER_245_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_246_172 ();
 DECAPx10_ASAP7_75t_R FILLER_246_194 ();
 DECAPx10_ASAP7_75t_R FILLER_246_216 ();
 DECAPx10_ASAP7_75t_R FILLER_246_238 ();
 DECAPx10_ASAP7_75t_R FILLER_246_260 ();
 DECAPx2_ASAP7_75t_R FILLER_246_282 ();
 FILLER_ASAP7_75t_R FILLER_246_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_290 ();
 FILLER_ASAP7_75t_R FILLER_246_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_321 ();
 FILLER_ASAP7_75t_R FILLER_246_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_330 ();
 DECAPx1_ASAP7_75t_R FILLER_246_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_347 ();
 DECAPx6_ASAP7_75t_R FILLER_246_366 ();
 DECAPx2_ASAP7_75t_R FILLER_246_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_386 ();
 FILLER_ASAP7_75t_R FILLER_246_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_395 ();
 DECAPx2_ASAP7_75t_R FILLER_246_410 ();
 DECAPx10_ASAP7_75t_R FILLER_246_424 ();
 DECAPx6_ASAP7_75t_R FILLER_246_446 ();
 DECAPx2_ASAP7_75t_R FILLER_246_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_466 ();
 DECAPx2_ASAP7_75t_R FILLER_246_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_481 ();
 DECAPx10_ASAP7_75t_R FILLER_246_490 ();
 DECAPx10_ASAP7_75t_R FILLER_246_512 ();
 DECAPx10_ASAP7_75t_R FILLER_246_534 ();
 DECAPx10_ASAP7_75t_R FILLER_246_556 ();
 DECAPx10_ASAP7_75t_R FILLER_246_578 ();
 DECAPx6_ASAP7_75t_R FILLER_246_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_614 ();
 FILLER_ASAP7_75t_R FILLER_246_622 ();
 FILLER_ASAP7_75t_R FILLER_246_634 ();
 FILLER_ASAP7_75t_R FILLER_246_652 ();
 DECAPx10_ASAP7_75t_R FILLER_246_678 ();
 FILLER_ASAP7_75t_R FILLER_246_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_702 ();
 DECAPx6_ASAP7_75t_R FILLER_246_711 ();
 FILLER_ASAP7_75t_R FILLER_246_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_727 ();
 DECAPx1_ASAP7_75t_R FILLER_246_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_770 ();
 DECAPx10_ASAP7_75t_R FILLER_246_779 ();
 DECAPx2_ASAP7_75t_R FILLER_246_801 ();
 FILLER_ASAP7_75t_R FILLER_246_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_809 ();
 DECAPx10_ASAP7_75t_R FILLER_246_824 ();
 DECAPx2_ASAP7_75t_R FILLER_246_846 ();
 DECAPx1_ASAP7_75t_R FILLER_246_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_863 ();
 DECAPx6_ASAP7_75t_R FILLER_246_880 ();
 DECAPx1_ASAP7_75t_R FILLER_246_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_898 ();
 FILLER_ASAP7_75t_R FILLER_246_907 ();
 DECAPx10_ASAP7_75t_R FILLER_246_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_934 ();
 DECAPx1_ASAP7_75t_R FILLER_246_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_943 ();
 DECAPx4_ASAP7_75t_R FILLER_246_965 ();
 FILLER_ASAP7_75t_R FILLER_246_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_246_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1269 ();
 FILLER_ASAP7_75t_R FILLER_246_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_247_172 ();
 DECAPx10_ASAP7_75t_R FILLER_247_194 ();
 DECAPx10_ASAP7_75t_R FILLER_247_216 ();
 DECAPx10_ASAP7_75t_R FILLER_247_238 ();
 DECAPx6_ASAP7_75t_R FILLER_247_260 ();
 DECAPx1_ASAP7_75t_R FILLER_247_274 ();
 DECAPx1_ASAP7_75t_R FILLER_247_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_288 ();
 DECAPx10_ASAP7_75t_R FILLER_247_299 ();
 DECAPx10_ASAP7_75t_R FILLER_247_321 ();
 DECAPx6_ASAP7_75t_R FILLER_247_343 ();
 DECAPx1_ASAP7_75t_R FILLER_247_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_361 ();
 DECAPx6_ASAP7_75t_R FILLER_247_374 ();
 DECAPx10_ASAP7_75t_R FILLER_247_400 ();
 DECAPx10_ASAP7_75t_R FILLER_247_422 ();
 DECAPx2_ASAP7_75t_R FILLER_247_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_450 ();
 DECAPx2_ASAP7_75t_R FILLER_247_459 ();
 FILLER_ASAP7_75t_R FILLER_247_465 ();
 DECAPx2_ASAP7_75t_R FILLER_247_491 ();
 DECAPx10_ASAP7_75t_R FILLER_247_511 ();
 DECAPx10_ASAP7_75t_R FILLER_247_533 ();
 DECAPx10_ASAP7_75t_R FILLER_247_555 ();
 DECAPx10_ASAP7_75t_R FILLER_247_577 ();
 DECAPx6_ASAP7_75t_R FILLER_247_599 ();
 DECAPx4_ASAP7_75t_R FILLER_247_636 ();
 DECAPx10_ASAP7_75t_R FILLER_247_666 ();
 DECAPx6_ASAP7_75t_R FILLER_247_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_731 ();
 DECAPx4_ASAP7_75t_R FILLER_247_741 ();
 DECAPx10_ASAP7_75t_R FILLER_247_757 ();
 DECAPx1_ASAP7_75t_R FILLER_247_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_783 ();
 FILLER_ASAP7_75t_R FILLER_247_792 ();
 DECAPx2_ASAP7_75t_R FILLER_247_797 ();
 DECAPx4_ASAP7_75t_R FILLER_247_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_825 ();
 DECAPx4_ASAP7_75t_R FILLER_247_834 ();
 FILLER_ASAP7_75t_R FILLER_247_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_846 ();
 DECAPx10_ASAP7_75t_R FILLER_247_855 ();
 DECAPx4_ASAP7_75t_R FILLER_247_877 ();
 FILLER_ASAP7_75t_R FILLER_247_887 ();
 DECAPx1_ASAP7_75t_R FILLER_247_910 ();
 DECAPx10_ASAP7_75t_R FILLER_247_935 ();
 DECAPx6_ASAP7_75t_R FILLER_247_957 ();
 DECAPx1_ASAP7_75t_R FILLER_247_971 ();
 DECAPx10_ASAP7_75t_R FILLER_247_979 ();
 DECAPx4_ASAP7_75t_R FILLER_247_1001 ();
 FILLER_ASAP7_75t_R FILLER_247_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_247_1050 ();
 FILLER_ASAP7_75t_R FILLER_247_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1066 ();
 FILLER_ASAP7_75t_R FILLER_247_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_247_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_247_1277 ();
 FILLER_ASAP7_75t_R FILLER_247_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_248_172 ();
 DECAPx10_ASAP7_75t_R FILLER_248_194 ();
 DECAPx10_ASAP7_75t_R FILLER_248_216 ();
 DECAPx10_ASAP7_75t_R FILLER_248_238 ();
 DECAPx6_ASAP7_75t_R FILLER_248_260 ();
 DECAPx1_ASAP7_75t_R FILLER_248_288 ();
 DECAPx1_ASAP7_75t_R FILLER_248_300 ();
 FILLER_ASAP7_75t_R FILLER_248_328 ();
 DECAPx6_ASAP7_75t_R FILLER_248_350 ();
 DECAPx1_ASAP7_75t_R FILLER_248_364 ();
 DECAPx2_ASAP7_75t_R FILLER_248_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_382 ();
 DECAPx1_ASAP7_75t_R FILLER_248_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_405 ();
 DECAPx1_ASAP7_75t_R FILLER_248_420 ();
 DECAPx2_ASAP7_75t_R FILLER_248_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_437 ();
 DECAPx1_ASAP7_75t_R FILLER_248_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_448 ();
 FILLER_ASAP7_75t_R FILLER_248_455 ();
 DECAPx2_ASAP7_75t_R FILLER_248_471 ();
 FILLER_ASAP7_75t_R FILLER_248_477 ();
 DECAPx10_ASAP7_75t_R FILLER_248_495 ();
 DECAPx10_ASAP7_75t_R FILLER_248_517 ();
 DECAPx10_ASAP7_75t_R FILLER_248_539 ();
 DECAPx10_ASAP7_75t_R FILLER_248_561 ();
 DECAPx10_ASAP7_75t_R FILLER_248_583 ();
 DECAPx10_ASAP7_75t_R FILLER_248_605 ();
 DECAPx1_ASAP7_75t_R FILLER_248_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_631 ();
 DECAPx6_ASAP7_75t_R FILLER_248_634 ();
 DECAPx1_ASAP7_75t_R FILLER_248_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_652 ();
 DECAPx10_ASAP7_75t_R FILLER_248_656 ();
 DECAPx10_ASAP7_75t_R FILLER_248_684 ();
 DECAPx6_ASAP7_75t_R FILLER_248_706 ();
 DECAPx1_ASAP7_75t_R FILLER_248_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_724 ();
 DECAPx6_ASAP7_75t_R FILLER_248_746 ();
 DECAPx1_ASAP7_75t_R FILLER_248_760 ();
 DECAPx2_ASAP7_75t_R FILLER_248_770 ();
 FILLER_ASAP7_75t_R FILLER_248_776 ();
 DECAPx10_ASAP7_75t_R FILLER_248_799 ();
 DECAPx2_ASAP7_75t_R FILLER_248_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_834 ();
 DECAPx1_ASAP7_75t_R FILLER_248_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_847 ();
 FILLER_ASAP7_75t_R FILLER_248_856 ();
 FILLER_ASAP7_75t_R FILLER_248_866 ();
 DECAPx10_ASAP7_75t_R FILLER_248_871 ();
 FILLER_ASAP7_75t_R FILLER_248_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_895 ();
 DECAPx4_ASAP7_75t_R FILLER_248_903 ();
 FILLER_ASAP7_75t_R FILLER_248_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_915 ();
 DECAPx6_ASAP7_75t_R FILLER_248_924 ();
 DECAPx4_ASAP7_75t_R FILLER_248_945 ();
 FILLER_ASAP7_75t_R FILLER_248_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_957 ();
 DECAPx4_ASAP7_75t_R FILLER_248_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_976 ();
 DECAPx10_ASAP7_75t_R FILLER_248_991 ();
 DECAPx6_ASAP7_75t_R FILLER_248_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_248_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_249_172 ();
 DECAPx10_ASAP7_75t_R FILLER_249_194 ();
 DECAPx10_ASAP7_75t_R FILLER_249_216 ();
 DECAPx10_ASAP7_75t_R FILLER_249_238 ();
 DECAPx10_ASAP7_75t_R FILLER_249_260 ();
 FILLER_ASAP7_75t_R FILLER_249_288 ();
 DECAPx10_ASAP7_75t_R FILLER_249_302 ();
 DECAPx4_ASAP7_75t_R FILLER_249_324 ();
 FILLER_ASAP7_75t_R FILLER_249_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_342 ();
 DECAPx10_ASAP7_75t_R FILLER_249_349 ();
 DECAPx10_ASAP7_75t_R FILLER_249_371 ();
 DECAPx6_ASAP7_75t_R FILLER_249_393 ();
 DECAPx1_ASAP7_75t_R FILLER_249_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_411 ();
 DECAPx2_ASAP7_75t_R FILLER_249_426 ();
 DECAPx10_ASAP7_75t_R FILLER_249_456 ();
 DECAPx10_ASAP7_75t_R FILLER_249_484 ();
 DECAPx10_ASAP7_75t_R FILLER_249_506 ();
 DECAPx10_ASAP7_75t_R FILLER_249_528 ();
 DECAPx10_ASAP7_75t_R FILLER_249_550 ();
 DECAPx10_ASAP7_75t_R FILLER_249_572 ();
 DECAPx10_ASAP7_75t_R FILLER_249_594 ();
 DECAPx4_ASAP7_75t_R FILLER_249_616 ();
 FILLER_ASAP7_75t_R FILLER_249_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_628 ();
 DECAPx4_ASAP7_75t_R FILLER_249_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_713 ();
 DECAPx2_ASAP7_75t_R FILLER_249_722 ();
 FILLER_ASAP7_75t_R FILLER_249_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_730 ();
 DECAPx1_ASAP7_75t_R FILLER_249_747 ();
 DECAPx2_ASAP7_75t_R FILLER_249_759 ();
 FILLER_ASAP7_75t_R FILLER_249_765 ();
 DECAPx1_ASAP7_75t_R FILLER_249_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_782 ();
 DECAPx1_ASAP7_75t_R FILLER_249_789 ();
 DECAPx2_ASAP7_75t_R FILLER_249_799 ();
 DECAPx2_ASAP7_75t_R FILLER_249_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_852 ();
 DECAPx4_ASAP7_75t_R FILLER_249_874 ();
 FILLER_ASAP7_75t_R FILLER_249_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_886 ();
 DECAPx10_ASAP7_75t_R FILLER_249_891 ();
 DECAPx1_ASAP7_75t_R FILLER_249_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_955 ();
 DECAPx10_ASAP7_75t_R FILLER_249_977 ();
 FILLER_ASAP7_75t_R FILLER_249_999 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1004 ();
 FILLER_ASAP7_75t_R FILLER_249_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1049 ();
 FILLER_ASAP7_75t_R FILLER_249_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_249_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_249_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_250_172 ();
 DECAPx10_ASAP7_75t_R FILLER_250_194 ();
 DECAPx10_ASAP7_75t_R FILLER_250_216 ();
 DECAPx10_ASAP7_75t_R FILLER_250_238 ();
 DECAPx10_ASAP7_75t_R FILLER_250_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_296 ();
 DECAPx2_ASAP7_75t_R FILLER_250_305 ();
 FILLER_ASAP7_75t_R FILLER_250_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_313 ();
 DECAPx4_ASAP7_75t_R FILLER_250_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_334 ();
 DECAPx10_ASAP7_75t_R FILLER_250_341 ();
 DECAPx6_ASAP7_75t_R FILLER_250_363 ();
 DECAPx1_ASAP7_75t_R FILLER_250_377 ();
 DECAPx10_ASAP7_75t_R FILLER_250_393 ();
 FILLER_ASAP7_75t_R FILLER_250_415 ();
 DECAPx6_ASAP7_75t_R FILLER_250_423 ();
 FILLER_ASAP7_75t_R FILLER_250_437 ();
 DECAPx6_ASAP7_75t_R FILLER_250_446 ();
 FILLER_ASAP7_75t_R FILLER_250_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_462 ();
 DECAPx2_ASAP7_75t_R FILLER_250_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_475 ();
 DECAPx1_ASAP7_75t_R FILLER_250_482 ();
 DECAPx10_ASAP7_75t_R FILLER_250_506 ();
 DECAPx10_ASAP7_75t_R FILLER_250_528 ();
 DECAPx10_ASAP7_75t_R FILLER_250_550 ();
 DECAPx10_ASAP7_75t_R FILLER_250_572 ();
 DECAPx6_ASAP7_75t_R FILLER_250_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_608 ();
 DECAPx4_ASAP7_75t_R FILLER_250_620 ();
 FILLER_ASAP7_75t_R FILLER_250_630 ();
 DECAPx1_ASAP7_75t_R FILLER_250_634 ();
 DECAPx6_ASAP7_75t_R FILLER_250_646 ();
 FILLER_ASAP7_75t_R FILLER_250_660 ();
 DECAPx1_ASAP7_75t_R FILLER_250_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_674 ();
 DECAPx4_ASAP7_75t_R FILLER_250_678 ();
 DECAPx10_ASAP7_75t_R FILLER_250_696 ();
 DECAPx6_ASAP7_75t_R FILLER_250_718 ();
 FILLER_ASAP7_75t_R FILLER_250_732 ();
 DECAPx2_ASAP7_75t_R FILLER_250_745 ();
 FILLER_ASAP7_75t_R FILLER_250_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_753 ();
 DECAPx6_ASAP7_75t_R FILLER_250_783 ();
 DECAPx1_ASAP7_75t_R FILLER_250_797 ();
 DECAPx10_ASAP7_75t_R FILLER_250_822 ();
 DECAPx10_ASAP7_75t_R FILLER_250_844 ();
 DECAPx4_ASAP7_75t_R FILLER_250_866 ();
 DECAPx6_ASAP7_75t_R FILLER_250_884 ();
 DECAPx1_ASAP7_75t_R FILLER_250_898 ();
 DECAPx10_ASAP7_75t_R FILLER_250_910 ();
 DECAPx2_ASAP7_75t_R FILLER_250_932 ();
 DECAPx10_ASAP7_75t_R FILLER_250_959 ();
 DECAPx1_ASAP7_75t_R FILLER_250_981 ();
 DECAPx4_ASAP7_75t_R FILLER_250_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1009 ();
 FILLER_ASAP7_75t_R FILLER_250_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1033 ();
 FILLER_ASAP7_75t_R FILLER_250_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_250_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_251_172 ();
 DECAPx10_ASAP7_75t_R FILLER_251_194 ();
 DECAPx10_ASAP7_75t_R FILLER_251_216 ();
 DECAPx10_ASAP7_75t_R FILLER_251_238 ();
 DECAPx4_ASAP7_75t_R FILLER_251_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_270 ();
 DECAPx6_ASAP7_75t_R FILLER_251_279 ();
 FILLER_ASAP7_75t_R FILLER_251_293 ();
 DECAPx1_ASAP7_75t_R FILLER_251_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_306 ();
 DECAPx2_ASAP7_75t_R FILLER_251_313 ();
 FILLER_ASAP7_75t_R FILLER_251_319 ();
 DECAPx10_ASAP7_75t_R FILLER_251_329 ();
 FILLER_ASAP7_75t_R FILLER_251_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_353 ();
 DECAPx6_ASAP7_75t_R FILLER_251_360 ();
 DECAPx4_ASAP7_75t_R FILLER_251_393 ();
 DECAPx10_ASAP7_75t_R FILLER_251_409 ();
 DECAPx10_ASAP7_75t_R FILLER_251_431 ();
 DECAPx2_ASAP7_75t_R FILLER_251_453 ();
 FILLER_ASAP7_75t_R FILLER_251_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_461 ();
 FILLER_ASAP7_75t_R FILLER_251_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_474 ();
 DECAPx10_ASAP7_75t_R FILLER_251_481 ();
 DECAPx10_ASAP7_75t_R FILLER_251_503 ();
 DECAPx10_ASAP7_75t_R FILLER_251_525 ();
 DECAPx10_ASAP7_75t_R FILLER_251_547 ();
 DECAPx10_ASAP7_75t_R FILLER_251_569 ();
 DECAPx2_ASAP7_75t_R FILLER_251_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_597 ();
 FILLER_ASAP7_75t_R FILLER_251_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_628 ();
 FILLER_ASAP7_75t_R FILLER_251_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_638 ();
 DECAPx6_ASAP7_75t_R FILLER_251_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_656 ();
 DECAPx10_ASAP7_75t_R FILLER_251_678 ();
 DECAPx4_ASAP7_75t_R FILLER_251_700 ();
 DECAPx4_ASAP7_75t_R FILLER_251_713 ();
 FILLER_ASAP7_75t_R FILLER_251_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_764 ();
 DECAPx10_ASAP7_75t_R FILLER_251_768 ();
 DECAPx6_ASAP7_75t_R FILLER_251_790 ();
 FILLER_ASAP7_75t_R FILLER_251_804 ();
 DECAPx10_ASAP7_75t_R FILLER_251_814 ();
 DECAPx10_ASAP7_75t_R FILLER_251_836 ();
 DECAPx1_ASAP7_75t_R FILLER_251_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_862 ();
 DECAPx1_ASAP7_75t_R FILLER_251_867 ();
 DECAPx1_ASAP7_75t_R FILLER_251_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_903 ();
 DECAPx10_ASAP7_75t_R FILLER_251_907 ();
 DECAPx10_ASAP7_75t_R FILLER_251_929 ();
 DECAPx10_ASAP7_75t_R FILLER_251_951 ();
 DECAPx4_ASAP7_75t_R FILLER_251_973 ();
 FILLER_ASAP7_75t_R FILLER_251_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_985 ();
 FILLER_ASAP7_75t_R FILLER_251_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1020 ();
 FILLER_ASAP7_75t_R FILLER_251_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_252_172 ();
 DECAPx10_ASAP7_75t_R FILLER_252_194 ();
 DECAPx10_ASAP7_75t_R FILLER_252_216 ();
 DECAPx10_ASAP7_75t_R FILLER_252_238 ();
 DECAPx6_ASAP7_75t_R FILLER_252_260 ();
 DECAPx1_ASAP7_75t_R FILLER_252_274 ();
 DECAPx2_ASAP7_75t_R FILLER_252_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_294 ();
 FILLER_ASAP7_75t_R FILLER_252_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_346 ();
 DECAPx2_ASAP7_75t_R FILLER_252_362 ();
 FILLER_ASAP7_75t_R FILLER_252_368 ();
 FILLER_ASAP7_75t_R FILLER_252_376 ();
 FILLER_ASAP7_75t_R FILLER_252_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_388 ();
 DECAPx2_ASAP7_75t_R FILLER_252_395 ();
 FILLER_ASAP7_75t_R FILLER_252_401 ();
 DECAPx2_ASAP7_75t_R FILLER_252_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_426 ();
 DECAPx10_ASAP7_75t_R FILLER_252_439 ();
 DECAPx2_ASAP7_75t_R FILLER_252_461 ();
 FILLER_ASAP7_75t_R FILLER_252_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_469 ();
 DECAPx10_ASAP7_75t_R FILLER_252_506 ();
 DECAPx10_ASAP7_75t_R FILLER_252_528 ();
 DECAPx10_ASAP7_75t_R FILLER_252_550 ();
 DECAPx10_ASAP7_75t_R FILLER_252_572 ();
 DECAPx6_ASAP7_75t_R FILLER_252_594 ();
 FILLER_ASAP7_75t_R FILLER_252_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_610 ();
 FILLER_ASAP7_75t_R FILLER_252_642 ();
 DECAPx1_ASAP7_75t_R FILLER_252_655 ();
 DECAPx6_ASAP7_75t_R FILLER_252_665 ();
 DECAPx1_ASAP7_75t_R FILLER_252_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_683 ();
 DECAPx1_ASAP7_75t_R FILLER_252_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_699 ();
 FILLER_ASAP7_75t_R FILLER_252_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_723 ();
 FILLER_ASAP7_75t_R FILLER_252_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_747 ();
 DECAPx10_ASAP7_75t_R FILLER_252_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_791 ();
 DECAPx10_ASAP7_75t_R FILLER_252_803 ();
 DECAPx4_ASAP7_75t_R FILLER_252_825 ();
 FILLER_ASAP7_75t_R FILLER_252_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_837 ();
 FILLER_ASAP7_75t_R FILLER_252_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_848 ();
 FILLER_ASAP7_75t_R FILLER_252_880 ();
 DECAPx10_ASAP7_75t_R FILLER_252_903 ();
 DECAPx10_ASAP7_75t_R FILLER_252_925 ();
 FILLER_ASAP7_75t_R FILLER_252_947 ();
 DECAPx2_ASAP7_75t_R FILLER_252_966 ();
 DECAPx1_ASAP7_75t_R FILLER_252_986 ();
 DECAPx2_ASAP7_75t_R FILLER_252_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_252_1022 ();
 FILLER_ASAP7_75t_R FILLER_252_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1285 ();
 FILLER_ASAP7_75t_R FILLER_252_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_253_172 ();
 DECAPx10_ASAP7_75t_R FILLER_253_194 ();
 DECAPx10_ASAP7_75t_R FILLER_253_216 ();
 DECAPx10_ASAP7_75t_R FILLER_253_238 ();
 DECAPx10_ASAP7_75t_R FILLER_253_260 ();
 DECAPx6_ASAP7_75t_R FILLER_253_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_296 ();
 DECAPx6_ASAP7_75t_R FILLER_253_313 ();
 DECAPx2_ASAP7_75t_R FILLER_253_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_333 ();
 DECAPx2_ASAP7_75t_R FILLER_253_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_346 ();
 DECAPx6_ASAP7_75t_R FILLER_253_355 ();
 DECAPx1_ASAP7_75t_R FILLER_253_375 ();
 DECAPx1_ASAP7_75t_R FILLER_253_386 ();
 DECAPx1_ASAP7_75t_R FILLER_253_396 ();
 FILLER_ASAP7_75t_R FILLER_253_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_442 ();
 DECAPx2_ASAP7_75t_R FILLER_253_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_466 ();
 FILLER_ASAP7_75t_R FILLER_253_473 ();
 FILLER_ASAP7_75t_R FILLER_253_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_483 ();
 DECAPx10_ASAP7_75t_R FILLER_253_494 ();
 DECAPx10_ASAP7_75t_R FILLER_253_516 ();
 DECAPx10_ASAP7_75t_R FILLER_253_538 ();
 DECAPx10_ASAP7_75t_R FILLER_253_560 ();
 DECAPx10_ASAP7_75t_R FILLER_253_582 ();
 DECAPx10_ASAP7_75t_R FILLER_253_604 ();
 DECAPx4_ASAP7_75t_R FILLER_253_626 ();
 DECAPx6_ASAP7_75t_R FILLER_253_657 ();
 DECAPx1_ASAP7_75t_R FILLER_253_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_675 ();
 FILLER_ASAP7_75t_R FILLER_253_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_699 ();
 DECAPx6_ASAP7_75t_R FILLER_253_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_728 ();
 DECAPx6_ASAP7_75t_R FILLER_253_735 ();
 FILLER_ASAP7_75t_R FILLER_253_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_751 ();
 DECAPx2_ASAP7_75t_R FILLER_253_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_764 ();
 DECAPx6_ASAP7_75t_R FILLER_253_807 ();
 DECAPx1_ASAP7_75t_R FILLER_253_829 ();
 DECAPx2_ASAP7_75t_R FILLER_253_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_868 ();
 DECAPx6_ASAP7_75t_R FILLER_253_875 ();
 DECAPx1_ASAP7_75t_R FILLER_253_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_893 ();
 FILLER_ASAP7_75t_R FILLER_253_901 ();
 FILLER_ASAP7_75t_R FILLER_253_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_929 ();
 DECAPx2_ASAP7_75t_R FILLER_253_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_998 ();
 DECAPx6_ASAP7_75t_R FILLER_253_1013 ();
 FILLER_ASAP7_75t_R FILLER_253_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_253_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_253_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_254_172 ();
 DECAPx10_ASAP7_75t_R FILLER_254_194 ();
 DECAPx10_ASAP7_75t_R FILLER_254_216 ();
 DECAPx10_ASAP7_75t_R FILLER_254_238 ();
 DECAPx10_ASAP7_75t_R FILLER_254_260 ();
 DECAPx10_ASAP7_75t_R FILLER_254_282 ();
 DECAPx10_ASAP7_75t_R FILLER_254_310 ();
 DECAPx2_ASAP7_75t_R FILLER_254_332 ();
 FILLER_ASAP7_75t_R FILLER_254_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_340 ();
 DECAPx6_ASAP7_75t_R FILLER_254_353 ();
 FILLER_ASAP7_75t_R FILLER_254_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_369 ();
 FILLER_ASAP7_75t_R FILLER_254_377 ();
 DECAPx6_ASAP7_75t_R FILLER_254_385 ();
 FILLER_ASAP7_75t_R FILLER_254_399 ();
 DECAPx10_ASAP7_75t_R FILLER_254_415 ();
 FILLER_ASAP7_75t_R FILLER_254_443 ();
 DECAPx2_ASAP7_75t_R FILLER_254_457 ();
 FILLER_ASAP7_75t_R FILLER_254_463 ();
 DECAPx1_ASAP7_75t_R FILLER_254_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_475 ();
 DECAPx10_ASAP7_75t_R FILLER_254_484 ();
 DECAPx10_ASAP7_75t_R FILLER_254_506 ();
 DECAPx10_ASAP7_75t_R FILLER_254_528 ();
 DECAPx10_ASAP7_75t_R FILLER_254_550 ();
 DECAPx10_ASAP7_75t_R FILLER_254_572 ();
 DECAPx4_ASAP7_75t_R FILLER_254_594 ();
 DECAPx2_ASAP7_75t_R FILLER_254_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_631 ();
 DECAPx2_ASAP7_75t_R FILLER_254_634 ();
 FILLER_ASAP7_75t_R FILLER_254_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_642 ();
 FILLER_ASAP7_75t_R FILLER_254_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_651 ();
 DECAPx2_ASAP7_75t_R FILLER_254_676 ();
 FILLER_ASAP7_75t_R FILLER_254_682 ();
 DECAPx10_ASAP7_75t_R FILLER_254_690 ();
 DECAPx10_ASAP7_75t_R FILLER_254_712 ();
 DECAPx10_ASAP7_75t_R FILLER_254_734 ();
 DECAPx2_ASAP7_75t_R FILLER_254_756 ();
 FILLER_ASAP7_75t_R FILLER_254_776 ();
 DECAPx2_ASAP7_75t_R FILLER_254_781 ();
 FILLER_ASAP7_75t_R FILLER_254_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_789 ();
 DECAPx4_ASAP7_75t_R FILLER_254_796 ();
 DECAPx4_ASAP7_75t_R FILLER_254_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_833 ();
 DECAPx6_ASAP7_75t_R FILLER_254_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_854 ();
 DECAPx4_ASAP7_75t_R FILLER_254_862 ();
 FILLER_ASAP7_75t_R FILLER_254_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_874 ();
 FILLER_ASAP7_75t_R FILLER_254_899 ();
 DECAPx4_ASAP7_75t_R FILLER_254_923 ();
 DECAPx10_ASAP7_75t_R FILLER_254_944 ();
 DECAPx6_ASAP7_75t_R FILLER_254_966 ();
 FILLER_ASAP7_75t_R FILLER_254_980 ();
 DECAPx10_ASAP7_75t_R FILLER_254_996 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_254_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_255_172 ();
 DECAPx10_ASAP7_75t_R FILLER_255_194 ();
 DECAPx10_ASAP7_75t_R FILLER_255_216 ();
 DECAPx10_ASAP7_75t_R FILLER_255_238 ();
 DECAPx10_ASAP7_75t_R FILLER_255_260 ();
 DECAPx4_ASAP7_75t_R FILLER_255_282 ();
 FILLER_ASAP7_75t_R FILLER_255_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_322 ();
 DECAPx10_ASAP7_75t_R FILLER_255_331 ();
 DECAPx10_ASAP7_75t_R FILLER_255_353 ();
 DECAPx1_ASAP7_75t_R FILLER_255_375 ();
 DECAPx2_ASAP7_75t_R FILLER_255_387 ();
 FILLER_ASAP7_75t_R FILLER_255_405 ();
 DECAPx6_ASAP7_75t_R FILLER_255_415 ();
 DECAPx1_ASAP7_75t_R FILLER_255_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_433 ();
 DECAPx10_ASAP7_75t_R FILLER_255_441 ();
 DECAPx10_ASAP7_75t_R FILLER_255_463 ();
 FILLER_ASAP7_75t_R FILLER_255_485 ();
 DECAPx10_ASAP7_75t_R FILLER_255_497 ();
 DECAPx10_ASAP7_75t_R FILLER_255_519 ();
 DECAPx10_ASAP7_75t_R FILLER_255_541 ();
 DECAPx10_ASAP7_75t_R FILLER_255_563 ();
 DECAPx10_ASAP7_75t_R FILLER_255_585 ();
 DECAPx4_ASAP7_75t_R FILLER_255_607 ();
 DECAPx6_ASAP7_75t_R FILLER_255_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_642 ();
 DECAPx1_ASAP7_75t_R FILLER_255_649 ();
 DECAPx10_ASAP7_75t_R FILLER_255_667 ();
 DECAPx4_ASAP7_75t_R FILLER_255_689 ();
 FILLER_ASAP7_75t_R FILLER_255_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_701 ();
 DECAPx4_ASAP7_75t_R FILLER_255_710 ();
 DECAPx2_ASAP7_75t_R FILLER_255_731 ();
 FILLER_ASAP7_75t_R FILLER_255_737 ();
 DECAPx10_ASAP7_75t_R FILLER_255_750 ();
 DECAPx10_ASAP7_75t_R FILLER_255_772 ();
 DECAPx6_ASAP7_75t_R FILLER_255_794 ();
 DECAPx2_ASAP7_75t_R FILLER_255_808 ();
 DECAPx10_ASAP7_75t_R FILLER_255_828 ();
 DECAPx4_ASAP7_75t_R FILLER_255_850 ();
 FILLER_ASAP7_75t_R FILLER_255_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_862 ();
 DECAPx10_ASAP7_75t_R FILLER_255_866 ();
 DECAPx4_ASAP7_75t_R FILLER_255_888 ();
 FILLER_ASAP7_75t_R FILLER_255_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_900 ();
 FILLER_ASAP7_75t_R FILLER_255_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_917 ();
 DECAPx10_ASAP7_75t_R FILLER_255_945 ();
 DECAPx6_ASAP7_75t_R FILLER_255_967 ();
 FILLER_ASAP7_75t_R FILLER_255_981 ();
 DECAPx6_ASAP7_75t_R FILLER_255_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_255_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_255_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_255_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_256_172 ();
 DECAPx10_ASAP7_75t_R FILLER_256_194 ();
 DECAPx10_ASAP7_75t_R FILLER_256_216 ();
 DECAPx10_ASAP7_75t_R FILLER_256_238 ();
 DECAPx10_ASAP7_75t_R FILLER_256_260 ();
 DECAPx10_ASAP7_75t_R FILLER_256_282 ();
 DECAPx6_ASAP7_75t_R FILLER_256_304 ();
 FILLER_ASAP7_75t_R FILLER_256_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_320 ();
 FILLER_ASAP7_75t_R FILLER_256_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_337 ();
 DECAPx4_ASAP7_75t_R FILLER_256_351 ();
 DECAPx10_ASAP7_75t_R FILLER_256_371 ();
 DECAPx1_ASAP7_75t_R FILLER_256_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_420 ();
 DECAPx2_ASAP7_75t_R FILLER_256_429 ();
 FILLER_ASAP7_75t_R FILLER_256_435 ();
 FILLER_ASAP7_75t_R FILLER_256_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_445 ();
 DECAPx2_ASAP7_75t_R FILLER_256_452 ();
 FILLER_ASAP7_75t_R FILLER_256_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_468 ();
 DECAPx2_ASAP7_75t_R FILLER_256_475 ();
 DECAPx10_ASAP7_75t_R FILLER_256_491 ();
 DECAPx10_ASAP7_75t_R FILLER_256_513 ();
 DECAPx10_ASAP7_75t_R FILLER_256_535 ();
 DECAPx10_ASAP7_75t_R FILLER_256_557 ();
 DECAPx10_ASAP7_75t_R FILLER_256_579 ();
 DECAPx6_ASAP7_75t_R FILLER_256_601 ();
 DECAPx2_ASAP7_75t_R FILLER_256_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_621 ();
 DECAPx1_ASAP7_75t_R FILLER_256_628 ();
 DECAPx2_ASAP7_75t_R FILLER_256_634 ();
 FILLER_ASAP7_75t_R FILLER_256_640 ();
 DECAPx6_ASAP7_75t_R FILLER_256_657 ();
 FILLER_ASAP7_75t_R FILLER_256_671 ();
 DECAPx1_ASAP7_75t_R FILLER_256_687 ();
 FILLER_ASAP7_75t_R FILLER_256_754 ();
 DECAPx10_ASAP7_75t_R FILLER_256_764 ();
 DECAPx2_ASAP7_75t_R FILLER_256_786 ();
 FILLER_ASAP7_75t_R FILLER_256_792 ();
 DECAPx6_ASAP7_75t_R FILLER_256_838 ();
 DECAPx1_ASAP7_75t_R FILLER_256_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_856 ();
 DECAPx6_ASAP7_75t_R FILLER_256_865 ();
 DECAPx2_ASAP7_75t_R FILLER_256_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_885 ();
 DECAPx10_ASAP7_75t_R FILLER_256_910 ();
 DECAPx2_ASAP7_75t_R FILLER_256_932 ();
 DECAPx2_ASAP7_75t_R FILLER_256_945 ();
 FILLER_ASAP7_75t_R FILLER_256_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_953 ();
 FILLER_ASAP7_75t_R FILLER_256_965 ();
 DECAPx10_ASAP7_75t_R FILLER_256_973 ();
 DECAPx6_ASAP7_75t_R FILLER_256_995 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_256_1034 ();
 FILLER_ASAP7_75t_R FILLER_256_1040 ();
 FILLER_ASAP7_75t_R FILLER_256_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_256_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_257_172 ();
 DECAPx10_ASAP7_75t_R FILLER_257_194 ();
 DECAPx10_ASAP7_75t_R FILLER_257_216 ();
 DECAPx10_ASAP7_75t_R FILLER_257_238 ();
 DECAPx10_ASAP7_75t_R FILLER_257_260 ();
 DECAPx2_ASAP7_75t_R FILLER_257_282 ();
 DECAPx6_ASAP7_75t_R FILLER_257_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_335 ();
 DECAPx10_ASAP7_75t_R FILLER_257_347 ();
 DECAPx4_ASAP7_75t_R FILLER_257_369 ();
 FILLER_ASAP7_75t_R FILLER_257_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_388 ();
 DECAPx6_ASAP7_75t_R FILLER_257_403 ();
 DECAPx1_ASAP7_75t_R FILLER_257_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_443 ();
 FILLER_ASAP7_75t_R FILLER_257_451 ();
 FILLER_ASAP7_75t_R FILLER_257_460 ();
 FILLER_ASAP7_75t_R FILLER_257_468 ();
 FILLER_ASAP7_75t_R FILLER_257_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_479 ();
 DECAPx10_ASAP7_75t_R FILLER_257_488 ();
 DECAPx10_ASAP7_75t_R FILLER_257_510 ();
 DECAPx10_ASAP7_75t_R FILLER_257_532 ();
 DECAPx10_ASAP7_75t_R FILLER_257_554 ();
 DECAPx10_ASAP7_75t_R FILLER_257_576 ();
 DECAPx4_ASAP7_75t_R FILLER_257_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_640 ();
 DECAPx1_ASAP7_75t_R FILLER_257_695 ();
 FILLER_ASAP7_75t_R FILLER_257_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_716 ();
 DECAPx4_ASAP7_75t_R FILLER_257_723 ();
 FILLER_ASAP7_75t_R FILLER_257_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_735 ();
 DECAPx2_ASAP7_75t_R FILLER_257_742 ();
 FILLER_ASAP7_75t_R FILLER_257_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_750 ();
 DECAPx2_ASAP7_75t_R FILLER_257_772 ();
 DECAPx4_ASAP7_75t_R FILLER_257_786 ();
 DECAPx6_ASAP7_75t_R FILLER_257_807 ();
 DECAPx2_ASAP7_75t_R FILLER_257_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_827 ();
 DECAPx1_ASAP7_75t_R FILLER_257_849 ();
 DECAPx10_ASAP7_75t_R FILLER_257_874 ();
 DECAPx6_ASAP7_75t_R FILLER_257_896 ();
 FILLER_ASAP7_75t_R FILLER_257_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_912 ();
 DECAPx10_ASAP7_75t_R FILLER_257_919 ();
 DECAPx4_ASAP7_75t_R FILLER_257_941 ();
 DECAPx10_ASAP7_75t_R FILLER_257_972 ();
 DECAPx1_ASAP7_75t_R FILLER_257_994 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_257_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_257_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_257_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_257_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_258_172 ();
 DECAPx10_ASAP7_75t_R FILLER_258_194 ();
 DECAPx10_ASAP7_75t_R FILLER_258_216 ();
 DECAPx10_ASAP7_75t_R FILLER_258_238 ();
 DECAPx10_ASAP7_75t_R FILLER_258_260 ();
 DECAPx10_ASAP7_75t_R FILLER_258_282 ();
 DECAPx10_ASAP7_75t_R FILLER_258_304 ();
 DECAPx6_ASAP7_75t_R FILLER_258_326 ();
 FILLER_ASAP7_75t_R FILLER_258_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_364 ();
 DECAPx1_ASAP7_75t_R FILLER_258_373 ();
 DECAPx4_ASAP7_75t_R FILLER_258_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_399 ();
 DECAPx1_ASAP7_75t_R FILLER_258_412 ();
 DECAPx1_ASAP7_75t_R FILLER_258_428 ();
 DECAPx1_ASAP7_75t_R FILLER_258_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_470 ();
 DECAPx10_ASAP7_75t_R FILLER_258_477 ();
 DECAPx10_ASAP7_75t_R FILLER_258_499 ();
 DECAPx10_ASAP7_75t_R FILLER_258_521 ();
 DECAPx10_ASAP7_75t_R FILLER_258_543 ();
 DECAPx10_ASAP7_75t_R FILLER_258_565 ();
 DECAPx10_ASAP7_75t_R FILLER_258_587 ();
 DECAPx6_ASAP7_75t_R FILLER_258_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_623 ();
 DECAPx1_ASAP7_75t_R FILLER_258_634 ();
 DECAPx1_ASAP7_75t_R FILLER_258_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_650 ();
 DECAPx10_ASAP7_75t_R FILLER_258_661 ();
 DECAPx10_ASAP7_75t_R FILLER_258_683 ();
 DECAPx10_ASAP7_75t_R FILLER_258_705 ();
 DECAPx10_ASAP7_75t_R FILLER_258_727 ();
 DECAPx1_ASAP7_75t_R FILLER_258_749 ();
 FILLER_ASAP7_75t_R FILLER_258_759 ();
 DECAPx2_ASAP7_75t_R FILLER_258_764 ();
 FILLER_ASAP7_75t_R FILLER_258_770 ();
 DECAPx6_ASAP7_75t_R FILLER_258_814 ();
 DECAPx1_ASAP7_75t_R FILLER_258_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_832 ();
 DECAPx10_ASAP7_75t_R FILLER_258_870 ();
 FILLER_ASAP7_75t_R FILLER_258_892 ();
 DECAPx2_ASAP7_75t_R FILLER_258_901 ();
 FILLER_ASAP7_75t_R FILLER_258_910 ();
 DECAPx1_ASAP7_75t_R FILLER_258_926 ();
 DECAPx1_ASAP7_75t_R FILLER_258_933 ();
 DECAPx2_ASAP7_75t_R FILLER_258_961 ();
 FILLER_ASAP7_75t_R FILLER_258_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_969 ();
 DECAPx2_ASAP7_75t_R FILLER_258_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_987 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_258_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_259_172 ();
 DECAPx10_ASAP7_75t_R FILLER_259_194 ();
 DECAPx10_ASAP7_75t_R FILLER_259_216 ();
 DECAPx10_ASAP7_75t_R FILLER_259_238 ();
 DECAPx10_ASAP7_75t_R FILLER_259_260 ();
 DECAPx10_ASAP7_75t_R FILLER_259_282 ();
 DECAPx4_ASAP7_75t_R FILLER_259_304 ();
 FILLER_ASAP7_75t_R FILLER_259_314 ();
 DECAPx6_ASAP7_75t_R FILLER_259_326 ();
 FILLER_ASAP7_75t_R FILLER_259_340 ();
 FILLER_ASAP7_75t_R FILLER_259_355 ();
 DECAPx4_ASAP7_75t_R FILLER_259_369 ();
 DECAPx6_ASAP7_75t_R FILLER_259_391 ();
 FILLER_ASAP7_75t_R FILLER_259_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_419 ();
 DECAPx10_ASAP7_75t_R FILLER_259_426 ();
 DECAPx6_ASAP7_75t_R FILLER_259_448 ();
 DECAPx1_ASAP7_75t_R FILLER_259_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_466 ();
 FILLER_ASAP7_75t_R FILLER_259_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_477 ();
 DECAPx10_ASAP7_75t_R FILLER_259_488 ();
 DECAPx10_ASAP7_75t_R FILLER_259_510 ();
 DECAPx10_ASAP7_75t_R FILLER_259_532 ();
 DECAPx10_ASAP7_75t_R FILLER_259_554 ();
 DECAPx10_ASAP7_75t_R FILLER_259_576 ();
 DECAPx10_ASAP7_75t_R FILLER_259_598 ();
 DECAPx4_ASAP7_75t_R FILLER_259_620 ();
 FILLER_ASAP7_75t_R FILLER_259_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_632 ();
 DECAPx10_ASAP7_75t_R FILLER_259_662 ();
 FILLER_ASAP7_75t_R FILLER_259_684 ();
 DECAPx2_ASAP7_75t_R FILLER_259_715 ();
 FILLER_ASAP7_75t_R FILLER_259_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_723 ();
 DECAPx6_ASAP7_75t_R FILLER_259_727 ();
 DECAPx10_ASAP7_75t_R FILLER_259_744 ();
 DECAPx2_ASAP7_75t_R FILLER_259_766 ();
 FILLER_ASAP7_75t_R FILLER_259_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_774 ();
 FILLER_ASAP7_75t_R FILLER_259_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_783 ();
 DECAPx10_ASAP7_75t_R FILLER_259_787 ();
 DECAPx6_ASAP7_75t_R FILLER_259_809 ();
 DECAPx4_ASAP7_75t_R FILLER_259_852 ();
 DECAPx6_ASAP7_75t_R FILLER_259_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_901 ();
 DECAPx1_ASAP7_75t_R FILLER_259_910 ();
 FILLER_ASAP7_75t_R FILLER_259_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_937 ();
 DECAPx4_ASAP7_75t_R FILLER_259_953 ();
 FILLER_ASAP7_75t_R FILLER_259_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_986 ();
 DECAPx6_ASAP7_75t_R FILLER_259_995 ();
 DECAPx1_ASAP7_75t_R FILLER_259_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_259_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_259_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_259_1082 ();
 FILLER_ASAP7_75t_R FILLER_259_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_259_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_259_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_260_172 ();
 DECAPx10_ASAP7_75t_R FILLER_260_194 ();
 DECAPx10_ASAP7_75t_R FILLER_260_216 ();
 DECAPx10_ASAP7_75t_R FILLER_260_238 ();
 DECAPx10_ASAP7_75t_R FILLER_260_260 ();
 DECAPx10_ASAP7_75t_R FILLER_260_282 ();
 DECAPx10_ASAP7_75t_R FILLER_260_304 ();
 DECAPx6_ASAP7_75t_R FILLER_260_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_340 ();
 FILLER_ASAP7_75t_R FILLER_260_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_353 ();
 DECAPx10_ASAP7_75t_R FILLER_260_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_390 ();
 DECAPx2_ASAP7_75t_R FILLER_260_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_405 ();
 DECAPx1_ASAP7_75t_R FILLER_260_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_422 ();
 DECAPx1_ASAP7_75t_R FILLER_260_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_433 ();
 FILLER_ASAP7_75t_R FILLER_260_446 ();
 DECAPx2_ASAP7_75t_R FILLER_260_456 ();
 DECAPx4_ASAP7_75t_R FILLER_260_472 ();
 DECAPx10_ASAP7_75t_R FILLER_260_500 ();
 DECAPx10_ASAP7_75t_R FILLER_260_522 ();
 DECAPx10_ASAP7_75t_R FILLER_260_544 ();
 DECAPx10_ASAP7_75t_R FILLER_260_566 ();
 DECAPx10_ASAP7_75t_R FILLER_260_588 ();
 DECAPx1_ASAP7_75t_R FILLER_260_610 ();
 FILLER_ASAP7_75t_R FILLER_260_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_624 ();
 DECAPx1_ASAP7_75t_R FILLER_260_628 ();
 DECAPx10_ASAP7_75t_R FILLER_260_634 ();
 DECAPx6_ASAP7_75t_R FILLER_260_656 ();
 DECAPx1_ASAP7_75t_R FILLER_260_694 ();
 DECAPx2_ASAP7_75t_R FILLER_260_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_757 ();
 DECAPx10_ASAP7_75t_R FILLER_260_769 ();
 DECAPx6_ASAP7_75t_R FILLER_260_791 ();
 DECAPx2_ASAP7_75t_R FILLER_260_805 ();
 DECAPx2_ASAP7_75t_R FILLER_260_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_847 ();
 DECAPx6_ASAP7_75t_R FILLER_260_851 ();
 DECAPx10_ASAP7_75t_R FILLER_260_907 ();
 DECAPx10_ASAP7_75t_R FILLER_260_929 ();
 DECAPx10_ASAP7_75t_R FILLER_260_951 ();
 DECAPx4_ASAP7_75t_R FILLER_260_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_983 ();
 DECAPx2_ASAP7_75t_R FILLER_260_990 ();
 FILLER_ASAP7_75t_R FILLER_260_996 ();
 DECAPx4_ASAP7_75t_R FILLER_260_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_260_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_260_1280 ();
 FILLER_ASAP7_75t_R FILLER_260_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_261_172 ();
 DECAPx10_ASAP7_75t_R FILLER_261_194 ();
 DECAPx10_ASAP7_75t_R FILLER_261_216 ();
 DECAPx10_ASAP7_75t_R FILLER_261_238 ();
 DECAPx10_ASAP7_75t_R FILLER_261_260 ();
 DECAPx10_ASAP7_75t_R FILLER_261_282 ();
 DECAPx10_ASAP7_75t_R FILLER_261_304 ();
 DECAPx10_ASAP7_75t_R FILLER_261_326 ();
 DECAPx10_ASAP7_75t_R FILLER_261_348 ();
 DECAPx1_ASAP7_75t_R FILLER_261_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_391 ();
 DECAPx4_ASAP7_75t_R FILLER_261_398 ();
 FILLER_ASAP7_75t_R FILLER_261_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_418 ();
 FILLER_ASAP7_75t_R FILLER_261_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_434 ();
 DECAPx2_ASAP7_75t_R FILLER_261_447 ();
 DECAPx10_ASAP7_75t_R FILLER_261_463 ();
 DECAPx10_ASAP7_75t_R FILLER_261_485 ();
 DECAPx10_ASAP7_75t_R FILLER_261_507 ();
 DECAPx10_ASAP7_75t_R FILLER_261_529 ();
 DECAPx10_ASAP7_75t_R FILLER_261_551 ();
 DECAPx10_ASAP7_75t_R FILLER_261_573 ();
 DECAPx4_ASAP7_75t_R FILLER_261_595 ();
 FILLER_ASAP7_75t_R FILLER_261_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_607 ();
 FILLER_ASAP7_75t_R FILLER_261_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_631 ();
 DECAPx2_ASAP7_75t_R FILLER_261_640 ();
 FILLER_ASAP7_75t_R FILLER_261_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_648 ();
 DECAPx2_ASAP7_75t_R FILLER_261_652 ();
 FILLER_ASAP7_75t_R FILLER_261_658 ();
 DECAPx6_ASAP7_75t_R FILLER_261_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_680 ();
 DECAPx2_ASAP7_75t_R FILLER_261_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_701 ();
 DECAPx1_ASAP7_75t_R FILLER_261_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_712 ();
 FILLER_ASAP7_75t_R FILLER_261_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_729 ();
 DECAPx2_ASAP7_75t_R FILLER_261_744 ();
 FILLER_ASAP7_75t_R FILLER_261_750 ();
 DECAPx2_ASAP7_75t_R FILLER_261_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_779 ();
 DECAPx6_ASAP7_75t_R FILLER_261_791 ();
 DECAPx1_ASAP7_75t_R FILLER_261_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_823 ();
 DECAPx10_ASAP7_75t_R FILLER_261_835 ();
 DECAPx10_ASAP7_75t_R FILLER_261_857 ();
 DECAPx2_ASAP7_75t_R FILLER_261_879 ();
 DECAPx10_ASAP7_75t_R FILLER_261_888 ();
 FILLER_ASAP7_75t_R FILLER_261_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_912 ();
 DECAPx10_ASAP7_75t_R FILLER_261_919 ();
 DECAPx10_ASAP7_75t_R FILLER_261_941 ();
 DECAPx10_ASAP7_75t_R FILLER_261_963 ();
 FILLER_ASAP7_75t_R FILLER_261_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1008 ();
 DECAPx4_ASAP7_75t_R FILLER_261_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1027 ();
 DECAPx6_ASAP7_75t_R FILLER_261_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_261_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_261_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_261_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_262_172 ();
 DECAPx10_ASAP7_75t_R FILLER_262_194 ();
 DECAPx10_ASAP7_75t_R FILLER_262_216 ();
 DECAPx10_ASAP7_75t_R FILLER_262_238 ();
 DECAPx10_ASAP7_75t_R FILLER_262_260 ();
 DECAPx10_ASAP7_75t_R FILLER_262_282 ();
 DECAPx10_ASAP7_75t_R FILLER_262_304 ();
 DECAPx10_ASAP7_75t_R FILLER_262_326 ();
 DECAPx10_ASAP7_75t_R FILLER_262_348 ();
 DECAPx2_ASAP7_75t_R FILLER_262_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_376 ();
 DECAPx6_ASAP7_75t_R FILLER_262_385 ();
 FILLER_ASAP7_75t_R FILLER_262_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_413 ();
 DECAPx2_ASAP7_75t_R FILLER_262_430 ();
 DECAPx2_ASAP7_75t_R FILLER_262_444 ();
 FILLER_ASAP7_75t_R FILLER_262_450 ();
 DECAPx10_ASAP7_75t_R FILLER_262_462 ();
 DECAPx10_ASAP7_75t_R FILLER_262_484 ();
 DECAPx10_ASAP7_75t_R FILLER_262_506 ();
 DECAPx10_ASAP7_75t_R FILLER_262_528 ();
 DECAPx10_ASAP7_75t_R FILLER_262_550 ();
 DECAPx10_ASAP7_75t_R FILLER_262_572 ();
 DECAPx6_ASAP7_75t_R FILLER_262_594 ();
 DECAPx1_ASAP7_75t_R FILLER_262_608 ();
 DECAPx2_ASAP7_75t_R FILLER_262_618 ();
 FILLER_ASAP7_75t_R FILLER_262_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_656 ();
 DECAPx10_ASAP7_75t_R FILLER_262_681 ();
 DECAPx1_ASAP7_75t_R FILLER_262_703 ();
 DECAPx10_ASAP7_75t_R FILLER_262_713 ();
 DECAPx6_ASAP7_75t_R FILLER_262_735 ();
 DECAPx2_ASAP7_75t_R FILLER_262_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_755 ();
 DECAPx4_ASAP7_75t_R FILLER_262_762 ();
 FILLER_ASAP7_75t_R FILLER_262_772 ();
 DECAPx1_ASAP7_75t_R FILLER_262_795 ();
 FILLER_ASAP7_75t_R FILLER_262_820 ();
 DECAPx10_ASAP7_75t_R FILLER_262_828 ();
 DECAPx10_ASAP7_75t_R FILLER_262_850 ();
 DECAPx2_ASAP7_75t_R FILLER_262_872 ();
 FILLER_ASAP7_75t_R FILLER_262_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_880 ();
 DECAPx4_ASAP7_75t_R FILLER_262_889 ();
 FILLER_ASAP7_75t_R FILLER_262_899 ();
 FILLER_ASAP7_75t_R FILLER_262_907 ();
 FILLER_ASAP7_75t_R FILLER_262_912 ();
 DECAPx1_ASAP7_75t_R FILLER_262_922 ();
 DECAPx1_ASAP7_75t_R FILLER_262_947 ();
 FILLER_ASAP7_75t_R FILLER_262_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_961 ();
 DECAPx1_ASAP7_75t_R FILLER_262_965 ();
 DECAPx1_ASAP7_75t_R FILLER_262_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_981 ();
 DECAPx1_ASAP7_75t_R FILLER_262_996 ();
 FILLER_ASAP7_75t_R FILLER_262_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1011 ();
 FILLER_ASAP7_75t_R FILLER_262_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_262_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_262_1277 ();
 FILLER_ASAP7_75t_R FILLER_262_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_263_172 ();
 DECAPx10_ASAP7_75t_R FILLER_263_194 ();
 DECAPx10_ASAP7_75t_R FILLER_263_216 ();
 DECAPx10_ASAP7_75t_R FILLER_263_238 ();
 DECAPx10_ASAP7_75t_R FILLER_263_260 ();
 DECAPx10_ASAP7_75t_R FILLER_263_282 ();
 DECAPx10_ASAP7_75t_R FILLER_263_304 ();
 DECAPx10_ASAP7_75t_R FILLER_263_326 ();
 DECAPx10_ASAP7_75t_R FILLER_263_348 ();
 DECAPx10_ASAP7_75t_R FILLER_263_370 ();
 DECAPx6_ASAP7_75t_R FILLER_263_392 ();
 DECAPx2_ASAP7_75t_R FILLER_263_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_412 ();
 DECAPx10_ASAP7_75t_R FILLER_263_419 ();
 DECAPx1_ASAP7_75t_R FILLER_263_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_445 ();
 DECAPx10_ASAP7_75t_R FILLER_263_456 ();
 DECAPx10_ASAP7_75t_R FILLER_263_478 ();
 DECAPx10_ASAP7_75t_R FILLER_263_500 ();
 DECAPx10_ASAP7_75t_R FILLER_263_522 ();
 DECAPx10_ASAP7_75t_R FILLER_263_544 ();
 DECAPx10_ASAP7_75t_R FILLER_263_566 ();
 DECAPx10_ASAP7_75t_R FILLER_263_588 ();
 DECAPx10_ASAP7_75t_R FILLER_263_610 ();
 DECAPx10_ASAP7_75t_R FILLER_263_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_654 ();
 DECAPx4_ASAP7_75t_R FILLER_263_669 ();
 DECAPx10_ASAP7_75t_R FILLER_263_687 ();
 DECAPx4_ASAP7_75t_R FILLER_263_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_727 ();
 DECAPx4_ASAP7_75t_R FILLER_263_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_744 ();
 DECAPx10_ASAP7_75t_R FILLER_263_751 ();
 DECAPx1_ASAP7_75t_R FILLER_263_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_777 ();
 DECAPx10_ASAP7_75t_R FILLER_263_792 ();
 DECAPx10_ASAP7_75t_R FILLER_263_814 ();
 DECAPx6_ASAP7_75t_R FILLER_263_836 ();
 FILLER_ASAP7_75t_R FILLER_263_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_852 ();
 DECAPx6_ASAP7_75t_R FILLER_263_870 ();
 DECAPx1_ASAP7_75t_R FILLER_263_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_888 ();
 DECAPx2_ASAP7_75t_R FILLER_263_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_943 ();
 DECAPx6_ASAP7_75t_R FILLER_263_986 ();
 FILLER_ASAP7_75t_R FILLER_263_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_263_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_263_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_263_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_263_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_263_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_264_172 ();
 DECAPx10_ASAP7_75t_R FILLER_264_194 ();
 DECAPx10_ASAP7_75t_R FILLER_264_216 ();
 DECAPx10_ASAP7_75t_R FILLER_264_238 ();
 DECAPx10_ASAP7_75t_R FILLER_264_260 ();
 DECAPx10_ASAP7_75t_R FILLER_264_282 ();
 DECAPx10_ASAP7_75t_R FILLER_264_304 ();
 DECAPx10_ASAP7_75t_R FILLER_264_326 ();
 DECAPx10_ASAP7_75t_R FILLER_264_348 ();
 DECAPx10_ASAP7_75t_R FILLER_264_370 ();
 DECAPx10_ASAP7_75t_R FILLER_264_392 ();
 DECAPx10_ASAP7_75t_R FILLER_264_414 ();
 DECAPx10_ASAP7_75t_R FILLER_264_436 ();
 DECAPx10_ASAP7_75t_R FILLER_264_458 ();
 DECAPx10_ASAP7_75t_R FILLER_264_480 ();
 DECAPx10_ASAP7_75t_R FILLER_264_502 ();
 DECAPx10_ASAP7_75t_R FILLER_264_524 ();
 DECAPx10_ASAP7_75t_R FILLER_264_546 ();
 DECAPx10_ASAP7_75t_R FILLER_264_568 ();
 DECAPx10_ASAP7_75t_R FILLER_264_590 ();
 DECAPx6_ASAP7_75t_R FILLER_264_612 ();
 DECAPx2_ASAP7_75t_R FILLER_264_626 ();
 DECAPx1_ASAP7_75t_R FILLER_264_634 ();
 DECAPx10_ASAP7_75t_R FILLER_264_667 ();
 FILLER_ASAP7_75t_R FILLER_264_689 ();
 DECAPx6_ASAP7_75t_R FILLER_264_699 ();
 FILLER_ASAP7_75t_R FILLER_264_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_715 ();
 DECAPx4_ASAP7_75t_R FILLER_264_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_738 ();
 DECAPx2_ASAP7_75t_R FILLER_264_742 ();
 DECAPx1_ASAP7_75t_R FILLER_264_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_763 ();
 DECAPx2_ASAP7_75t_R FILLER_264_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_794 ();
 DECAPx6_ASAP7_75t_R FILLER_264_801 ();
 DECAPx1_ASAP7_75t_R FILLER_264_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_819 ();
 DECAPx1_ASAP7_75t_R FILLER_264_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_849 ();
 FILLER_ASAP7_75t_R FILLER_264_853 ();
 DECAPx10_ASAP7_75t_R FILLER_264_897 ();
 DECAPx6_ASAP7_75t_R FILLER_264_919 ();
 DECAPx1_ASAP7_75t_R FILLER_264_933 ();
 DECAPx6_ASAP7_75t_R FILLER_264_981 ();
 FILLER_ASAP7_75t_R FILLER_264_995 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_264_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_265_172 ();
 DECAPx10_ASAP7_75t_R FILLER_265_194 ();
 DECAPx10_ASAP7_75t_R FILLER_265_216 ();
 DECAPx10_ASAP7_75t_R FILLER_265_238 ();
 DECAPx10_ASAP7_75t_R FILLER_265_260 ();
 DECAPx10_ASAP7_75t_R FILLER_265_282 ();
 DECAPx10_ASAP7_75t_R FILLER_265_304 ();
 DECAPx10_ASAP7_75t_R FILLER_265_326 ();
 DECAPx10_ASAP7_75t_R FILLER_265_348 ();
 DECAPx10_ASAP7_75t_R FILLER_265_370 ();
 DECAPx10_ASAP7_75t_R FILLER_265_392 ();
 DECAPx10_ASAP7_75t_R FILLER_265_414 ();
 DECAPx10_ASAP7_75t_R FILLER_265_436 ();
 DECAPx10_ASAP7_75t_R FILLER_265_458 ();
 DECAPx10_ASAP7_75t_R FILLER_265_480 ();
 DECAPx10_ASAP7_75t_R FILLER_265_502 ();
 DECAPx10_ASAP7_75t_R FILLER_265_524 ();
 DECAPx10_ASAP7_75t_R FILLER_265_546 ();
 DECAPx10_ASAP7_75t_R FILLER_265_568 ();
 DECAPx10_ASAP7_75t_R FILLER_265_590 ();
 DECAPx10_ASAP7_75t_R FILLER_265_612 ();
 DECAPx10_ASAP7_75t_R FILLER_265_634 ();
 DECAPx1_ASAP7_75t_R FILLER_265_656 ();
 DECAPx4_ASAP7_75t_R FILLER_265_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_673 ();
 FILLER_ASAP7_75t_R FILLER_265_677 ();
 DECAPx2_ASAP7_75t_R FILLER_265_763 ();
 FILLER_ASAP7_75t_R FILLER_265_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_771 ();
 DECAPx4_ASAP7_75t_R FILLER_265_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_790 ();
 DECAPx4_ASAP7_75t_R FILLER_265_812 ();
 DECAPx10_ASAP7_75t_R FILLER_265_864 ();
 DECAPx6_ASAP7_75t_R FILLER_265_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_900 ();
 DECAPx10_ASAP7_75t_R FILLER_265_907 ();
 DECAPx6_ASAP7_75t_R FILLER_265_929 ();
 DECAPx1_ASAP7_75t_R FILLER_265_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_947 ();
 DECAPx10_ASAP7_75t_R FILLER_265_954 ();
 DECAPx10_ASAP7_75t_R FILLER_265_976 ();
 DECAPx10_ASAP7_75t_R FILLER_265_998 ();
 DECAPx6_ASAP7_75t_R FILLER_265_1020 ();
 FILLER_ASAP7_75t_R FILLER_265_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_265_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_265_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_265_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_265_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_266_172 ();
 DECAPx10_ASAP7_75t_R FILLER_266_194 ();
 DECAPx10_ASAP7_75t_R FILLER_266_216 ();
 DECAPx10_ASAP7_75t_R FILLER_266_238 ();
 DECAPx10_ASAP7_75t_R FILLER_266_260 ();
 DECAPx10_ASAP7_75t_R FILLER_266_282 ();
 DECAPx10_ASAP7_75t_R FILLER_266_304 ();
 DECAPx10_ASAP7_75t_R FILLER_266_326 ();
 DECAPx10_ASAP7_75t_R FILLER_266_348 ();
 DECAPx10_ASAP7_75t_R FILLER_266_370 ();
 DECAPx10_ASAP7_75t_R FILLER_266_392 ();
 DECAPx10_ASAP7_75t_R FILLER_266_414 ();
 DECAPx10_ASAP7_75t_R FILLER_266_436 ();
 DECAPx10_ASAP7_75t_R FILLER_266_458 ();
 DECAPx10_ASAP7_75t_R FILLER_266_480 ();
 DECAPx10_ASAP7_75t_R FILLER_266_502 ();
 DECAPx10_ASAP7_75t_R FILLER_266_524 ();
 DECAPx10_ASAP7_75t_R FILLER_266_546 ();
 DECAPx10_ASAP7_75t_R FILLER_266_568 ();
 DECAPx10_ASAP7_75t_R FILLER_266_590 ();
 DECAPx6_ASAP7_75t_R FILLER_266_612 ();
 DECAPx2_ASAP7_75t_R FILLER_266_626 ();
 DECAPx10_ASAP7_75t_R FILLER_266_634 ();
 DECAPx4_ASAP7_75t_R FILLER_266_656 ();
 FILLER_ASAP7_75t_R FILLER_266_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_677 ();
 DECAPx2_ASAP7_75t_R FILLER_266_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_690 ();
 DECAPx10_ASAP7_75t_R FILLER_266_700 ();
 DECAPx10_ASAP7_75t_R FILLER_266_722 ();
 DECAPx10_ASAP7_75t_R FILLER_266_744 ();
 DECAPx1_ASAP7_75t_R FILLER_266_766 ();
 DECAPx6_ASAP7_75t_R FILLER_266_776 ();
 DECAPx2_ASAP7_75t_R FILLER_266_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_796 ();
 DECAPx6_ASAP7_75t_R FILLER_266_808 ();
 DECAPx10_ASAP7_75t_R FILLER_266_828 ();
 DECAPx10_ASAP7_75t_R FILLER_266_850 ();
 DECAPx10_ASAP7_75t_R FILLER_266_872 ();
 DECAPx2_ASAP7_75t_R FILLER_266_894 ();
 FILLER_ASAP7_75t_R FILLER_266_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_908 ();
 DECAPx10_ASAP7_75t_R FILLER_266_929 ();
 DECAPx10_ASAP7_75t_R FILLER_266_951 ();
 FILLER_ASAP7_75t_R FILLER_266_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_975 ();
 DECAPx10_ASAP7_75t_R FILLER_266_979 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_266_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_267_172 ();
 DECAPx10_ASAP7_75t_R FILLER_267_194 ();
 DECAPx10_ASAP7_75t_R FILLER_267_216 ();
 DECAPx10_ASAP7_75t_R FILLER_267_238 ();
 DECAPx10_ASAP7_75t_R FILLER_267_260 ();
 DECAPx10_ASAP7_75t_R FILLER_267_282 ();
 DECAPx10_ASAP7_75t_R FILLER_267_304 ();
 DECAPx10_ASAP7_75t_R FILLER_267_326 ();
 DECAPx10_ASAP7_75t_R FILLER_267_348 ();
 DECAPx10_ASAP7_75t_R FILLER_267_370 ();
 DECAPx10_ASAP7_75t_R FILLER_267_392 ();
 DECAPx10_ASAP7_75t_R FILLER_267_414 ();
 DECAPx10_ASAP7_75t_R FILLER_267_436 ();
 DECAPx10_ASAP7_75t_R FILLER_267_458 ();
 DECAPx10_ASAP7_75t_R FILLER_267_480 ();
 DECAPx10_ASAP7_75t_R FILLER_267_502 ();
 DECAPx10_ASAP7_75t_R FILLER_267_524 ();
 DECAPx10_ASAP7_75t_R FILLER_267_546 ();
 DECAPx10_ASAP7_75t_R FILLER_267_568 ();
 DECAPx10_ASAP7_75t_R FILLER_267_590 ();
 DECAPx10_ASAP7_75t_R FILLER_267_612 ();
 FILLER_ASAP7_75t_R FILLER_267_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_636 ();
 DECAPx10_ASAP7_75t_R FILLER_267_679 ();
 DECAPx4_ASAP7_75t_R FILLER_267_701 ();
 FILLER_ASAP7_75t_R FILLER_267_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_713 ();
 DECAPx10_ASAP7_75t_R FILLER_267_717 ();
 DECAPx6_ASAP7_75t_R FILLER_267_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_753 ();
 DECAPx10_ASAP7_75t_R FILLER_267_757 ();
 DECAPx10_ASAP7_75t_R FILLER_267_779 ();
 DECAPx10_ASAP7_75t_R FILLER_267_801 ();
 DECAPx6_ASAP7_75t_R FILLER_267_823 ();
 DECAPx4_ASAP7_75t_R FILLER_267_840 ();
 FILLER_ASAP7_75t_R FILLER_267_850 ();
 DECAPx10_ASAP7_75t_R FILLER_267_860 ();
 FILLER_ASAP7_75t_R FILLER_267_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_913 ();
 DECAPx1_ASAP7_75t_R FILLER_267_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_939 ();
 DECAPx2_ASAP7_75t_R FILLER_267_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_978 ();
 FILLER_ASAP7_75t_R FILLER_267_985 ();
 FILLER_ASAP7_75t_R FILLER_267_995 ();
 FILLER_ASAP7_75t_R FILLER_267_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_267_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1030 ();
 FILLER_ASAP7_75t_R FILLER_267_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_267_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_267_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_267_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_268_172 ();
 DECAPx10_ASAP7_75t_R FILLER_268_194 ();
 DECAPx10_ASAP7_75t_R FILLER_268_216 ();
 DECAPx10_ASAP7_75t_R FILLER_268_238 ();
 DECAPx10_ASAP7_75t_R FILLER_268_260 ();
 DECAPx10_ASAP7_75t_R FILLER_268_282 ();
 DECAPx10_ASAP7_75t_R FILLER_268_304 ();
 DECAPx10_ASAP7_75t_R FILLER_268_326 ();
 DECAPx10_ASAP7_75t_R FILLER_268_348 ();
 DECAPx10_ASAP7_75t_R FILLER_268_370 ();
 DECAPx10_ASAP7_75t_R FILLER_268_392 ();
 DECAPx10_ASAP7_75t_R FILLER_268_414 ();
 DECAPx10_ASAP7_75t_R FILLER_268_436 ();
 DECAPx10_ASAP7_75t_R FILLER_268_458 ();
 DECAPx10_ASAP7_75t_R FILLER_268_480 ();
 DECAPx10_ASAP7_75t_R FILLER_268_502 ();
 DECAPx10_ASAP7_75t_R FILLER_268_524 ();
 DECAPx10_ASAP7_75t_R FILLER_268_546 ();
 DECAPx10_ASAP7_75t_R FILLER_268_568 ();
 DECAPx10_ASAP7_75t_R FILLER_268_590 ();
 DECAPx6_ASAP7_75t_R FILLER_268_612 ();
 DECAPx2_ASAP7_75t_R FILLER_268_626 ();
 DECAPx1_ASAP7_75t_R FILLER_268_634 ();
 DECAPx10_ASAP7_75t_R FILLER_268_649 ();
 DECAPx6_ASAP7_75t_R FILLER_268_671 ();
 DECAPx2_ASAP7_75t_R FILLER_268_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_691 ();
 DECAPx4_ASAP7_75t_R FILLER_268_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_710 ();
 DECAPx4_ASAP7_75t_R FILLER_268_719 ();
 FILLER_ASAP7_75t_R FILLER_268_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_731 ();
 DECAPx2_ASAP7_75t_R FILLER_268_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_749 ();
 DECAPx6_ASAP7_75t_R FILLER_268_758 ();
 DECAPx4_ASAP7_75t_R FILLER_268_783 ();
 FILLER_ASAP7_75t_R FILLER_268_793 ();
 DECAPx4_ASAP7_75t_R FILLER_268_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_808 ();
 DECAPx4_ASAP7_75t_R FILLER_268_820 ();
 FILLER_ASAP7_75t_R FILLER_268_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_832 ();
 DECAPx10_ASAP7_75t_R FILLER_268_841 ();
 DECAPx10_ASAP7_75t_R FILLER_268_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_885 ();
 DECAPx2_ASAP7_75t_R FILLER_268_894 ();
 FILLER_ASAP7_75t_R FILLER_268_900 ();
 DECAPx1_ASAP7_75t_R FILLER_268_919 ();
 DECAPx1_ASAP7_75t_R FILLER_268_929 ();
 DECAPx4_ASAP7_75t_R FILLER_268_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_954 ();
 DECAPx1_ASAP7_75t_R FILLER_268_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_967 ();
 DECAPx2_ASAP7_75t_R FILLER_268_974 ();
 FILLER_ASAP7_75t_R FILLER_268_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_982 ();
 FILLER_ASAP7_75t_R FILLER_268_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_268_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_268_1280 ();
 FILLER_ASAP7_75t_R FILLER_268_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_269_172 ();
 DECAPx10_ASAP7_75t_R FILLER_269_194 ();
 DECAPx10_ASAP7_75t_R FILLER_269_216 ();
 DECAPx10_ASAP7_75t_R FILLER_269_238 ();
 DECAPx10_ASAP7_75t_R FILLER_269_260 ();
 DECAPx10_ASAP7_75t_R FILLER_269_282 ();
 DECAPx10_ASAP7_75t_R FILLER_269_304 ();
 DECAPx10_ASAP7_75t_R FILLER_269_326 ();
 DECAPx10_ASAP7_75t_R FILLER_269_348 ();
 DECAPx10_ASAP7_75t_R FILLER_269_370 ();
 DECAPx10_ASAP7_75t_R FILLER_269_392 ();
 DECAPx10_ASAP7_75t_R FILLER_269_414 ();
 DECAPx10_ASAP7_75t_R FILLER_269_436 ();
 DECAPx10_ASAP7_75t_R FILLER_269_458 ();
 DECAPx10_ASAP7_75t_R FILLER_269_480 ();
 DECAPx10_ASAP7_75t_R FILLER_269_502 ();
 DECAPx10_ASAP7_75t_R FILLER_269_524 ();
 DECAPx10_ASAP7_75t_R FILLER_269_546 ();
 DECAPx10_ASAP7_75t_R FILLER_269_568 ();
 DECAPx10_ASAP7_75t_R FILLER_269_590 ();
 DECAPx10_ASAP7_75t_R FILLER_269_612 ();
 DECAPx1_ASAP7_75t_R FILLER_269_634 ();
 DECAPx6_ASAP7_75t_R FILLER_269_644 ();
 FILLER_ASAP7_75t_R FILLER_269_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_660 ();
 DECAPx2_ASAP7_75t_R FILLER_269_814 ();
 FILLER_ASAP7_75t_R FILLER_269_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_822 ();
 DECAPx10_ASAP7_75t_R FILLER_269_850 ();
 DECAPx10_ASAP7_75t_R FILLER_269_872 ();
 DECAPx6_ASAP7_75t_R FILLER_269_894 ();
 DECAPx1_ASAP7_75t_R FILLER_269_916 ();
 FILLER_ASAP7_75t_R FILLER_269_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_928 ();
 DECAPx4_ASAP7_75t_R FILLER_269_956 ();
 DECAPx10_ASAP7_75t_R FILLER_269_987 ();
 DECAPx6_ASAP7_75t_R FILLER_269_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_269_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1069 ();
 FILLER_ASAP7_75t_R FILLER_269_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_269_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_269_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_270_172 ();
 DECAPx10_ASAP7_75t_R FILLER_270_194 ();
 DECAPx10_ASAP7_75t_R FILLER_270_216 ();
 DECAPx10_ASAP7_75t_R FILLER_270_238 ();
 DECAPx10_ASAP7_75t_R FILLER_270_260 ();
 DECAPx10_ASAP7_75t_R FILLER_270_282 ();
 DECAPx10_ASAP7_75t_R FILLER_270_304 ();
 DECAPx10_ASAP7_75t_R FILLER_270_326 ();
 DECAPx10_ASAP7_75t_R FILLER_270_348 ();
 DECAPx10_ASAP7_75t_R FILLER_270_370 ();
 DECAPx10_ASAP7_75t_R FILLER_270_392 ();
 DECAPx10_ASAP7_75t_R FILLER_270_414 ();
 DECAPx10_ASAP7_75t_R FILLER_270_436 ();
 DECAPx10_ASAP7_75t_R FILLER_270_458 ();
 DECAPx10_ASAP7_75t_R FILLER_270_480 ();
 DECAPx10_ASAP7_75t_R FILLER_270_502 ();
 DECAPx10_ASAP7_75t_R FILLER_270_524 ();
 DECAPx10_ASAP7_75t_R FILLER_270_546 ();
 DECAPx10_ASAP7_75t_R FILLER_270_568 ();
 DECAPx10_ASAP7_75t_R FILLER_270_590 ();
 DECAPx6_ASAP7_75t_R FILLER_270_612 ();
 DECAPx2_ASAP7_75t_R FILLER_270_626 ();
 DECAPx10_ASAP7_75t_R FILLER_270_634 ();
 DECAPx6_ASAP7_75t_R FILLER_270_656 ();
 FILLER_ASAP7_75t_R FILLER_270_670 ();
 DECAPx4_ASAP7_75t_R FILLER_270_675 ();
 FILLER_ASAP7_75t_R FILLER_270_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_687 ();
 FILLER_ASAP7_75t_R FILLER_270_694 ();
 DECAPx4_ASAP7_75t_R FILLER_270_699 ();
 FILLER_ASAP7_75t_R FILLER_270_709 ();
 DECAPx4_ASAP7_75t_R FILLER_270_717 ();
 FILLER_ASAP7_75t_R FILLER_270_727 ();
 DECAPx6_ASAP7_75t_R FILLER_270_735 ();
 DECAPx6_ASAP7_75t_R FILLER_270_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_769 ();
 DECAPx6_ASAP7_75t_R FILLER_270_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_790 ();
 FILLER_ASAP7_75t_R FILLER_270_799 ();
 DECAPx2_ASAP7_75t_R FILLER_270_822 ();
 FILLER_ASAP7_75t_R FILLER_270_828 ();
 DECAPx10_ASAP7_75t_R FILLER_270_836 ();
 DECAPx10_ASAP7_75t_R FILLER_270_858 ();
 DECAPx10_ASAP7_75t_R FILLER_270_880 ();
 DECAPx2_ASAP7_75t_R FILLER_270_902 ();
 FILLER_ASAP7_75t_R FILLER_270_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_910 ();
 DECAPx6_ASAP7_75t_R FILLER_270_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_933 ();
 DECAPx6_ASAP7_75t_R FILLER_270_937 ();
 DECAPx1_ASAP7_75t_R FILLER_270_951 ();
 DECAPx10_ASAP7_75t_R FILLER_270_958 ();
 DECAPx10_ASAP7_75t_R FILLER_270_980 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_270_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_271_172 ();
 DECAPx10_ASAP7_75t_R FILLER_271_194 ();
 DECAPx10_ASAP7_75t_R FILLER_271_216 ();
 DECAPx10_ASAP7_75t_R FILLER_271_238 ();
 DECAPx10_ASAP7_75t_R FILLER_271_260 ();
 DECAPx10_ASAP7_75t_R FILLER_271_282 ();
 DECAPx10_ASAP7_75t_R FILLER_271_304 ();
 DECAPx10_ASAP7_75t_R FILLER_271_326 ();
 DECAPx10_ASAP7_75t_R FILLER_271_348 ();
 DECAPx10_ASAP7_75t_R FILLER_271_370 ();
 DECAPx10_ASAP7_75t_R FILLER_271_392 ();
 DECAPx10_ASAP7_75t_R FILLER_271_414 ();
 DECAPx10_ASAP7_75t_R FILLER_271_436 ();
 DECAPx10_ASAP7_75t_R FILLER_271_458 ();
 DECAPx10_ASAP7_75t_R FILLER_271_480 ();
 DECAPx6_ASAP7_75t_R FILLER_271_502 ();
 DECAPx2_ASAP7_75t_R FILLER_271_516 ();
 DECAPx10_ASAP7_75t_R FILLER_271_532 ();
 DECAPx10_ASAP7_75t_R FILLER_271_554 ();
 DECAPx10_ASAP7_75t_R FILLER_271_576 ();
 DECAPx10_ASAP7_75t_R FILLER_271_598 ();
 DECAPx10_ASAP7_75t_R FILLER_271_620 ();
 DECAPx10_ASAP7_75t_R FILLER_271_642 ();
 DECAPx6_ASAP7_75t_R FILLER_271_664 ();
 FILLER_ASAP7_75t_R FILLER_271_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_680 ();
 DECAPx10_ASAP7_75t_R FILLER_271_684 ();
 DECAPx1_ASAP7_75t_R FILLER_271_706 ();
 DECAPx2_ASAP7_75t_R FILLER_271_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_722 ();
 DECAPx4_ASAP7_75t_R FILLER_271_729 ();
 FILLER_ASAP7_75t_R FILLER_271_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_741 ();
 DECAPx6_ASAP7_75t_R FILLER_271_778 ();
 DECAPx10_ASAP7_75t_R FILLER_271_798 ();
 DECAPx10_ASAP7_75t_R FILLER_271_820 ();
 DECAPx10_ASAP7_75t_R FILLER_271_842 ();
 DECAPx10_ASAP7_75t_R FILLER_271_864 ();
 DECAPx4_ASAP7_75t_R FILLER_271_886 ();
 DECAPx4_ASAP7_75t_R FILLER_271_917 ();
 FILLER_ASAP7_75t_R FILLER_271_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_929 ();
 DECAPx2_ASAP7_75t_R FILLER_271_938 ();
 DECAPx4_ASAP7_75t_R FILLER_271_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_968 ();
 FILLER_ASAP7_75t_R FILLER_271_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_985 ();
 DECAPx4_ASAP7_75t_R FILLER_271_997 ();
 FILLER_ASAP7_75t_R FILLER_271_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_271_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1069 ();
 FILLER_ASAP7_75t_R FILLER_271_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_271_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_271_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_272_172 ();
 DECAPx10_ASAP7_75t_R FILLER_272_194 ();
 DECAPx10_ASAP7_75t_R FILLER_272_216 ();
 DECAPx10_ASAP7_75t_R FILLER_272_238 ();
 DECAPx10_ASAP7_75t_R FILLER_272_260 ();
 DECAPx10_ASAP7_75t_R FILLER_272_282 ();
 DECAPx10_ASAP7_75t_R FILLER_272_304 ();
 DECAPx10_ASAP7_75t_R FILLER_272_326 ();
 DECAPx10_ASAP7_75t_R FILLER_272_348 ();
 DECAPx10_ASAP7_75t_R FILLER_272_370 ();
 DECAPx10_ASAP7_75t_R FILLER_272_392 ();
 DECAPx10_ASAP7_75t_R FILLER_272_414 ();
 DECAPx10_ASAP7_75t_R FILLER_272_436 ();
 DECAPx10_ASAP7_75t_R FILLER_272_458 ();
 DECAPx10_ASAP7_75t_R FILLER_272_480 ();
 DECAPx10_ASAP7_75t_R FILLER_272_502 ();
 DECAPx10_ASAP7_75t_R FILLER_272_524 ();
 DECAPx10_ASAP7_75t_R FILLER_272_546 ();
 DECAPx10_ASAP7_75t_R FILLER_272_568 ();
 DECAPx10_ASAP7_75t_R FILLER_272_590 ();
 DECAPx6_ASAP7_75t_R FILLER_272_612 ();
 DECAPx2_ASAP7_75t_R FILLER_272_626 ();
 DECAPx10_ASAP7_75t_R FILLER_272_634 ();
 DECAPx6_ASAP7_75t_R FILLER_272_656 ();
 DECAPx2_ASAP7_75t_R FILLER_272_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_676 ();
 FILLER_ASAP7_75t_R FILLER_272_691 ();
 DECAPx2_ASAP7_75t_R FILLER_272_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_708 ();
 DECAPx2_ASAP7_75t_R FILLER_272_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_726 ();
 DECAPx4_ASAP7_75t_R FILLER_272_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_753 ();
 DECAPx1_ASAP7_75t_R FILLER_272_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_769 ();
 FILLER_ASAP7_75t_R FILLER_272_776 ();
 DECAPx4_ASAP7_75t_R FILLER_272_784 ();
 FILLER_ASAP7_75t_R FILLER_272_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_796 ();
 DECAPx4_ASAP7_75t_R FILLER_272_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_822 ();
 DECAPx2_ASAP7_75t_R FILLER_272_840 ();
 FILLER_ASAP7_75t_R FILLER_272_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_848 ();
 DECAPx10_ASAP7_75t_R FILLER_272_859 ();
 DECAPx10_ASAP7_75t_R FILLER_272_881 ();
 DECAPx6_ASAP7_75t_R FILLER_272_903 ();
 DECAPx1_ASAP7_75t_R FILLER_272_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_921 ();
 DECAPx1_ASAP7_75t_R FILLER_272_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_974 ();
 DECAPx2_ASAP7_75t_R FILLER_272_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_272_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_272_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_272_1281 ();
 FILLER_ASAP7_75t_R FILLER_272_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_273_172 ();
 DECAPx10_ASAP7_75t_R FILLER_273_194 ();
 DECAPx10_ASAP7_75t_R FILLER_273_216 ();
 DECAPx10_ASAP7_75t_R FILLER_273_238 ();
 DECAPx10_ASAP7_75t_R FILLER_273_260 ();
 DECAPx10_ASAP7_75t_R FILLER_273_282 ();
 DECAPx10_ASAP7_75t_R FILLER_273_304 ();
 DECAPx10_ASAP7_75t_R FILLER_273_326 ();
 DECAPx10_ASAP7_75t_R FILLER_273_348 ();
 DECAPx10_ASAP7_75t_R FILLER_273_370 ();
 DECAPx10_ASAP7_75t_R FILLER_273_392 ();
 DECAPx10_ASAP7_75t_R FILLER_273_414 ();
 DECAPx10_ASAP7_75t_R FILLER_273_436 ();
 DECAPx10_ASAP7_75t_R FILLER_273_458 ();
 DECAPx10_ASAP7_75t_R FILLER_273_480 ();
 DECAPx10_ASAP7_75t_R FILLER_273_502 ();
 DECAPx10_ASAP7_75t_R FILLER_273_524 ();
 DECAPx10_ASAP7_75t_R FILLER_273_546 ();
 DECAPx10_ASAP7_75t_R FILLER_273_568 ();
 DECAPx10_ASAP7_75t_R FILLER_273_590 ();
 DECAPx10_ASAP7_75t_R FILLER_273_612 ();
 DECAPx10_ASAP7_75t_R FILLER_273_634 ();
 DECAPx4_ASAP7_75t_R FILLER_273_656 ();
 DECAPx2_ASAP7_75t_R FILLER_273_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_693 ();
 DECAPx6_ASAP7_75t_R FILLER_273_702 ();
 DECAPx1_ASAP7_75t_R FILLER_273_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_720 ();
 DECAPx2_ASAP7_75t_R FILLER_273_742 ();
 DECAPx2_ASAP7_75t_R FILLER_273_791 ();
 FILLER_ASAP7_75t_R FILLER_273_797 ();
 DECAPx1_ASAP7_75t_R FILLER_273_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_814 ();
 DECAPx10_ASAP7_75t_R FILLER_273_844 ();
 DECAPx10_ASAP7_75t_R FILLER_273_866 ();
 DECAPx10_ASAP7_75t_R FILLER_273_888 ();
 DECAPx10_ASAP7_75t_R FILLER_273_910 ();
 DECAPx10_ASAP7_75t_R FILLER_273_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_954 ();
 DECAPx10_ASAP7_75t_R FILLER_273_976 ();
 DECAPx2_ASAP7_75t_R FILLER_273_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_273_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_273_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_273_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_273_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_273_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_274_172 ();
 DECAPx10_ASAP7_75t_R FILLER_274_194 ();
 DECAPx10_ASAP7_75t_R FILLER_274_216 ();
 DECAPx10_ASAP7_75t_R FILLER_274_238 ();
 DECAPx10_ASAP7_75t_R FILLER_274_260 ();
 DECAPx10_ASAP7_75t_R FILLER_274_282 ();
 DECAPx10_ASAP7_75t_R FILLER_274_304 ();
 DECAPx10_ASAP7_75t_R FILLER_274_326 ();
 DECAPx10_ASAP7_75t_R FILLER_274_348 ();
 DECAPx10_ASAP7_75t_R FILLER_274_370 ();
 DECAPx10_ASAP7_75t_R FILLER_274_392 ();
 DECAPx10_ASAP7_75t_R FILLER_274_414 ();
 DECAPx10_ASAP7_75t_R FILLER_274_436 ();
 DECAPx10_ASAP7_75t_R FILLER_274_458 ();
 DECAPx10_ASAP7_75t_R FILLER_274_480 ();
 DECAPx10_ASAP7_75t_R FILLER_274_502 ();
 DECAPx10_ASAP7_75t_R FILLER_274_524 ();
 DECAPx10_ASAP7_75t_R FILLER_274_546 ();
 DECAPx10_ASAP7_75t_R FILLER_274_568 ();
 DECAPx10_ASAP7_75t_R FILLER_274_590 ();
 DECAPx6_ASAP7_75t_R FILLER_274_612 ();
 DECAPx2_ASAP7_75t_R FILLER_274_626 ();
 DECAPx10_ASAP7_75t_R FILLER_274_634 ();
 DECAPx10_ASAP7_75t_R FILLER_274_656 ();
 FILLER_ASAP7_75t_R FILLER_274_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_680 ();
 DECAPx4_ASAP7_75t_R FILLER_274_723 ();
 FILLER_ASAP7_75t_R FILLER_274_733 ();
 DECAPx6_ASAP7_75t_R FILLER_274_738 ();
 DECAPx1_ASAP7_75t_R FILLER_274_752 ();
 DECAPx6_ASAP7_75t_R FILLER_274_777 ();
 FILLER_ASAP7_75t_R FILLER_274_791 ();
 DECAPx10_ASAP7_75t_R FILLER_274_835 ();
 DECAPx10_ASAP7_75t_R FILLER_274_857 ();
 DECAPx10_ASAP7_75t_R FILLER_274_879 ();
 DECAPx10_ASAP7_75t_R FILLER_274_901 ();
 DECAPx10_ASAP7_75t_R FILLER_274_923 ();
 DECAPx10_ASAP7_75t_R FILLER_274_945 ();
 DECAPx10_ASAP7_75t_R FILLER_274_967 ();
 DECAPx10_ASAP7_75t_R FILLER_274_989 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_274_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_274_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_275_172 ();
 DECAPx10_ASAP7_75t_R FILLER_275_194 ();
 DECAPx10_ASAP7_75t_R FILLER_275_216 ();
 DECAPx10_ASAP7_75t_R FILLER_275_238 ();
 DECAPx10_ASAP7_75t_R FILLER_275_260 ();
 DECAPx10_ASAP7_75t_R FILLER_275_282 ();
 DECAPx10_ASAP7_75t_R FILLER_275_304 ();
 DECAPx10_ASAP7_75t_R FILLER_275_326 ();
 DECAPx10_ASAP7_75t_R FILLER_275_348 ();
 DECAPx10_ASAP7_75t_R FILLER_275_370 ();
 DECAPx10_ASAP7_75t_R FILLER_275_392 ();
 DECAPx10_ASAP7_75t_R FILLER_275_414 ();
 DECAPx10_ASAP7_75t_R FILLER_275_436 ();
 DECAPx10_ASAP7_75t_R FILLER_275_458 ();
 DECAPx10_ASAP7_75t_R FILLER_275_480 ();
 DECAPx10_ASAP7_75t_R FILLER_275_502 ();
 DECAPx10_ASAP7_75t_R FILLER_275_524 ();
 DECAPx10_ASAP7_75t_R FILLER_275_546 ();
 DECAPx10_ASAP7_75t_R FILLER_275_568 ();
 DECAPx10_ASAP7_75t_R FILLER_275_590 ();
 DECAPx10_ASAP7_75t_R FILLER_275_612 ();
 DECAPx10_ASAP7_75t_R FILLER_275_634 ();
 DECAPx10_ASAP7_75t_R FILLER_275_656 ();
 DECAPx10_ASAP7_75t_R FILLER_275_678 ();
 DECAPx10_ASAP7_75t_R FILLER_275_700 ();
 DECAPx2_ASAP7_75t_R FILLER_275_722 ();
 FILLER_ASAP7_75t_R FILLER_275_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_730 ();
 DECAPx10_ASAP7_75t_R FILLER_275_752 ();
 DECAPx10_ASAP7_75t_R FILLER_275_774 ();
 DECAPx10_ASAP7_75t_R FILLER_275_796 ();
 DECAPx10_ASAP7_75t_R FILLER_275_818 ();
 DECAPx10_ASAP7_75t_R FILLER_275_840 ();
 DECAPx10_ASAP7_75t_R FILLER_275_862 ();
 DECAPx10_ASAP7_75t_R FILLER_275_884 ();
 DECAPx10_ASAP7_75t_R FILLER_275_906 ();
 DECAPx10_ASAP7_75t_R FILLER_275_928 ();
 DECAPx10_ASAP7_75t_R FILLER_275_950 ();
 DECAPx10_ASAP7_75t_R FILLER_275_972 ();
 DECAPx10_ASAP7_75t_R FILLER_275_994 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_275_1082 ();
 FILLER_ASAP7_75t_R FILLER_275_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_275_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_275_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_276_172 ();
 DECAPx10_ASAP7_75t_R FILLER_276_194 ();
 DECAPx10_ASAP7_75t_R FILLER_276_216 ();
 DECAPx10_ASAP7_75t_R FILLER_276_238 ();
 DECAPx10_ASAP7_75t_R FILLER_276_260 ();
 DECAPx10_ASAP7_75t_R FILLER_276_282 ();
 DECAPx10_ASAP7_75t_R FILLER_276_304 ();
 DECAPx10_ASAP7_75t_R FILLER_276_326 ();
 DECAPx10_ASAP7_75t_R FILLER_276_348 ();
 DECAPx10_ASAP7_75t_R FILLER_276_370 ();
 DECAPx10_ASAP7_75t_R FILLER_276_392 ();
 DECAPx10_ASAP7_75t_R FILLER_276_414 ();
 DECAPx10_ASAP7_75t_R FILLER_276_436 ();
 DECAPx10_ASAP7_75t_R FILLER_276_458 ();
 DECAPx10_ASAP7_75t_R FILLER_276_480 ();
 DECAPx10_ASAP7_75t_R FILLER_276_502 ();
 DECAPx10_ASAP7_75t_R FILLER_276_524 ();
 DECAPx10_ASAP7_75t_R FILLER_276_546 ();
 DECAPx10_ASAP7_75t_R FILLER_276_568 ();
 DECAPx10_ASAP7_75t_R FILLER_276_590 ();
 DECAPx6_ASAP7_75t_R FILLER_276_612 ();
 DECAPx2_ASAP7_75t_R FILLER_276_626 ();
 DECAPx10_ASAP7_75t_R FILLER_276_634 ();
 DECAPx10_ASAP7_75t_R FILLER_276_656 ();
 DECAPx10_ASAP7_75t_R FILLER_276_678 ();
 DECAPx10_ASAP7_75t_R FILLER_276_700 ();
 DECAPx10_ASAP7_75t_R FILLER_276_722 ();
 DECAPx10_ASAP7_75t_R FILLER_276_744 ();
 DECAPx2_ASAP7_75t_R FILLER_276_766 ();
 FILLER_ASAP7_75t_R FILLER_276_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_774 ();
 DECAPx10_ASAP7_75t_R FILLER_276_796 ();
 DECAPx10_ASAP7_75t_R FILLER_276_818 ();
 DECAPx10_ASAP7_75t_R FILLER_276_840 ();
 DECAPx10_ASAP7_75t_R FILLER_276_862 ();
 DECAPx10_ASAP7_75t_R FILLER_276_884 ();
 DECAPx10_ASAP7_75t_R FILLER_276_906 ();
 DECAPx10_ASAP7_75t_R FILLER_276_928 ();
 DECAPx10_ASAP7_75t_R FILLER_276_950 ();
 DECAPx10_ASAP7_75t_R FILLER_276_972 ();
 DECAPx10_ASAP7_75t_R FILLER_276_994 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_276_1280 ();
 FILLER_ASAP7_75t_R FILLER_276_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_277_172 ();
 DECAPx10_ASAP7_75t_R FILLER_277_194 ();
 DECAPx10_ASAP7_75t_R FILLER_277_216 ();
 DECAPx10_ASAP7_75t_R FILLER_277_238 ();
 DECAPx10_ASAP7_75t_R FILLER_277_260 ();
 DECAPx10_ASAP7_75t_R FILLER_277_282 ();
 DECAPx10_ASAP7_75t_R FILLER_277_304 ();
 DECAPx10_ASAP7_75t_R FILLER_277_326 ();
 DECAPx10_ASAP7_75t_R FILLER_277_348 ();
 DECAPx10_ASAP7_75t_R FILLER_277_370 ();
 DECAPx10_ASAP7_75t_R FILLER_277_392 ();
 DECAPx10_ASAP7_75t_R FILLER_277_414 ();
 DECAPx10_ASAP7_75t_R FILLER_277_436 ();
 DECAPx10_ASAP7_75t_R FILLER_277_458 ();
 DECAPx10_ASAP7_75t_R FILLER_277_480 ();
 DECAPx10_ASAP7_75t_R FILLER_277_502 ();
 DECAPx10_ASAP7_75t_R FILLER_277_524 ();
 DECAPx10_ASAP7_75t_R FILLER_277_546 ();
 DECAPx10_ASAP7_75t_R FILLER_277_568 ();
 DECAPx10_ASAP7_75t_R FILLER_277_590 ();
 DECAPx10_ASAP7_75t_R FILLER_277_612 ();
 DECAPx10_ASAP7_75t_R FILLER_277_634 ();
 DECAPx10_ASAP7_75t_R FILLER_277_656 ();
 DECAPx10_ASAP7_75t_R FILLER_277_678 ();
 DECAPx10_ASAP7_75t_R FILLER_277_700 ();
 DECAPx10_ASAP7_75t_R FILLER_277_722 ();
 DECAPx10_ASAP7_75t_R FILLER_277_744 ();
 DECAPx10_ASAP7_75t_R FILLER_277_766 ();
 DECAPx10_ASAP7_75t_R FILLER_277_788 ();
 DECAPx10_ASAP7_75t_R FILLER_277_810 ();
 DECAPx10_ASAP7_75t_R FILLER_277_832 ();
 DECAPx10_ASAP7_75t_R FILLER_277_854 ();
 DECAPx10_ASAP7_75t_R FILLER_277_876 ();
 DECAPx10_ASAP7_75t_R FILLER_277_898 ();
 DECAPx10_ASAP7_75t_R FILLER_277_920 ();
 DECAPx10_ASAP7_75t_R FILLER_277_942 ();
 DECAPx10_ASAP7_75t_R FILLER_277_964 ();
 DECAPx10_ASAP7_75t_R FILLER_277_986 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_277_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_277_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_277_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_277_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_278_172 ();
 DECAPx10_ASAP7_75t_R FILLER_278_194 ();
 DECAPx10_ASAP7_75t_R FILLER_278_216 ();
 DECAPx10_ASAP7_75t_R FILLER_278_238 ();
 DECAPx10_ASAP7_75t_R FILLER_278_260 ();
 DECAPx10_ASAP7_75t_R FILLER_278_282 ();
 DECAPx10_ASAP7_75t_R FILLER_278_304 ();
 DECAPx10_ASAP7_75t_R FILLER_278_326 ();
 DECAPx10_ASAP7_75t_R FILLER_278_348 ();
 DECAPx10_ASAP7_75t_R FILLER_278_370 ();
 DECAPx10_ASAP7_75t_R FILLER_278_392 ();
 DECAPx10_ASAP7_75t_R FILLER_278_414 ();
 DECAPx10_ASAP7_75t_R FILLER_278_436 ();
 DECAPx10_ASAP7_75t_R FILLER_278_458 ();
 DECAPx10_ASAP7_75t_R FILLER_278_480 ();
 DECAPx10_ASAP7_75t_R FILLER_278_502 ();
 DECAPx10_ASAP7_75t_R FILLER_278_524 ();
 DECAPx10_ASAP7_75t_R FILLER_278_546 ();
 DECAPx10_ASAP7_75t_R FILLER_278_568 ();
 DECAPx10_ASAP7_75t_R FILLER_278_590 ();
 DECAPx6_ASAP7_75t_R FILLER_278_612 ();
 DECAPx2_ASAP7_75t_R FILLER_278_626 ();
 DECAPx10_ASAP7_75t_R FILLER_278_634 ();
 DECAPx10_ASAP7_75t_R FILLER_278_656 ();
 DECAPx10_ASAP7_75t_R FILLER_278_678 ();
 DECAPx10_ASAP7_75t_R FILLER_278_700 ();
 DECAPx10_ASAP7_75t_R FILLER_278_722 ();
 DECAPx10_ASAP7_75t_R FILLER_278_744 ();
 DECAPx10_ASAP7_75t_R FILLER_278_766 ();
 DECAPx10_ASAP7_75t_R FILLER_278_788 ();
 DECAPx10_ASAP7_75t_R FILLER_278_810 ();
 DECAPx10_ASAP7_75t_R FILLER_278_832 ();
 DECAPx10_ASAP7_75t_R FILLER_278_854 ();
 DECAPx10_ASAP7_75t_R FILLER_278_876 ();
 DECAPx10_ASAP7_75t_R FILLER_278_898 ();
 DECAPx10_ASAP7_75t_R FILLER_278_920 ();
 DECAPx10_ASAP7_75t_R FILLER_278_942 ();
 DECAPx10_ASAP7_75t_R FILLER_278_964 ();
 DECAPx10_ASAP7_75t_R FILLER_278_986 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_278_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_278_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_279_172 ();
 DECAPx10_ASAP7_75t_R FILLER_279_194 ();
 DECAPx10_ASAP7_75t_R FILLER_279_216 ();
 DECAPx10_ASAP7_75t_R FILLER_279_238 ();
 DECAPx10_ASAP7_75t_R FILLER_279_260 ();
 DECAPx10_ASAP7_75t_R FILLER_279_282 ();
 DECAPx10_ASAP7_75t_R FILLER_279_304 ();
 DECAPx10_ASAP7_75t_R FILLER_279_326 ();
 DECAPx10_ASAP7_75t_R FILLER_279_348 ();
 DECAPx10_ASAP7_75t_R FILLER_279_370 ();
 DECAPx10_ASAP7_75t_R FILLER_279_392 ();
 DECAPx10_ASAP7_75t_R FILLER_279_414 ();
 DECAPx10_ASAP7_75t_R FILLER_279_436 ();
 DECAPx10_ASAP7_75t_R FILLER_279_458 ();
 DECAPx10_ASAP7_75t_R FILLER_279_480 ();
 DECAPx10_ASAP7_75t_R FILLER_279_502 ();
 DECAPx10_ASAP7_75t_R FILLER_279_524 ();
 DECAPx10_ASAP7_75t_R FILLER_279_546 ();
 DECAPx10_ASAP7_75t_R FILLER_279_568 ();
 DECAPx10_ASAP7_75t_R FILLER_279_590 ();
 DECAPx10_ASAP7_75t_R FILLER_279_612 ();
 DECAPx10_ASAP7_75t_R FILLER_279_634 ();
 DECAPx10_ASAP7_75t_R FILLER_279_656 ();
 DECAPx10_ASAP7_75t_R FILLER_279_678 ();
 DECAPx10_ASAP7_75t_R FILLER_279_700 ();
 DECAPx10_ASAP7_75t_R FILLER_279_722 ();
 DECAPx10_ASAP7_75t_R FILLER_279_744 ();
 DECAPx10_ASAP7_75t_R FILLER_279_766 ();
 DECAPx10_ASAP7_75t_R FILLER_279_788 ();
 DECAPx10_ASAP7_75t_R FILLER_279_810 ();
 DECAPx10_ASAP7_75t_R FILLER_279_832 ();
 DECAPx10_ASAP7_75t_R FILLER_279_854 ();
 DECAPx10_ASAP7_75t_R FILLER_279_876 ();
 DECAPx10_ASAP7_75t_R FILLER_279_898 ();
 DECAPx10_ASAP7_75t_R FILLER_279_920 ();
 DECAPx10_ASAP7_75t_R FILLER_279_942 ();
 DECAPx10_ASAP7_75t_R FILLER_279_964 ();
 DECAPx10_ASAP7_75t_R FILLER_279_986 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_279_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_279_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_279_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_279_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_280_172 ();
 DECAPx10_ASAP7_75t_R FILLER_280_194 ();
 DECAPx10_ASAP7_75t_R FILLER_280_216 ();
 DECAPx10_ASAP7_75t_R FILLER_280_238 ();
 DECAPx10_ASAP7_75t_R FILLER_280_260 ();
 DECAPx10_ASAP7_75t_R FILLER_280_282 ();
 DECAPx10_ASAP7_75t_R FILLER_280_304 ();
 DECAPx10_ASAP7_75t_R FILLER_280_326 ();
 DECAPx10_ASAP7_75t_R FILLER_280_348 ();
 DECAPx10_ASAP7_75t_R FILLER_280_370 ();
 DECAPx10_ASAP7_75t_R FILLER_280_392 ();
 DECAPx10_ASAP7_75t_R FILLER_280_414 ();
 DECAPx10_ASAP7_75t_R FILLER_280_436 ();
 DECAPx10_ASAP7_75t_R FILLER_280_458 ();
 DECAPx10_ASAP7_75t_R FILLER_280_480 ();
 DECAPx10_ASAP7_75t_R FILLER_280_502 ();
 DECAPx10_ASAP7_75t_R FILLER_280_524 ();
 DECAPx10_ASAP7_75t_R FILLER_280_546 ();
 DECAPx10_ASAP7_75t_R FILLER_280_568 ();
 DECAPx10_ASAP7_75t_R FILLER_280_590 ();
 DECAPx6_ASAP7_75t_R FILLER_280_612 ();
 DECAPx2_ASAP7_75t_R FILLER_280_626 ();
 DECAPx10_ASAP7_75t_R FILLER_280_634 ();
 DECAPx10_ASAP7_75t_R FILLER_280_656 ();
 DECAPx10_ASAP7_75t_R FILLER_280_678 ();
 DECAPx10_ASAP7_75t_R FILLER_280_700 ();
 DECAPx10_ASAP7_75t_R FILLER_280_722 ();
 DECAPx10_ASAP7_75t_R FILLER_280_744 ();
 DECAPx10_ASAP7_75t_R FILLER_280_766 ();
 DECAPx10_ASAP7_75t_R FILLER_280_788 ();
 DECAPx10_ASAP7_75t_R FILLER_280_810 ();
 DECAPx10_ASAP7_75t_R FILLER_280_832 ();
 DECAPx10_ASAP7_75t_R FILLER_280_854 ();
 DECAPx10_ASAP7_75t_R FILLER_280_876 ();
 DECAPx10_ASAP7_75t_R FILLER_280_898 ();
 DECAPx10_ASAP7_75t_R FILLER_280_920 ();
 DECAPx10_ASAP7_75t_R FILLER_280_942 ();
 DECAPx10_ASAP7_75t_R FILLER_280_964 ();
 DECAPx10_ASAP7_75t_R FILLER_280_986 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_280_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_280_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_281_172 ();
 DECAPx10_ASAP7_75t_R FILLER_281_194 ();
 DECAPx10_ASAP7_75t_R FILLER_281_216 ();
 DECAPx10_ASAP7_75t_R FILLER_281_238 ();
 DECAPx10_ASAP7_75t_R FILLER_281_260 ();
 DECAPx10_ASAP7_75t_R FILLER_281_282 ();
 DECAPx10_ASAP7_75t_R FILLER_281_304 ();
 DECAPx10_ASAP7_75t_R FILLER_281_326 ();
 DECAPx10_ASAP7_75t_R FILLER_281_348 ();
 DECAPx10_ASAP7_75t_R FILLER_281_370 ();
 DECAPx10_ASAP7_75t_R FILLER_281_392 ();
 DECAPx10_ASAP7_75t_R FILLER_281_414 ();
 DECAPx10_ASAP7_75t_R FILLER_281_436 ();
 DECAPx10_ASAP7_75t_R FILLER_281_458 ();
 DECAPx10_ASAP7_75t_R FILLER_281_480 ();
 DECAPx10_ASAP7_75t_R FILLER_281_502 ();
 DECAPx10_ASAP7_75t_R FILLER_281_524 ();
 DECAPx10_ASAP7_75t_R FILLER_281_546 ();
 DECAPx10_ASAP7_75t_R FILLER_281_568 ();
 DECAPx10_ASAP7_75t_R FILLER_281_590 ();
 DECAPx10_ASAP7_75t_R FILLER_281_612 ();
 DECAPx10_ASAP7_75t_R FILLER_281_634 ();
 DECAPx10_ASAP7_75t_R FILLER_281_656 ();
 DECAPx10_ASAP7_75t_R FILLER_281_678 ();
 DECAPx10_ASAP7_75t_R FILLER_281_700 ();
 DECAPx10_ASAP7_75t_R FILLER_281_722 ();
 DECAPx10_ASAP7_75t_R FILLER_281_744 ();
 DECAPx10_ASAP7_75t_R FILLER_281_766 ();
 DECAPx10_ASAP7_75t_R FILLER_281_788 ();
 DECAPx10_ASAP7_75t_R FILLER_281_810 ();
 DECAPx10_ASAP7_75t_R FILLER_281_832 ();
 DECAPx10_ASAP7_75t_R FILLER_281_854 ();
 DECAPx10_ASAP7_75t_R FILLER_281_876 ();
 DECAPx10_ASAP7_75t_R FILLER_281_898 ();
 DECAPx10_ASAP7_75t_R FILLER_281_920 ();
 DECAPx10_ASAP7_75t_R FILLER_281_942 ();
 DECAPx10_ASAP7_75t_R FILLER_281_964 ();
 DECAPx10_ASAP7_75t_R FILLER_281_986 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_281_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_281_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_281_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_281_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_282_172 ();
 DECAPx10_ASAP7_75t_R FILLER_282_194 ();
 DECAPx10_ASAP7_75t_R FILLER_282_216 ();
 DECAPx10_ASAP7_75t_R FILLER_282_238 ();
 DECAPx10_ASAP7_75t_R FILLER_282_260 ();
 DECAPx10_ASAP7_75t_R FILLER_282_282 ();
 DECAPx10_ASAP7_75t_R FILLER_282_304 ();
 DECAPx10_ASAP7_75t_R FILLER_282_326 ();
 DECAPx10_ASAP7_75t_R FILLER_282_348 ();
 DECAPx10_ASAP7_75t_R FILLER_282_370 ();
 DECAPx10_ASAP7_75t_R FILLER_282_392 ();
 DECAPx10_ASAP7_75t_R FILLER_282_414 ();
 DECAPx10_ASAP7_75t_R FILLER_282_436 ();
 DECAPx10_ASAP7_75t_R FILLER_282_458 ();
 DECAPx10_ASAP7_75t_R FILLER_282_480 ();
 DECAPx10_ASAP7_75t_R FILLER_282_502 ();
 DECAPx10_ASAP7_75t_R FILLER_282_524 ();
 DECAPx10_ASAP7_75t_R FILLER_282_546 ();
 DECAPx10_ASAP7_75t_R FILLER_282_568 ();
 DECAPx10_ASAP7_75t_R FILLER_282_590 ();
 DECAPx6_ASAP7_75t_R FILLER_282_612 ();
 DECAPx2_ASAP7_75t_R FILLER_282_626 ();
 DECAPx10_ASAP7_75t_R FILLER_282_634 ();
 DECAPx10_ASAP7_75t_R FILLER_282_656 ();
 DECAPx10_ASAP7_75t_R FILLER_282_678 ();
 DECAPx10_ASAP7_75t_R FILLER_282_700 ();
 DECAPx10_ASAP7_75t_R FILLER_282_722 ();
 DECAPx10_ASAP7_75t_R FILLER_282_744 ();
 DECAPx10_ASAP7_75t_R FILLER_282_766 ();
 DECAPx10_ASAP7_75t_R FILLER_282_788 ();
 DECAPx10_ASAP7_75t_R FILLER_282_810 ();
 DECAPx10_ASAP7_75t_R FILLER_282_832 ();
 DECAPx10_ASAP7_75t_R FILLER_282_854 ();
 DECAPx10_ASAP7_75t_R FILLER_282_876 ();
 DECAPx10_ASAP7_75t_R FILLER_282_898 ();
 DECAPx10_ASAP7_75t_R FILLER_282_920 ();
 DECAPx10_ASAP7_75t_R FILLER_282_942 ();
 DECAPx10_ASAP7_75t_R FILLER_282_964 ();
 DECAPx10_ASAP7_75t_R FILLER_282_986 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_282_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_282_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_283_172 ();
 DECAPx10_ASAP7_75t_R FILLER_283_194 ();
 DECAPx10_ASAP7_75t_R FILLER_283_216 ();
 DECAPx10_ASAP7_75t_R FILLER_283_238 ();
 DECAPx10_ASAP7_75t_R FILLER_283_260 ();
 DECAPx10_ASAP7_75t_R FILLER_283_282 ();
 DECAPx10_ASAP7_75t_R FILLER_283_304 ();
 DECAPx10_ASAP7_75t_R FILLER_283_326 ();
 DECAPx10_ASAP7_75t_R FILLER_283_348 ();
 DECAPx10_ASAP7_75t_R FILLER_283_370 ();
 DECAPx10_ASAP7_75t_R FILLER_283_392 ();
 DECAPx10_ASAP7_75t_R FILLER_283_414 ();
 DECAPx10_ASAP7_75t_R FILLER_283_436 ();
 DECAPx10_ASAP7_75t_R FILLER_283_458 ();
 DECAPx10_ASAP7_75t_R FILLER_283_480 ();
 DECAPx10_ASAP7_75t_R FILLER_283_502 ();
 DECAPx10_ASAP7_75t_R FILLER_283_524 ();
 DECAPx10_ASAP7_75t_R FILLER_283_546 ();
 DECAPx10_ASAP7_75t_R FILLER_283_568 ();
 DECAPx10_ASAP7_75t_R FILLER_283_590 ();
 DECAPx10_ASAP7_75t_R FILLER_283_612 ();
 DECAPx10_ASAP7_75t_R FILLER_283_634 ();
 DECAPx10_ASAP7_75t_R FILLER_283_656 ();
 DECAPx10_ASAP7_75t_R FILLER_283_678 ();
 DECAPx10_ASAP7_75t_R FILLER_283_700 ();
 DECAPx10_ASAP7_75t_R FILLER_283_722 ();
 DECAPx10_ASAP7_75t_R FILLER_283_744 ();
 DECAPx10_ASAP7_75t_R FILLER_283_766 ();
 DECAPx10_ASAP7_75t_R FILLER_283_788 ();
 DECAPx10_ASAP7_75t_R FILLER_283_810 ();
 DECAPx10_ASAP7_75t_R FILLER_283_832 ();
 DECAPx10_ASAP7_75t_R FILLER_283_854 ();
 DECAPx10_ASAP7_75t_R FILLER_283_876 ();
 DECAPx10_ASAP7_75t_R FILLER_283_898 ();
 DECAPx10_ASAP7_75t_R FILLER_283_920 ();
 DECAPx10_ASAP7_75t_R FILLER_283_942 ();
 DECAPx10_ASAP7_75t_R FILLER_283_964 ();
 DECAPx10_ASAP7_75t_R FILLER_283_986 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_283_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_283_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_283_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_283_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_284_172 ();
 DECAPx10_ASAP7_75t_R FILLER_284_194 ();
 DECAPx10_ASAP7_75t_R FILLER_284_216 ();
 DECAPx10_ASAP7_75t_R FILLER_284_238 ();
 DECAPx10_ASAP7_75t_R FILLER_284_260 ();
 DECAPx10_ASAP7_75t_R FILLER_284_282 ();
 DECAPx10_ASAP7_75t_R FILLER_284_304 ();
 DECAPx10_ASAP7_75t_R FILLER_284_326 ();
 DECAPx10_ASAP7_75t_R FILLER_284_348 ();
 DECAPx10_ASAP7_75t_R FILLER_284_370 ();
 DECAPx10_ASAP7_75t_R FILLER_284_392 ();
 DECAPx10_ASAP7_75t_R FILLER_284_414 ();
 DECAPx10_ASAP7_75t_R FILLER_284_436 ();
 DECAPx10_ASAP7_75t_R FILLER_284_458 ();
 DECAPx10_ASAP7_75t_R FILLER_284_480 ();
 DECAPx10_ASAP7_75t_R FILLER_284_502 ();
 DECAPx10_ASAP7_75t_R FILLER_284_524 ();
 DECAPx10_ASAP7_75t_R FILLER_284_546 ();
 DECAPx10_ASAP7_75t_R FILLER_284_568 ();
 DECAPx10_ASAP7_75t_R FILLER_284_590 ();
 DECAPx6_ASAP7_75t_R FILLER_284_612 ();
 DECAPx2_ASAP7_75t_R FILLER_284_626 ();
 DECAPx10_ASAP7_75t_R FILLER_284_634 ();
 DECAPx10_ASAP7_75t_R FILLER_284_656 ();
 DECAPx10_ASAP7_75t_R FILLER_284_678 ();
 DECAPx10_ASAP7_75t_R FILLER_284_700 ();
 DECAPx10_ASAP7_75t_R FILLER_284_722 ();
 DECAPx10_ASAP7_75t_R FILLER_284_744 ();
 DECAPx10_ASAP7_75t_R FILLER_284_766 ();
 DECAPx10_ASAP7_75t_R FILLER_284_788 ();
 DECAPx10_ASAP7_75t_R FILLER_284_810 ();
 DECAPx10_ASAP7_75t_R FILLER_284_832 ();
 DECAPx10_ASAP7_75t_R FILLER_284_854 ();
 DECAPx10_ASAP7_75t_R FILLER_284_876 ();
 DECAPx10_ASAP7_75t_R FILLER_284_898 ();
 DECAPx10_ASAP7_75t_R FILLER_284_920 ();
 DECAPx10_ASAP7_75t_R FILLER_284_942 ();
 DECAPx10_ASAP7_75t_R FILLER_284_964 ();
 DECAPx10_ASAP7_75t_R FILLER_284_986 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_284_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_284_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_285_172 ();
 DECAPx10_ASAP7_75t_R FILLER_285_194 ();
 DECAPx10_ASAP7_75t_R FILLER_285_216 ();
 DECAPx10_ASAP7_75t_R FILLER_285_238 ();
 DECAPx10_ASAP7_75t_R FILLER_285_260 ();
 DECAPx10_ASAP7_75t_R FILLER_285_282 ();
 DECAPx10_ASAP7_75t_R FILLER_285_304 ();
 DECAPx10_ASAP7_75t_R FILLER_285_326 ();
 DECAPx10_ASAP7_75t_R FILLER_285_348 ();
 DECAPx10_ASAP7_75t_R FILLER_285_370 ();
 DECAPx10_ASAP7_75t_R FILLER_285_392 ();
 DECAPx10_ASAP7_75t_R FILLER_285_414 ();
 DECAPx10_ASAP7_75t_R FILLER_285_436 ();
 DECAPx10_ASAP7_75t_R FILLER_285_458 ();
 DECAPx10_ASAP7_75t_R FILLER_285_480 ();
 DECAPx10_ASAP7_75t_R FILLER_285_502 ();
 DECAPx10_ASAP7_75t_R FILLER_285_524 ();
 DECAPx10_ASAP7_75t_R FILLER_285_546 ();
 DECAPx10_ASAP7_75t_R FILLER_285_568 ();
 DECAPx10_ASAP7_75t_R FILLER_285_590 ();
 DECAPx10_ASAP7_75t_R FILLER_285_612 ();
 DECAPx10_ASAP7_75t_R FILLER_285_634 ();
 DECAPx10_ASAP7_75t_R FILLER_285_656 ();
 DECAPx10_ASAP7_75t_R FILLER_285_678 ();
 DECAPx10_ASAP7_75t_R FILLER_285_700 ();
 DECAPx10_ASAP7_75t_R FILLER_285_722 ();
 DECAPx10_ASAP7_75t_R FILLER_285_744 ();
 DECAPx10_ASAP7_75t_R FILLER_285_766 ();
 DECAPx10_ASAP7_75t_R FILLER_285_788 ();
 DECAPx10_ASAP7_75t_R FILLER_285_810 ();
 DECAPx10_ASAP7_75t_R FILLER_285_832 ();
 DECAPx10_ASAP7_75t_R FILLER_285_854 ();
 DECAPx10_ASAP7_75t_R FILLER_285_876 ();
 DECAPx10_ASAP7_75t_R FILLER_285_898 ();
 DECAPx10_ASAP7_75t_R FILLER_285_920 ();
 DECAPx10_ASAP7_75t_R FILLER_285_942 ();
 DECAPx10_ASAP7_75t_R FILLER_285_964 ();
 DECAPx10_ASAP7_75t_R FILLER_285_986 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_285_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_285_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_285_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_285_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_286_172 ();
 DECAPx10_ASAP7_75t_R FILLER_286_194 ();
 DECAPx10_ASAP7_75t_R FILLER_286_216 ();
 DECAPx10_ASAP7_75t_R FILLER_286_238 ();
 DECAPx10_ASAP7_75t_R FILLER_286_260 ();
 DECAPx10_ASAP7_75t_R FILLER_286_282 ();
 DECAPx10_ASAP7_75t_R FILLER_286_304 ();
 DECAPx10_ASAP7_75t_R FILLER_286_326 ();
 DECAPx10_ASAP7_75t_R FILLER_286_348 ();
 DECAPx10_ASAP7_75t_R FILLER_286_370 ();
 DECAPx10_ASAP7_75t_R FILLER_286_392 ();
 DECAPx10_ASAP7_75t_R FILLER_286_414 ();
 DECAPx10_ASAP7_75t_R FILLER_286_436 ();
 DECAPx10_ASAP7_75t_R FILLER_286_458 ();
 DECAPx10_ASAP7_75t_R FILLER_286_480 ();
 DECAPx10_ASAP7_75t_R FILLER_286_502 ();
 DECAPx10_ASAP7_75t_R FILLER_286_524 ();
 DECAPx10_ASAP7_75t_R FILLER_286_546 ();
 DECAPx10_ASAP7_75t_R FILLER_286_568 ();
 DECAPx10_ASAP7_75t_R FILLER_286_590 ();
 DECAPx6_ASAP7_75t_R FILLER_286_612 ();
 DECAPx2_ASAP7_75t_R FILLER_286_626 ();
 DECAPx10_ASAP7_75t_R FILLER_286_634 ();
 DECAPx10_ASAP7_75t_R FILLER_286_656 ();
 DECAPx10_ASAP7_75t_R FILLER_286_678 ();
 DECAPx10_ASAP7_75t_R FILLER_286_700 ();
 DECAPx10_ASAP7_75t_R FILLER_286_722 ();
 DECAPx10_ASAP7_75t_R FILLER_286_744 ();
 DECAPx10_ASAP7_75t_R FILLER_286_766 ();
 DECAPx10_ASAP7_75t_R FILLER_286_788 ();
 DECAPx10_ASAP7_75t_R FILLER_286_810 ();
 DECAPx10_ASAP7_75t_R FILLER_286_832 ();
 DECAPx10_ASAP7_75t_R FILLER_286_854 ();
 DECAPx10_ASAP7_75t_R FILLER_286_876 ();
 DECAPx10_ASAP7_75t_R FILLER_286_898 ();
 DECAPx10_ASAP7_75t_R FILLER_286_920 ();
 DECAPx10_ASAP7_75t_R FILLER_286_942 ();
 DECAPx10_ASAP7_75t_R FILLER_286_964 ();
 DECAPx10_ASAP7_75t_R FILLER_286_986 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_286_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_286_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_287_172 ();
 DECAPx10_ASAP7_75t_R FILLER_287_194 ();
 DECAPx10_ASAP7_75t_R FILLER_287_216 ();
 DECAPx10_ASAP7_75t_R FILLER_287_238 ();
 DECAPx10_ASAP7_75t_R FILLER_287_260 ();
 DECAPx10_ASAP7_75t_R FILLER_287_282 ();
 DECAPx10_ASAP7_75t_R FILLER_287_304 ();
 DECAPx10_ASAP7_75t_R FILLER_287_326 ();
 DECAPx10_ASAP7_75t_R FILLER_287_348 ();
 DECAPx10_ASAP7_75t_R FILLER_287_370 ();
 DECAPx10_ASAP7_75t_R FILLER_287_392 ();
 DECAPx10_ASAP7_75t_R FILLER_287_414 ();
 DECAPx10_ASAP7_75t_R FILLER_287_436 ();
 DECAPx10_ASAP7_75t_R FILLER_287_458 ();
 DECAPx10_ASAP7_75t_R FILLER_287_480 ();
 DECAPx10_ASAP7_75t_R FILLER_287_502 ();
 DECAPx10_ASAP7_75t_R FILLER_287_524 ();
 DECAPx10_ASAP7_75t_R FILLER_287_546 ();
 DECAPx10_ASAP7_75t_R FILLER_287_568 ();
 DECAPx10_ASAP7_75t_R FILLER_287_590 ();
 DECAPx10_ASAP7_75t_R FILLER_287_612 ();
 DECAPx10_ASAP7_75t_R FILLER_287_634 ();
 DECAPx10_ASAP7_75t_R FILLER_287_656 ();
 DECAPx10_ASAP7_75t_R FILLER_287_678 ();
 DECAPx10_ASAP7_75t_R FILLER_287_700 ();
 DECAPx10_ASAP7_75t_R FILLER_287_722 ();
 DECAPx10_ASAP7_75t_R FILLER_287_744 ();
 DECAPx10_ASAP7_75t_R FILLER_287_766 ();
 DECAPx10_ASAP7_75t_R FILLER_287_788 ();
 DECAPx10_ASAP7_75t_R FILLER_287_810 ();
 DECAPx10_ASAP7_75t_R FILLER_287_832 ();
 DECAPx10_ASAP7_75t_R FILLER_287_854 ();
 DECAPx10_ASAP7_75t_R FILLER_287_876 ();
 DECAPx10_ASAP7_75t_R FILLER_287_898 ();
 DECAPx10_ASAP7_75t_R FILLER_287_920 ();
 DECAPx10_ASAP7_75t_R FILLER_287_942 ();
 DECAPx10_ASAP7_75t_R FILLER_287_964 ();
 DECAPx10_ASAP7_75t_R FILLER_287_986 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_287_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_287_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_287_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_287_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_288_172 ();
 DECAPx10_ASAP7_75t_R FILLER_288_194 ();
 DECAPx10_ASAP7_75t_R FILLER_288_216 ();
 DECAPx10_ASAP7_75t_R FILLER_288_238 ();
 DECAPx10_ASAP7_75t_R FILLER_288_260 ();
 DECAPx10_ASAP7_75t_R FILLER_288_282 ();
 DECAPx10_ASAP7_75t_R FILLER_288_304 ();
 DECAPx10_ASAP7_75t_R FILLER_288_326 ();
 DECAPx10_ASAP7_75t_R FILLER_288_348 ();
 DECAPx10_ASAP7_75t_R FILLER_288_370 ();
 DECAPx10_ASAP7_75t_R FILLER_288_392 ();
 DECAPx10_ASAP7_75t_R FILLER_288_414 ();
 DECAPx10_ASAP7_75t_R FILLER_288_436 ();
 DECAPx10_ASAP7_75t_R FILLER_288_458 ();
 DECAPx10_ASAP7_75t_R FILLER_288_480 ();
 DECAPx10_ASAP7_75t_R FILLER_288_502 ();
 DECAPx10_ASAP7_75t_R FILLER_288_524 ();
 DECAPx10_ASAP7_75t_R FILLER_288_546 ();
 DECAPx10_ASAP7_75t_R FILLER_288_568 ();
 DECAPx10_ASAP7_75t_R FILLER_288_590 ();
 DECAPx6_ASAP7_75t_R FILLER_288_612 ();
 DECAPx2_ASAP7_75t_R FILLER_288_626 ();
 DECAPx10_ASAP7_75t_R FILLER_288_634 ();
 DECAPx10_ASAP7_75t_R FILLER_288_656 ();
 DECAPx10_ASAP7_75t_R FILLER_288_678 ();
 DECAPx10_ASAP7_75t_R FILLER_288_700 ();
 DECAPx10_ASAP7_75t_R FILLER_288_722 ();
 DECAPx10_ASAP7_75t_R FILLER_288_744 ();
 DECAPx10_ASAP7_75t_R FILLER_288_766 ();
 DECAPx10_ASAP7_75t_R FILLER_288_788 ();
 DECAPx10_ASAP7_75t_R FILLER_288_810 ();
 DECAPx10_ASAP7_75t_R FILLER_288_832 ();
 DECAPx10_ASAP7_75t_R FILLER_288_854 ();
 DECAPx10_ASAP7_75t_R FILLER_288_876 ();
 DECAPx10_ASAP7_75t_R FILLER_288_898 ();
 DECAPx10_ASAP7_75t_R FILLER_288_920 ();
 DECAPx10_ASAP7_75t_R FILLER_288_942 ();
 DECAPx10_ASAP7_75t_R FILLER_288_964 ();
 DECAPx10_ASAP7_75t_R FILLER_288_986 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_288_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_288_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_289_172 ();
 DECAPx10_ASAP7_75t_R FILLER_289_194 ();
 DECAPx10_ASAP7_75t_R FILLER_289_216 ();
 DECAPx10_ASAP7_75t_R FILLER_289_238 ();
 DECAPx10_ASAP7_75t_R FILLER_289_260 ();
 DECAPx10_ASAP7_75t_R FILLER_289_282 ();
 DECAPx10_ASAP7_75t_R FILLER_289_304 ();
 DECAPx10_ASAP7_75t_R FILLER_289_326 ();
 DECAPx10_ASAP7_75t_R FILLER_289_348 ();
 DECAPx10_ASAP7_75t_R FILLER_289_370 ();
 DECAPx10_ASAP7_75t_R FILLER_289_392 ();
 DECAPx10_ASAP7_75t_R FILLER_289_414 ();
 DECAPx10_ASAP7_75t_R FILLER_289_436 ();
 DECAPx10_ASAP7_75t_R FILLER_289_458 ();
 DECAPx10_ASAP7_75t_R FILLER_289_480 ();
 DECAPx10_ASAP7_75t_R FILLER_289_502 ();
 DECAPx10_ASAP7_75t_R FILLER_289_524 ();
 DECAPx10_ASAP7_75t_R FILLER_289_546 ();
 DECAPx10_ASAP7_75t_R FILLER_289_568 ();
 DECAPx10_ASAP7_75t_R FILLER_289_590 ();
 DECAPx10_ASAP7_75t_R FILLER_289_612 ();
 DECAPx10_ASAP7_75t_R FILLER_289_634 ();
 DECAPx10_ASAP7_75t_R FILLER_289_656 ();
 DECAPx10_ASAP7_75t_R FILLER_289_678 ();
 DECAPx10_ASAP7_75t_R FILLER_289_700 ();
 DECAPx10_ASAP7_75t_R FILLER_289_722 ();
 DECAPx10_ASAP7_75t_R FILLER_289_744 ();
 DECAPx10_ASAP7_75t_R FILLER_289_766 ();
 DECAPx10_ASAP7_75t_R FILLER_289_788 ();
 DECAPx10_ASAP7_75t_R FILLER_289_810 ();
 DECAPx10_ASAP7_75t_R FILLER_289_832 ();
 DECAPx10_ASAP7_75t_R FILLER_289_854 ();
 DECAPx10_ASAP7_75t_R FILLER_289_876 ();
 DECAPx10_ASAP7_75t_R FILLER_289_898 ();
 DECAPx10_ASAP7_75t_R FILLER_289_920 ();
 DECAPx10_ASAP7_75t_R FILLER_289_942 ();
 DECAPx10_ASAP7_75t_R FILLER_289_964 ();
 DECAPx10_ASAP7_75t_R FILLER_289_986 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_289_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_289_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_289_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_289_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_290_172 ();
 DECAPx10_ASAP7_75t_R FILLER_290_194 ();
 DECAPx10_ASAP7_75t_R FILLER_290_216 ();
 DECAPx10_ASAP7_75t_R FILLER_290_238 ();
 DECAPx10_ASAP7_75t_R FILLER_290_260 ();
 DECAPx10_ASAP7_75t_R FILLER_290_282 ();
 DECAPx10_ASAP7_75t_R FILLER_290_304 ();
 DECAPx10_ASAP7_75t_R FILLER_290_326 ();
 DECAPx10_ASAP7_75t_R FILLER_290_348 ();
 DECAPx10_ASAP7_75t_R FILLER_290_370 ();
 DECAPx10_ASAP7_75t_R FILLER_290_392 ();
 DECAPx10_ASAP7_75t_R FILLER_290_414 ();
 DECAPx10_ASAP7_75t_R FILLER_290_436 ();
 DECAPx10_ASAP7_75t_R FILLER_290_458 ();
 DECAPx10_ASAP7_75t_R FILLER_290_480 ();
 DECAPx10_ASAP7_75t_R FILLER_290_502 ();
 DECAPx10_ASAP7_75t_R FILLER_290_524 ();
 DECAPx10_ASAP7_75t_R FILLER_290_546 ();
 DECAPx10_ASAP7_75t_R FILLER_290_568 ();
 DECAPx10_ASAP7_75t_R FILLER_290_590 ();
 DECAPx6_ASAP7_75t_R FILLER_290_612 ();
 DECAPx2_ASAP7_75t_R FILLER_290_626 ();
 DECAPx10_ASAP7_75t_R FILLER_290_634 ();
 DECAPx10_ASAP7_75t_R FILLER_290_656 ();
 DECAPx10_ASAP7_75t_R FILLER_290_678 ();
 DECAPx10_ASAP7_75t_R FILLER_290_700 ();
 DECAPx10_ASAP7_75t_R FILLER_290_722 ();
 DECAPx10_ASAP7_75t_R FILLER_290_744 ();
 DECAPx10_ASAP7_75t_R FILLER_290_766 ();
 DECAPx10_ASAP7_75t_R FILLER_290_788 ();
 DECAPx10_ASAP7_75t_R FILLER_290_810 ();
 DECAPx10_ASAP7_75t_R FILLER_290_832 ();
 DECAPx10_ASAP7_75t_R FILLER_290_854 ();
 DECAPx10_ASAP7_75t_R FILLER_290_876 ();
 DECAPx10_ASAP7_75t_R FILLER_290_898 ();
 DECAPx10_ASAP7_75t_R FILLER_290_920 ();
 DECAPx10_ASAP7_75t_R FILLER_290_942 ();
 DECAPx10_ASAP7_75t_R FILLER_290_964 ();
 DECAPx10_ASAP7_75t_R FILLER_290_986 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_290_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_290_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_291_172 ();
 DECAPx10_ASAP7_75t_R FILLER_291_194 ();
 DECAPx10_ASAP7_75t_R FILLER_291_216 ();
 DECAPx10_ASAP7_75t_R FILLER_291_238 ();
 DECAPx10_ASAP7_75t_R FILLER_291_260 ();
 DECAPx10_ASAP7_75t_R FILLER_291_282 ();
 DECAPx10_ASAP7_75t_R FILLER_291_304 ();
 DECAPx10_ASAP7_75t_R FILLER_291_326 ();
 DECAPx10_ASAP7_75t_R FILLER_291_348 ();
 DECAPx10_ASAP7_75t_R FILLER_291_370 ();
 DECAPx10_ASAP7_75t_R FILLER_291_392 ();
 DECAPx10_ASAP7_75t_R FILLER_291_414 ();
 DECAPx10_ASAP7_75t_R FILLER_291_436 ();
 DECAPx10_ASAP7_75t_R FILLER_291_458 ();
 DECAPx10_ASAP7_75t_R FILLER_291_480 ();
 DECAPx10_ASAP7_75t_R FILLER_291_502 ();
 DECAPx10_ASAP7_75t_R FILLER_291_524 ();
 DECAPx10_ASAP7_75t_R FILLER_291_546 ();
 DECAPx10_ASAP7_75t_R FILLER_291_568 ();
 DECAPx10_ASAP7_75t_R FILLER_291_590 ();
 DECAPx10_ASAP7_75t_R FILLER_291_612 ();
 DECAPx10_ASAP7_75t_R FILLER_291_634 ();
 DECAPx10_ASAP7_75t_R FILLER_291_656 ();
 DECAPx10_ASAP7_75t_R FILLER_291_678 ();
 DECAPx10_ASAP7_75t_R FILLER_291_700 ();
 DECAPx10_ASAP7_75t_R FILLER_291_722 ();
 DECAPx10_ASAP7_75t_R FILLER_291_744 ();
 DECAPx10_ASAP7_75t_R FILLER_291_766 ();
 DECAPx10_ASAP7_75t_R FILLER_291_788 ();
 DECAPx10_ASAP7_75t_R FILLER_291_810 ();
 DECAPx10_ASAP7_75t_R FILLER_291_832 ();
 DECAPx10_ASAP7_75t_R FILLER_291_854 ();
 DECAPx10_ASAP7_75t_R FILLER_291_876 ();
 DECAPx10_ASAP7_75t_R FILLER_291_898 ();
 DECAPx10_ASAP7_75t_R FILLER_291_920 ();
 DECAPx10_ASAP7_75t_R FILLER_291_942 ();
 DECAPx10_ASAP7_75t_R FILLER_291_964 ();
 DECAPx10_ASAP7_75t_R FILLER_291_986 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_291_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_291_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_291_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_291_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_292_172 ();
 DECAPx10_ASAP7_75t_R FILLER_292_194 ();
 DECAPx10_ASAP7_75t_R FILLER_292_216 ();
 DECAPx10_ASAP7_75t_R FILLER_292_238 ();
 DECAPx10_ASAP7_75t_R FILLER_292_260 ();
 DECAPx10_ASAP7_75t_R FILLER_292_282 ();
 DECAPx10_ASAP7_75t_R FILLER_292_304 ();
 DECAPx10_ASAP7_75t_R FILLER_292_326 ();
 DECAPx10_ASAP7_75t_R FILLER_292_348 ();
 DECAPx10_ASAP7_75t_R FILLER_292_370 ();
 DECAPx10_ASAP7_75t_R FILLER_292_392 ();
 DECAPx10_ASAP7_75t_R FILLER_292_414 ();
 DECAPx10_ASAP7_75t_R FILLER_292_436 ();
 DECAPx10_ASAP7_75t_R FILLER_292_458 ();
 DECAPx10_ASAP7_75t_R FILLER_292_480 ();
 DECAPx10_ASAP7_75t_R FILLER_292_502 ();
 DECAPx10_ASAP7_75t_R FILLER_292_524 ();
 DECAPx10_ASAP7_75t_R FILLER_292_546 ();
 DECAPx10_ASAP7_75t_R FILLER_292_568 ();
 DECAPx10_ASAP7_75t_R FILLER_292_590 ();
 DECAPx6_ASAP7_75t_R FILLER_292_612 ();
 DECAPx2_ASAP7_75t_R FILLER_292_626 ();
 DECAPx10_ASAP7_75t_R FILLER_292_634 ();
 DECAPx10_ASAP7_75t_R FILLER_292_656 ();
 DECAPx10_ASAP7_75t_R FILLER_292_678 ();
 DECAPx10_ASAP7_75t_R FILLER_292_700 ();
 DECAPx10_ASAP7_75t_R FILLER_292_722 ();
 DECAPx10_ASAP7_75t_R FILLER_292_744 ();
 DECAPx10_ASAP7_75t_R FILLER_292_766 ();
 DECAPx10_ASAP7_75t_R FILLER_292_788 ();
 DECAPx10_ASAP7_75t_R FILLER_292_810 ();
 DECAPx10_ASAP7_75t_R FILLER_292_832 ();
 DECAPx10_ASAP7_75t_R FILLER_292_854 ();
 DECAPx10_ASAP7_75t_R FILLER_292_876 ();
 DECAPx10_ASAP7_75t_R FILLER_292_898 ();
 DECAPx10_ASAP7_75t_R FILLER_292_920 ();
 DECAPx10_ASAP7_75t_R FILLER_292_942 ();
 DECAPx10_ASAP7_75t_R FILLER_292_964 ();
 DECAPx10_ASAP7_75t_R FILLER_292_986 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_292_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_292_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_293_172 ();
 DECAPx10_ASAP7_75t_R FILLER_293_194 ();
 DECAPx10_ASAP7_75t_R FILLER_293_216 ();
 DECAPx10_ASAP7_75t_R FILLER_293_238 ();
 DECAPx10_ASAP7_75t_R FILLER_293_260 ();
 DECAPx10_ASAP7_75t_R FILLER_293_282 ();
 DECAPx10_ASAP7_75t_R FILLER_293_304 ();
 DECAPx10_ASAP7_75t_R FILLER_293_326 ();
 DECAPx10_ASAP7_75t_R FILLER_293_348 ();
 DECAPx10_ASAP7_75t_R FILLER_293_370 ();
 DECAPx10_ASAP7_75t_R FILLER_293_392 ();
 DECAPx10_ASAP7_75t_R FILLER_293_414 ();
 DECAPx10_ASAP7_75t_R FILLER_293_436 ();
 DECAPx10_ASAP7_75t_R FILLER_293_458 ();
 DECAPx10_ASAP7_75t_R FILLER_293_480 ();
 DECAPx10_ASAP7_75t_R FILLER_293_502 ();
 DECAPx10_ASAP7_75t_R FILLER_293_524 ();
 DECAPx10_ASAP7_75t_R FILLER_293_546 ();
 DECAPx10_ASAP7_75t_R FILLER_293_568 ();
 DECAPx10_ASAP7_75t_R FILLER_293_590 ();
 DECAPx10_ASAP7_75t_R FILLER_293_612 ();
 DECAPx10_ASAP7_75t_R FILLER_293_634 ();
 DECAPx10_ASAP7_75t_R FILLER_293_656 ();
 DECAPx10_ASAP7_75t_R FILLER_293_678 ();
 DECAPx10_ASAP7_75t_R FILLER_293_700 ();
 DECAPx10_ASAP7_75t_R FILLER_293_722 ();
 DECAPx10_ASAP7_75t_R FILLER_293_744 ();
 DECAPx10_ASAP7_75t_R FILLER_293_766 ();
 DECAPx10_ASAP7_75t_R FILLER_293_788 ();
 DECAPx10_ASAP7_75t_R FILLER_293_810 ();
 DECAPx10_ASAP7_75t_R FILLER_293_832 ();
 DECAPx10_ASAP7_75t_R FILLER_293_854 ();
 DECAPx10_ASAP7_75t_R FILLER_293_876 ();
 DECAPx10_ASAP7_75t_R FILLER_293_898 ();
 DECAPx10_ASAP7_75t_R FILLER_293_920 ();
 DECAPx10_ASAP7_75t_R FILLER_293_942 ();
 DECAPx10_ASAP7_75t_R FILLER_293_964 ();
 DECAPx10_ASAP7_75t_R FILLER_293_986 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_293_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_293_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_293_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_293_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_294_172 ();
 DECAPx10_ASAP7_75t_R FILLER_294_194 ();
 DECAPx10_ASAP7_75t_R FILLER_294_216 ();
 DECAPx10_ASAP7_75t_R FILLER_294_238 ();
 DECAPx10_ASAP7_75t_R FILLER_294_260 ();
 DECAPx10_ASAP7_75t_R FILLER_294_282 ();
 DECAPx10_ASAP7_75t_R FILLER_294_304 ();
 DECAPx10_ASAP7_75t_R FILLER_294_326 ();
 DECAPx10_ASAP7_75t_R FILLER_294_348 ();
 DECAPx10_ASAP7_75t_R FILLER_294_370 ();
 DECAPx10_ASAP7_75t_R FILLER_294_392 ();
 DECAPx10_ASAP7_75t_R FILLER_294_414 ();
 DECAPx10_ASAP7_75t_R FILLER_294_436 ();
 DECAPx10_ASAP7_75t_R FILLER_294_458 ();
 DECAPx10_ASAP7_75t_R FILLER_294_480 ();
 DECAPx10_ASAP7_75t_R FILLER_294_502 ();
 DECAPx10_ASAP7_75t_R FILLER_294_524 ();
 DECAPx10_ASAP7_75t_R FILLER_294_546 ();
 DECAPx10_ASAP7_75t_R FILLER_294_568 ();
 DECAPx10_ASAP7_75t_R FILLER_294_590 ();
 DECAPx6_ASAP7_75t_R FILLER_294_612 ();
 DECAPx2_ASAP7_75t_R FILLER_294_626 ();
 DECAPx10_ASAP7_75t_R FILLER_294_634 ();
 DECAPx10_ASAP7_75t_R FILLER_294_656 ();
 DECAPx10_ASAP7_75t_R FILLER_294_678 ();
 DECAPx10_ASAP7_75t_R FILLER_294_700 ();
 DECAPx10_ASAP7_75t_R FILLER_294_722 ();
 DECAPx10_ASAP7_75t_R FILLER_294_744 ();
 DECAPx10_ASAP7_75t_R FILLER_294_766 ();
 DECAPx10_ASAP7_75t_R FILLER_294_788 ();
 DECAPx10_ASAP7_75t_R FILLER_294_810 ();
 DECAPx10_ASAP7_75t_R FILLER_294_832 ();
 DECAPx10_ASAP7_75t_R FILLER_294_854 ();
 DECAPx10_ASAP7_75t_R FILLER_294_876 ();
 DECAPx10_ASAP7_75t_R FILLER_294_898 ();
 DECAPx10_ASAP7_75t_R FILLER_294_920 ();
 DECAPx10_ASAP7_75t_R FILLER_294_942 ();
 DECAPx10_ASAP7_75t_R FILLER_294_964 ();
 DECAPx10_ASAP7_75t_R FILLER_294_986 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_294_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_294_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_294_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_294_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_1292 ();
endmodule
