VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA ibex_alu_via2_3_1600_480_1_5_320_320
  VIARULE M1M2_PR ;
  CUTSIZE 0.15 0.15 ;
  LAYERS met1 via met2 ;
  CUTSPACING 0.17 0.17 ;
  ENCLOSURE 0.085 0.165 0.055 0.085 ;
  ROWCOL 1 5 ;
END ibex_alu_via2_3_1600_480_1_5_320_320

VIA ibex_alu_via3_4_1600_480_1_4_400_400
  VIARULE M2M3_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met2 via2 met3 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.04 0.085 0.065 0.065 ;
  ROWCOL 1 4 ;
END ibex_alu_via3_4_1600_480_1_4_400_400

VIA ibex_alu_via4_5_1600_480_1_4_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.06 0.1 0.065 ;
  ROWCOL 1 4 ;
END ibex_alu_via4_5_1600_480_1_4_400_400

VIA ibex_alu_via5_6_1600_1600_1_1_1600_1600
  VIARULE M4M5_PR ;
  CUTSIZE 0.8 0.8 ;
  LAYERS met4 via4 met5 ;
  CUTSPACING 0.8 0.8 ;
  ENCLOSURE 0.4 0.19 0.31 0.4 ;
END ibex_alu_via5_6_1600_1600_1_1_1600_1600

MACRO ibex_alu
  FOREIGN ibex_alu 0 0 ;
  CLASS BLOCK ;
  SIZE 149.39 BY 149.39 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  27.72 137.92 137.88 139.52 ;
        RECT  27.72 110.72 137.88 112.32 ;
        RECT  27.72 83.52 137.88 85.12 ;
        RECT  27.72 56.32 137.88 57.92 ;
        RECT  27.72 29.12 137.88 30.72 ;
      LAYER met4 ;
        RECT  136.28 5.2 137.88 147.12 ;
        RECT  109.14 5.2 110.74 147.12 ;
        RECT  82 5.2 83.6 147.12 ;
        RECT  54.86 5.2 56.46 147.12 ;
        RECT  27.72 5.2 29.32 147.12 ;
      LAYER met1 ;
        RECT  1.38 146.64 148.12 147.12 ;
        RECT  1.38 141.2 148.12 141.68 ;
        RECT  1.38 135.76 148.12 136.24 ;
        RECT  1.38 130.32 148.12 130.8 ;
        RECT  1.38 124.88 148.12 125.36 ;
        RECT  1.38 119.44 148.12 119.92 ;
        RECT  1.38 114 148.12 114.48 ;
        RECT  1.38 108.56 148.12 109.04 ;
        RECT  1.38 103.12 148.12 103.6 ;
        RECT  1.38 97.68 148.12 98.16 ;
        RECT  1.38 92.24 148.12 92.72 ;
        RECT  1.38 86.8 148.12 87.28 ;
        RECT  1.38 81.36 148.12 81.84 ;
        RECT  1.38 75.92 148.12 76.4 ;
        RECT  1.38 70.48 148.12 70.96 ;
        RECT  1.38 65.04 148.12 65.52 ;
        RECT  1.38 59.6 148.12 60.08 ;
        RECT  1.38 54.16 148.12 54.64 ;
        RECT  1.38 48.72 148.12 49.2 ;
        RECT  1.38 43.28 148.12 43.76 ;
        RECT  1.38 37.84 148.12 38.32 ;
        RECT  1.38 32.4 148.12 32.88 ;
        RECT  1.38 26.96 148.12 27.44 ;
        RECT  1.38 21.52 148.12 22 ;
        RECT  1.38 16.08 148.12 16.56 ;
        RECT  1.38 10.64 148.12 11.12 ;
        RECT  1.38 5.2 148.12 5.68 ;
      VIA 137.08 138.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 111.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 84.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 57.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 29.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 138.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 111.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 84.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 57.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 29.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 138.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 111.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 84.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 57.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 29.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 138.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 111.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 84.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 57.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 29.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 138.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 111.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 84.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 57.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 29.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  136.29 146.715 137.87 147.045 ;
      VIA 137.08 146.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 146.695 137.85 147.065 ;
      VIA 137.08 146.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 146.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 141.275 137.87 141.605 ;
      VIA 137.08 141.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 141.255 137.85 141.625 ;
      VIA 137.08 141.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 141.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 135.835 137.87 136.165 ;
      VIA 137.08 136 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 135.815 137.85 136.185 ;
      VIA 137.08 136 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 136 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 130.395 137.87 130.725 ;
      VIA 137.08 130.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 130.375 137.85 130.745 ;
      VIA 137.08 130.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 130.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 124.955 137.87 125.285 ;
      VIA 137.08 125.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 124.935 137.85 125.305 ;
      VIA 137.08 125.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 125.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 119.515 137.87 119.845 ;
      VIA 137.08 119.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 119.495 137.85 119.865 ;
      VIA 137.08 119.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 119.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 114.075 137.87 114.405 ;
      VIA 137.08 114.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 114.055 137.85 114.425 ;
      VIA 137.08 114.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 114.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 108.635 137.87 108.965 ;
      VIA 137.08 108.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 108.615 137.85 108.985 ;
      VIA 137.08 108.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 108.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 103.195 137.87 103.525 ;
      VIA 137.08 103.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 103.175 137.85 103.545 ;
      VIA 137.08 103.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 103.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 97.755 137.87 98.085 ;
      VIA 137.08 97.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 97.735 137.85 98.105 ;
      VIA 137.08 97.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 97.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 92.315 137.87 92.645 ;
      VIA 137.08 92.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 92.295 137.85 92.665 ;
      VIA 137.08 92.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 92.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 86.875 137.87 87.205 ;
      VIA 137.08 87.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 86.855 137.85 87.225 ;
      VIA 137.08 87.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 87.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 81.435 137.87 81.765 ;
      VIA 137.08 81.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 81.415 137.85 81.785 ;
      VIA 137.08 81.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 81.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 75.995 137.87 76.325 ;
      VIA 137.08 76.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 75.975 137.85 76.345 ;
      VIA 137.08 76.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 76.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 70.555 137.87 70.885 ;
      VIA 137.08 70.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 70.535 137.85 70.905 ;
      VIA 137.08 70.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 70.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 65.115 137.87 65.445 ;
      VIA 137.08 65.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 65.095 137.85 65.465 ;
      VIA 137.08 65.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 65.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 59.675 137.87 60.005 ;
      VIA 137.08 59.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 59.655 137.85 60.025 ;
      VIA 137.08 59.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 59.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 54.235 137.87 54.565 ;
      VIA 137.08 54.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 54.215 137.85 54.585 ;
      VIA 137.08 54.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 54.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 48.795 137.87 49.125 ;
      VIA 137.08 48.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 48.775 137.85 49.145 ;
      VIA 137.08 48.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 48.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 43.355 137.87 43.685 ;
      VIA 137.08 43.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 43.335 137.85 43.705 ;
      VIA 137.08 43.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 43.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 37.915 137.87 38.245 ;
      VIA 137.08 38.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 37.895 137.85 38.265 ;
      VIA 137.08 38.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 38.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 32.475 137.87 32.805 ;
      VIA 137.08 32.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 32.455 137.85 32.825 ;
      VIA 137.08 32.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 32.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 27.035 137.87 27.365 ;
      VIA 137.08 27.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 27.015 137.85 27.385 ;
      VIA 137.08 27.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 27.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 21.595 137.87 21.925 ;
      VIA 137.08 21.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 21.575 137.85 21.945 ;
      VIA 137.08 21.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 21.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 16.155 137.87 16.485 ;
      VIA 137.08 16.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 16.135 137.85 16.505 ;
      VIA 137.08 16.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 16.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 10.715 137.87 11.045 ;
      VIA 137.08 10.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 10.695 137.85 11.065 ;
      VIA 137.08 10.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 10.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 5.275 137.87 5.605 ;
      VIA 137.08 5.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 5.255 137.85 5.625 ;
      VIA 137.08 5.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 5.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 146.715 110.73 147.045 ;
      VIA 109.94 146.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 146.695 110.71 147.065 ;
      VIA 109.94 146.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 146.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 141.275 110.73 141.605 ;
      VIA 109.94 141.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 141.255 110.71 141.625 ;
      VIA 109.94 141.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 141.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 135.835 110.73 136.165 ;
      VIA 109.94 136 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 135.815 110.71 136.185 ;
      VIA 109.94 136 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 136 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 130.395 110.73 130.725 ;
      VIA 109.94 130.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 130.375 110.71 130.745 ;
      VIA 109.94 130.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 130.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 124.955 110.73 125.285 ;
      VIA 109.94 125.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 124.935 110.71 125.305 ;
      VIA 109.94 125.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 125.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 119.515 110.73 119.845 ;
      VIA 109.94 119.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 119.495 110.71 119.865 ;
      VIA 109.94 119.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 119.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 114.075 110.73 114.405 ;
      VIA 109.94 114.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 114.055 110.71 114.425 ;
      VIA 109.94 114.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 114.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 108.635 110.73 108.965 ;
      VIA 109.94 108.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 108.615 110.71 108.985 ;
      VIA 109.94 108.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 108.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 103.195 110.73 103.525 ;
      VIA 109.94 103.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 103.175 110.71 103.545 ;
      VIA 109.94 103.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 103.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 97.755 110.73 98.085 ;
      VIA 109.94 97.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 97.735 110.71 98.105 ;
      VIA 109.94 97.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 97.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 92.315 110.73 92.645 ;
      VIA 109.94 92.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 92.295 110.71 92.665 ;
      VIA 109.94 92.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 92.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 86.875 110.73 87.205 ;
      VIA 109.94 87.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 86.855 110.71 87.225 ;
      VIA 109.94 87.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 87.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 81.435 110.73 81.765 ;
      VIA 109.94 81.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 81.415 110.71 81.785 ;
      VIA 109.94 81.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 81.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 75.995 110.73 76.325 ;
      VIA 109.94 76.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 75.975 110.71 76.345 ;
      VIA 109.94 76.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 76.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 70.555 110.73 70.885 ;
      VIA 109.94 70.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 70.535 110.71 70.905 ;
      VIA 109.94 70.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 70.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 65.115 110.73 65.445 ;
      VIA 109.94 65.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 65.095 110.71 65.465 ;
      VIA 109.94 65.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 65.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 59.675 110.73 60.005 ;
      VIA 109.94 59.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 59.655 110.71 60.025 ;
      VIA 109.94 59.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 59.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 54.235 110.73 54.565 ;
      VIA 109.94 54.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 54.215 110.71 54.585 ;
      VIA 109.94 54.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 54.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 48.795 110.73 49.125 ;
      VIA 109.94 48.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 48.775 110.71 49.145 ;
      VIA 109.94 48.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 48.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 43.355 110.73 43.685 ;
      VIA 109.94 43.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 43.335 110.71 43.705 ;
      VIA 109.94 43.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 43.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 37.915 110.73 38.245 ;
      VIA 109.94 38.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 37.895 110.71 38.265 ;
      VIA 109.94 38.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 38.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 32.475 110.73 32.805 ;
      VIA 109.94 32.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 32.455 110.71 32.825 ;
      VIA 109.94 32.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 32.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 27.035 110.73 27.365 ;
      VIA 109.94 27.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 27.015 110.71 27.385 ;
      VIA 109.94 27.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 27.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 21.595 110.73 21.925 ;
      VIA 109.94 21.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 21.575 110.71 21.945 ;
      VIA 109.94 21.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 21.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 16.155 110.73 16.485 ;
      VIA 109.94 16.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 16.135 110.71 16.505 ;
      VIA 109.94 16.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 16.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 10.715 110.73 11.045 ;
      VIA 109.94 10.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 10.695 110.71 11.065 ;
      VIA 109.94 10.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 10.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 5.275 110.73 5.605 ;
      VIA 109.94 5.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 5.255 110.71 5.625 ;
      VIA 109.94 5.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 5.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 146.715 83.59 147.045 ;
      VIA 82.8 146.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 146.695 83.57 147.065 ;
      VIA 82.8 146.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 146.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 141.275 83.59 141.605 ;
      VIA 82.8 141.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 141.255 83.57 141.625 ;
      VIA 82.8 141.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 141.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 135.835 83.59 136.165 ;
      VIA 82.8 136 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 135.815 83.57 136.185 ;
      VIA 82.8 136 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 136 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 130.395 83.59 130.725 ;
      VIA 82.8 130.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 130.375 83.57 130.745 ;
      VIA 82.8 130.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 130.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 124.955 83.59 125.285 ;
      VIA 82.8 125.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 124.935 83.57 125.305 ;
      VIA 82.8 125.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 125.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 119.515 83.59 119.845 ;
      VIA 82.8 119.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 119.495 83.57 119.865 ;
      VIA 82.8 119.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 119.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 114.075 83.59 114.405 ;
      VIA 82.8 114.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 114.055 83.57 114.425 ;
      VIA 82.8 114.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 114.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 108.635 83.59 108.965 ;
      VIA 82.8 108.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 108.615 83.57 108.985 ;
      VIA 82.8 108.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 108.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 103.195 83.59 103.525 ;
      VIA 82.8 103.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 103.175 83.57 103.545 ;
      VIA 82.8 103.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 103.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 97.755 83.59 98.085 ;
      VIA 82.8 97.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 97.735 83.57 98.105 ;
      VIA 82.8 97.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 97.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 92.315 83.59 92.645 ;
      VIA 82.8 92.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 92.295 83.57 92.665 ;
      VIA 82.8 92.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 92.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 86.875 83.59 87.205 ;
      VIA 82.8 87.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 86.855 83.57 87.225 ;
      VIA 82.8 87.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 87.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 81.435 83.59 81.765 ;
      VIA 82.8 81.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 81.415 83.57 81.785 ;
      VIA 82.8 81.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 81.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 75.995 83.59 76.325 ;
      VIA 82.8 76.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 75.975 83.57 76.345 ;
      VIA 82.8 76.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 76.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 70.555 83.59 70.885 ;
      VIA 82.8 70.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 70.535 83.57 70.905 ;
      VIA 82.8 70.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 70.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 65.115 83.59 65.445 ;
      VIA 82.8 65.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 65.095 83.57 65.465 ;
      VIA 82.8 65.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 65.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 59.675 83.59 60.005 ;
      VIA 82.8 59.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 59.655 83.57 60.025 ;
      VIA 82.8 59.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 59.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 54.235 83.59 54.565 ;
      VIA 82.8 54.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 54.215 83.57 54.585 ;
      VIA 82.8 54.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 54.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 48.795 83.59 49.125 ;
      VIA 82.8 48.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 48.775 83.57 49.145 ;
      VIA 82.8 48.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 48.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 43.355 83.59 43.685 ;
      VIA 82.8 43.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 43.335 83.57 43.705 ;
      VIA 82.8 43.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 43.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 37.915 83.59 38.245 ;
      VIA 82.8 38.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 37.895 83.57 38.265 ;
      VIA 82.8 38.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 38.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 32.475 83.59 32.805 ;
      VIA 82.8 32.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 32.455 83.57 32.825 ;
      VIA 82.8 32.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 32.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 27.035 83.59 27.365 ;
      VIA 82.8 27.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 27.015 83.57 27.385 ;
      VIA 82.8 27.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 27.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 21.595 83.59 21.925 ;
      VIA 82.8 21.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 21.575 83.57 21.945 ;
      VIA 82.8 21.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 21.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 16.155 83.59 16.485 ;
      VIA 82.8 16.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 16.135 83.57 16.505 ;
      VIA 82.8 16.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 16.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 10.715 83.59 11.045 ;
      VIA 82.8 10.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 10.695 83.57 11.065 ;
      VIA 82.8 10.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 10.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 5.275 83.59 5.605 ;
      VIA 82.8 5.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 5.255 83.57 5.625 ;
      VIA 82.8 5.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 5.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 146.715 56.45 147.045 ;
      VIA 55.66 146.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 146.695 56.43 147.065 ;
      VIA 55.66 146.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 146.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 141.275 56.45 141.605 ;
      VIA 55.66 141.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 141.255 56.43 141.625 ;
      VIA 55.66 141.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 141.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 135.835 56.45 136.165 ;
      VIA 55.66 136 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 135.815 56.43 136.185 ;
      VIA 55.66 136 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 136 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 130.395 56.45 130.725 ;
      VIA 55.66 130.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 130.375 56.43 130.745 ;
      VIA 55.66 130.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 130.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 124.955 56.45 125.285 ;
      VIA 55.66 125.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 124.935 56.43 125.305 ;
      VIA 55.66 125.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 125.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 119.515 56.45 119.845 ;
      VIA 55.66 119.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 119.495 56.43 119.865 ;
      VIA 55.66 119.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 119.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 114.075 56.45 114.405 ;
      VIA 55.66 114.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 114.055 56.43 114.425 ;
      VIA 55.66 114.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 114.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 108.635 56.45 108.965 ;
      VIA 55.66 108.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 108.615 56.43 108.985 ;
      VIA 55.66 108.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 108.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 103.195 56.45 103.525 ;
      VIA 55.66 103.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 103.175 56.43 103.545 ;
      VIA 55.66 103.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 103.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 97.755 56.45 98.085 ;
      VIA 55.66 97.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 97.735 56.43 98.105 ;
      VIA 55.66 97.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 97.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 92.315 56.45 92.645 ;
      VIA 55.66 92.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 92.295 56.43 92.665 ;
      VIA 55.66 92.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 92.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 86.875 56.45 87.205 ;
      VIA 55.66 87.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 86.855 56.43 87.225 ;
      VIA 55.66 87.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 87.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 81.435 56.45 81.765 ;
      VIA 55.66 81.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 81.415 56.43 81.785 ;
      VIA 55.66 81.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 81.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 75.995 56.45 76.325 ;
      VIA 55.66 76.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 75.975 56.43 76.345 ;
      VIA 55.66 76.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 76.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 70.555 56.45 70.885 ;
      VIA 55.66 70.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 70.535 56.43 70.905 ;
      VIA 55.66 70.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 70.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 65.115 56.45 65.445 ;
      VIA 55.66 65.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 65.095 56.43 65.465 ;
      VIA 55.66 65.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 65.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 59.675 56.45 60.005 ;
      VIA 55.66 59.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 59.655 56.43 60.025 ;
      VIA 55.66 59.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 59.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 54.235 56.45 54.565 ;
      VIA 55.66 54.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 54.215 56.43 54.585 ;
      VIA 55.66 54.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 54.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 48.795 56.45 49.125 ;
      VIA 55.66 48.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 48.775 56.43 49.145 ;
      VIA 55.66 48.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 48.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 43.355 56.45 43.685 ;
      VIA 55.66 43.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 43.335 56.43 43.705 ;
      VIA 55.66 43.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 43.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 37.915 56.45 38.245 ;
      VIA 55.66 38.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 37.895 56.43 38.265 ;
      VIA 55.66 38.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 38.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 32.475 56.45 32.805 ;
      VIA 55.66 32.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 32.455 56.43 32.825 ;
      VIA 55.66 32.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 32.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 27.035 56.45 27.365 ;
      VIA 55.66 27.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 27.015 56.43 27.385 ;
      VIA 55.66 27.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 27.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 21.595 56.45 21.925 ;
      VIA 55.66 21.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 21.575 56.43 21.945 ;
      VIA 55.66 21.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 21.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 16.155 56.45 16.485 ;
      VIA 55.66 16.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 16.135 56.43 16.505 ;
      VIA 55.66 16.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 16.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 10.715 56.45 11.045 ;
      VIA 55.66 10.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 10.695 56.43 11.065 ;
      VIA 55.66 10.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 10.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 5.275 56.45 5.605 ;
      VIA 55.66 5.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 5.255 56.43 5.625 ;
      VIA 55.66 5.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 5.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 146.715 29.31 147.045 ;
      VIA 28.52 146.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 146.695 29.29 147.065 ;
      VIA 28.52 146.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 146.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 141.275 29.31 141.605 ;
      VIA 28.52 141.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 141.255 29.29 141.625 ;
      VIA 28.52 141.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 141.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 135.835 29.31 136.165 ;
      VIA 28.52 136 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 135.815 29.29 136.185 ;
      VIA 28.52 136 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 136 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 130.395 29.31 130.725 ;
      VIA 28.52 130.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 130.375 29.29 130.745 ;
      VIA 28.52 130.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 130.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 124.955 29.31 125.285 ;
      VIA 28.52 125.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 124.935 29.29 125.305 ;
      VIA 28.52 125.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 125.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 119.515 29.31 119.845 ;
      VIA 28.52 119.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 119.495 29.29 119.865 ;
      VIA 28.52 119.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 119.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 114.075 29.31 114.405 ;
      VIA 28.52 114.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 114.055 29.29 114.425 ;
      VIA 28.52 114.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 114.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 108.635 29.31 108.965 ;
      VIA 28.52 108.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 108.615 29.29 108.985 ;
      VIA 28.52 108.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 108.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 103.195 29.31 103.525 ;
      VIA 28.52 103.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 103.175 29.29 103.545 ;
      VIA 28.52 103.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 103.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 97.755 29.31 98.085 ;
      VIA 28.52 97.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 97.735 29.29 98.105 ;
      VIA 28.52 97.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 97.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 92.315 29.31 92.645 ;
      VIA 28.52 92.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 92.295 29.29 92.665 ;
      VIA 28.52 92.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 92.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 86.875 29.31 87.205 ;
      VIA 28.52 87.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 86.855 29.29 87.225 ;
      VIA 28.52 87.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 87.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 81.435 29.31 81.765 ;
      VIA 28.52 81.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 81.415 29.29 81.785 ;
      VIA 28.52 81.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 81.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 75.995 29.31 76.325 ;
      VIA 28.52 76.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 75.975 29.29 76.345 ;
      VIA 28.52 76.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 76.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 70.555 29.31 70.885 ;
      VIA 28.52 70.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 70.535 29.29 70.905 ;
      VIA 28.52 70.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 70.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 65.115 29.31 65.445 ;
      VIA 28.52 65.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 65.095 29.29 65.465 ;
      VIA 28.52 65.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 65.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 59.675 29.31 60.005 ;
      VIA 28.52 59.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 59.655 29.29 60.025 ;
      VIA 28.52 59.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 59.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 54.235 29.31 54.565 ;
      VIA 28.52 54.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 54.215 29.29 54.585 ;
      VIA 28.52 54.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 54.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 48.795 29.31 49.125 ;
      VIA 28.52 48.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 48.775 29.29 49.145 ;
      VIA 28.52 48.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 48.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 43.355 29.31 43.685 ;
      VIA 28.52 43.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 43.335 29.29 43.705 ;
      VIA 28.52 43.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 43.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 37.915 29.31 38.245 ;
      VIA 28.52 38.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 37.895 29.29 38.265 ;
      VIA 28.52 38.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 38.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 32.475 29.31 32.805 ;
      VIA 28.52 32.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 32.455 29.29 32.825 ;
      VIA 28.52 32.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 32.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 27.035 29.31 27.365 ;
      VIA 28.52 27.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 27.015 29.29 27.385 ;
      VIA 28.52 27.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 27.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 21.595 29.31 21.925 ;
      VIA 28.52 21.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 21.575 29.29 21.945 ;
      VIA 28.52 21.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 21.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 16.155 29.31 16.485 ;
      VIA 28.52 16.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 16.135 29.29 16.505 ;
      VIA 28.52 16.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 16.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 10.715 29.31 11.045 ;
      VIA 28.52 10.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 10.695 29.29 11.065 ;
      VIA 28.52 10.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 10.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 5.275 29.31 5.605 ;
      VIA 28.52 5.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 5.255 29.29 5.625 ;
      VIA 28.52 5.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 5.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  14.15 124.32 124.31 125.92 ;
        RECT  14.15 97.12 124.31 98.72 ;
        RECT  14.15 69.92 124.31 71.52 ;
        RECT  14.15 42.72 124.31 44.32 ;
        RECT  14.15 15.52 124.31 17.12 ;
      LAYER met4 ;
        RECT  122.71 2.48 124.31 144.4 ;
        RECT  95.57 2.48 97.17 144.4 ;
        RECT  68.43 2.48 70.03 144.4 ;
        RECT  41.29 2.48 42.89 144.4 ;
        RECT  14.15 2.48 15.75 144.4 ;
      LAYER met1 ;
        RECT  1.38 143.92 148.12 144.4 ;
        RECT  1.38 138.48 148.12 138.96 ;
        RECT  1.38 133.04 148.12 133.52 ;
        RECT  1.38 127.6 148.12 128.08 ;
        RECT  1.38 122.16 148.12 122.64 ;
        RECT  1.38 116.72 148.12 117.2 ;
        RECT  1.38 111.28 148.12 111.76 ;
        RECT  1.38 105.84 148.12 106.32 ;
        RECT  1.38 100.4 148.12 100.88 ;
        RECT  1.38 94.96 148.12 95.44 ;
        RECT  1.38 89.52 148.12 90 ;
        RECT  1.38 84.08 148.12 84.56 ;
        RECT  1.38 78.64 148.12 79.12 ;
        RECT  1.38 73.2 148.12 73.68 ;
        RECT  1.38 67.76 148.12 68.24 ;
        RECT  1.38 62.32 148.12 62.8 ;
        RECT  1.38 56.88 148.12 57.36 ;
        RECT  1.38 51.44 148.12 51.92 ;
        RECT  1.38 46 148.12 46.48 ;
        RECT  1.38 40.56 148.12 41.04 ;
        RECT  1.38 35.12 148.12 35.6 ;
        RECT  1.38 29.68 148.12 30.16 ;
        RECT  1.38 24.24 148.12 24.72 ;
        RECT  1.38 18.8 148.12 19.28 ;
        RECT  1.38 13.36 148.12 13.84 ;
        RECT  1.38 7.92 148.12 8.4 ;
        RECT  1.38 2.48 148.12 2.96 ;
      VIA 123.51 125.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 97.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 70.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 43.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 16.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 125.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 97.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 70.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 43.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 16.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 125.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 97.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 70.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 43.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 16.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 125.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 97.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 70.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 43.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 16.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 125.12 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 97.92 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 70.72 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 43.52 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 16.32 ibex_alu_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  122.72 143.995 124.3 144.325 ;
      VIA 123.51 144.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 143.975 124.28 144.345 ;
      VIA 123.51 144.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 144.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 138.555 124.3 138.885 ;
      VIA 123.51 138.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 138.535 124.28 138.905 ;
      VIA 123.51 138.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 138.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 133.115 124.3 133.445 ;
      VIA 123.51 133.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 133.095 124.28 133.465 ;
      VIA 123.51 133.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 133.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 127.675 124.3 128.005 ;
      VIA 123.51 127.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 127.655 124.28 128.025 ;
      VIA 123.51 127.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 127.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 122.235 124.3 122.565 ;
      VIA 123.51 122.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 122.215 124.28 122.585 ;
      VIA 123.51 122.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 122.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 116.795 124.3 117.125 ;
      VIA 123.51 116.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 116.775 124.28 117.145 ;
      VIA 123.51 116.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 116.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 111.355 124.3 111.685 ;
      VIA 123.51 111.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 111.335 124.28 111.705 ;
      VIA 123.51 111.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 111.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 105.915 124.3 106.245 ;
      VIA 123.51 106.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 105.895 124.28 106.265 ;
      VIA 123.51 106.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 106.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 100.475 124.3 100.805 ;
      VIA 123.51 100.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 100.455 124.28 100.825 ;
      VIA 123.51 100.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 100.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 95.035 124.3 95.365 ;
      VIA 123.51 95.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 95.015 124.28 95.385 ;
      VIA 123.51 95.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 95.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 89.595 124.3 89.925 ;
      VIA 123.51 89.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 89.575 124.28 89.945 ;
      VIA 123.51 89.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 89.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 84.155 124.3 84.485 ;
      VIA 123.51 84.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 84.135 124.28 84.505 ;
      VIA 123.51 84.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 84.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 78.715 124.3 79.045 ;
      VIA 123.51 78.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 78.695 124.28 79.065 ;
      VIA 123.51 78.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 78.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 73.275 124.3 73.605 ;
      VIA 123.51 73.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 73.255 124.28 73.625 ;
      VIA 123.51 73.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 73.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 67.835 124.3 68.165 ;
      VIA 123.51 68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 67.815 124.28 68.185 ;
      VIA 123.51 68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 62.395 124.3 62.725 ;
      VIA 123.51 62.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 62.375 124.28 62.745 ;
      VIA 123.51 62.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 62.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 56.955 124.3 57.285 ;
      VIA 123.51 57.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 56.935 124.28 57.305 ;
      VIA 123.51 57.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 57.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 51.515 124.3 51.845 ;
      VIA 123.51 51.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 51.495 124.28 51.865 ;
      VIA 123.51 51.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 51.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 46.075 124.3 46.405 ;
      VIA 123.51 46.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 46.055 124.28 46.425 ;
      VIA 123.51 46.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 46.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 40.635 124.3 40.965 ;
      VIA 123.51 40.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 40.615 124.28 40.985 ;
      VIA 123.51 40.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 40.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 35.195 124.3 35.525 ;
      VIA 123.51 35.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 35.175 124.28 35.545 ;
      VIA 123.51 35.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 35.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 29.755 124.3 30.085 ;
      VIA 123.51 29.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 29.735 124.28 30.105 ;
      VIA 123.51 29.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 29.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 24.315 124.3 24.645 ;
      VIA 123.51 24.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 24.295 124.28 24.665 ;
      VIA 123.51 24.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 24.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 18.875 124.3 19.205 ;
      VIA 123.51 19.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 18.855 124.28 19.225 ;
      VIA 123.51 19.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 19.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 13.435 124.3 13.765 ;
      VIA 123.51 13.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 13.415 124.28 13.785 ;
      VIA 123.51 13.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 13.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 7.995 124.3 8.325 ;
      VIA 123.51 8.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 7.975 124.28 8.345 ;
      VIA 123.51 8.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 8.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 2.555 124.3 2.885 ;
      VIA 123.51 2.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 2.535 124.28 2.905 ;
      VIA 123.51 2.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 2.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 143.995 97.16 144.325 ;
      VIA 96.37 144.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 143.975 97.14 144.345 ;
      VIA 96.37 144.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 144.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 138.555 97.16 138.885 ;
      VIA 96.37 138.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 138.535 97.14 138.905 ;
      VIA 96.37 138.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 138.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 133.115 97.16 133.445 ;
      VIA 96.37 133.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 133.095 97.14 133.465 ;
      VIA 96.37 133.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 133.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 127.675 97.16 128.005 ;
      VIA 96.37 127.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 127.655 97.14 128.025 ;
      VIA 96.37 127.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 127.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 122.235 97.16 122.565 ;
      VIA 96.37 122.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 122.215 97.14 122.585 ;
      VIA 96.37 122.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 122.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 116.795 97.16 117.125 ;
      VIA 96.37 116.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 116.775 97.14 117.145 ;
      VIA 96.37 116.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 116.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 111.355 97.16 111.685 ;
      VIA 96.37 111.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 111.335 97.14 111.705 ;
      VIA 96.37 111.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 111.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 105.915 97.16 106.245 ;
      VIA 96.37 106.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 105.895 97.14 106.265 ;
      VIA 96.37 106.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 106.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 100.475 97.16 100.805 ;
      VIA 96.37 100.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 100.455 97.14 100.825 ;
      VIA 96.37 100.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 100.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 95.035 97.16 95.365 ;
      VIA 96.37 95.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 95.015 97.14 95.385 ;
      VIA 96.37 95.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 95.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 89.595 97.16 89.925 ;
      VIA 96.37 89.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 89.575 97.14 89.945 ;
      VIA 96.37 89.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 89.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 84.155 97.16 84.485 ;
      VIA 96.37 84.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 84.135 97.14 84.505 ;
      VIA 96.37 84.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 84.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 78.715 97.16 79.045 ;
      VIA 96.37 78.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 78.695 97.14 79.065 ;
      VIA 96.37 78.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 78.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 73.275 97.16 73.605 ;
      VIA 96.37 73.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 73.255 97.14 73.625 ;
      VIA 96.37 73.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 73.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 67.835 97.16 68.165 ;
      VIA 96.37 68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 67.815 97.14 68.185 ;
      VIA 96.37 68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 62.395 97.16 62.725 ;
      VIA 96.37 62.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 62.375 97.14 62.745 ;
      VIA 96.37 62.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 62.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 56.955 97.16 57.285 ;
      VIA 96.37 57.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 56.935 97.14 57.305 ;
      VIA 96.37 57.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 57.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 51.515 97.16 51.845 ;
      VIA 96.37 51.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 51.495 97.14 51.865 ;
      VIA 96.37 51.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 51.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 46.075 97.16 46.405 ;
      VIA 96.37 46.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 46.055 97.14 46.425 ;
      VIA 96.37 46.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 46.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 40.635 97.16 40.965 ;
      VIA 96.37 40.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 40.615 97.14 40.985 ;
      VIA 96.37 40.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 40.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 35.195 97.16 35.525 ;
      VIA 96.37 35.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 35.175 97.14 35.545 ;
      VIA 96.37 35.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 35.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 29.755 97.16 30.085 ;
      VIA 96.37 29.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 29.735 97.14 30.105 ;
      VIA 96.37 29.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 29.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 24.315 97.16 24.645 ;
      VIA 96.37 24.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 24.295 97.14 24.665 ;
      VIA 96.37 24.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 24.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 18.875 97.16 19.205 ;
      VIA 96.37 19.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 18.855 97.14 19.225 ;
      VIA 96.37 19.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 19.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 13.435 97.16 13.765 ;
      VIA 96.37 13.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 13.415 97.14 13.785 ;
      VIA 96.37 13.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 13.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 7.995 97.16 8.325 ;
      VIA 96.37 8.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 7.975 97.14 8.345 ;
      VIA 96.37 8.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 8.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 2.555 97.16 2.885 ;
      VIA 96.37 2.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 2.535 97.14 2.905 ;
      VIA 96.37 2.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 2.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 143.995 70.02 144.325 ;
      VIA 69.23 144.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 143.975 70 144.345 ;
      VIA 69.23 144.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 144.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 138.555 70.02 138.885 ;
      VIA 69.23 138.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 138.535 70 138.905 ;
      VIA 69.23 138.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 138.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 133.115 70.02 133.445 ;
      VIA 69.23 133.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 133.095 70 133.465 ;
      VIA 69.23 133.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 133.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 127.675 70.02 128.005 ;
      VIA 69.23 127.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 127.655 70 128.025 ;
      VIA 69.23 127.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 127.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 122.235 70.02 122.565 ;
      VIA 69.23 122.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 122.215 70 122.585 ;
      VIA 69.23 122.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 122.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 116.795 70.02 117.125 ;
      VIA 69.23 116.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 116.775 70 117.145 ;
      VIA 69.23 116.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 116.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 111.355 70.02 111.685 ;
      VIA 69.23 111.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 111.335 70 111.705 ;
      VIA 69.23 111.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 111.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 105.915 70.02 106.245 ;
      VIA 69.23 106.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 105.895 70 106.265 ;
      VIA 69.23 106.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 106.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 100.475 70.02 100.805 ;
      VIA 69.23 100.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 100.455 70 100.825 ;
      VIA 69.23 100.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 100.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 95.035 70.02 95.365 ;
      VIA 69.23 95.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 95.015 70 95.385 ;
      VIA 69.23 95.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 95.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 89.595 70.02 89.925 ;
      VIA 69.23 89.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 89.575 70 89.945 ;
      VIA 69.23 89.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 89.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 84.155 70.02 84.485 ;
      VIA 69.23 84.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 84.135 70 84.505 ;
      VIA 69.23 84.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 84.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 78.715 70.02 79.045 ;
      VIA 69.23 78.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 78.695 70 79.065 ;
      VIA 69.23 78.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 78.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 73.275 70.02 73.605 ;
      VIA 69.23 73.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 73.255 70 73.625 ;
      VIA 69.23 73.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 73.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 67.835 70.02 68.165 ;
      VIA 69.23 68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 67.815 70 68.185 ;
      VIA 69.23 68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 62.395 70.02 62.725 ;
      VIA 69.23 62.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 62.375 70 62.745 ;
      VIA 69.23 62.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 62.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 56.955 70.02 57.285 ;
      VIA 69.23 57.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 56.935 70 57.305 ;
      VIA 69.23 57.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 57.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 51.515 70.02 51.845 ;
      VIA 69.23 51.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 51.495 70 51.865 ;
      VIA 69.23 51.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 51.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 46.075 70.02 46.405 ;
      VIA 69.23 46.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 46.055 70 46.425 ;
      VIA 69.23 46.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 46.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 40.635 70.02 40.965 ;
      VIA 69.23 40.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 40.615 70 40.985 ;
      VIA 69.23 40.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 40.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 35.195 70.02 35.525 ;
      VIA 69.23 35.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 35.175 70 35.545 ;
      VIA 69.23 35.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 35.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 29.755 70.02 30.085 ;
      VIA 69.23 29.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 29.735 70 30.105 ;
      VIA 69.23 29.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 29.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 24.315 70.02 24.645 ;
      VIA 69.23 24.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 24.295 70 24.665 ;
      VIA 69.23 24.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 24.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 18.875 70.02 19.205 ;
      VIA 69.23 19.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 18.855 70 19.225 ;
      VIA 69.23 19.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 19.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 13.435 70.02 13.765 ;
      VIA 69.23 13.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 13.415 70 13.785 ;
      VIA 69.23 13.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 13.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 7.995 70.02 8.325 ;
      VIA 69.23 8.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 7.975 70 8.345 ;
      VIA 69.23 8.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 8.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 2.555 70.02 2.885 ;
      VIA 69.23 2.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 2.535 70 2.905 ;
      VIA 69.23 2.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 2.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 143.995 42.88 144.325 ;
      VIA 42.09 144.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 143.975 42.86 144.345 ;
      VIA 42.09 144.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 144.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 138.555 42.88 138.885 ;
      VIA 42.09 138.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 138.535 42.86 138.905 ;
      VIA 42.09 138.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 138.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 133.115 42.88 133.445 ;
      VIA 42.09 133.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 133.095 42.86 133.465 ;
      VIA 42.09 133.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 133.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 127.675 42.88 128.005 ;
      VIA 42.09 127.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 127.655 42.86 128.025 ;
      VIA 42.09 127.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 127.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 122.235 42.88 122.565 ;
      VIA 42.09 122.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 122.215 42.86 122.585 ;
      VIA 42.09 122.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 122.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 116.795 42.88 117.125 ;
      VIA 42.09 116.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 116.775 42.86 117.145 ;
      VIA 42.09 116.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 116.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 111.355 42.88 111.685 ;
      VIA 42.09 111.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 111.335 42.86 111.705 ;
      VIA 42.09 111.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 111.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 105.915 42.88 106.245 ;
      VIA 42.09 106.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 105.895 42.86 106.265 ;
      VIA 42.09 106.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 106.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 100.475 42.88 100.805 ;
      VIA 42.09 100.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 100.455 42.86 100.825 ;
      VIA 42.09 100.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 100.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 95.035 42.88 95.365 ;
      VIA 42.09 95.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 95.015 42.86 95.385 ;
      VIA 42.09 95.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 95.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 89.595 42.88 89.925 ;
      VIA 42.09 89.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 89.575 42.86 89.945 ;
      VIA 42.09 89.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 89.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 84.155 42.88 84.485 ;
      VIA 42.09 84.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 84.135 42.86 84.505 ;
      VIA 42.09 84.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 84.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 78.715 42.88 79.045 ;
      VIA 42.09 78.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 78.695 42.86 79.065 ;
      VIA 42.09 78.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 78.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 73.275 42.88 73.605 ;
      VIA 42.09 73.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 73.255 42.86 73.625 ;
      VIA 42.09 73.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 73.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 67.835 42.88 68.165 ;
      VIA 42.09 68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 67.815 42.86 68.185 ;
      VIA 42.09 68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 62.395 42.88 62.725 ;
      VIA 42.09 62.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 62.375 42.86 62.745 ;
      VIA 42.09 62.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 62.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 56.955 42.88 57.285 ;
      VIA 42.09 57.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 56.935 42.86 57.305 ;
      VIA 42.09 57.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 57.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 51.515 42.88 51.845 ;
      VIA 42.09 51.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 51.495 42.86 51.865 ;
      VIA 42.09 51.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 51.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 46.075 42.88 46.405 ;
      VIA 42.09 46.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 46.055 42.86 46.425 ;
      VIA 42.09 46.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 46.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 40.635 42.88 40.965 ;
      VIA 42.09 40.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 40.615 42.86 40.985 ;
      VIA 42.09 40.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 40.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 35.195 42.88 35.525 ;
      VIA 42.09 35.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 35.175 42.86 35.545 ;
      VIA 42.09 35.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 35.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 29.755 42.88 30.085 ;
      VIA 42.09 29.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 29.735 42.86 30.105 ;
      VIA 42.09 29.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 29.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 24.315 42.88 24.645 ;
      VIA 42.09 24.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 24.295 42.86 24.665 ;
      VIA 42.09 24.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 24.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 18.875 42.88 19.205 ;
      VIA 42.09 19.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 18.855 42.86 19.225 ;
      VIA 42.09 19.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 19.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 13.435 42.88 13.765 ;
      VIA 42.09 13.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 13.415 42.86 13.785 ;
      VIA 42.09 13.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 13.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 7.995 42.88 8.325 ;
      VIA 42.09 8.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 7.975 42.86 8.345 ;
      VIA 42.09 8.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 8.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 2.555 42.88 2.885 ;
      VIA 42.09 2.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 2.535 42.86 2.905 ;
      VIA 42.09 2.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 2.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 143.995 15.74 144.325 ;
      VIA 14.95 144.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 143.975 15.72 144.345 ;
      VIA 14.95 144.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 144.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 138.555 15.74 138.885 ;
      VIA 14.95 138.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 138.535 15.72 138.905 ;
      VIA 14.95 138.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 138.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 133.115 15.74 133.445 ;
      VIA 14.95 133.28 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 133.095 15.72 133.465 ;
      VIA 14.95 133.28 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 133.28 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 127.675 15.74 128.005 ;
      VIA 14.95 127.84 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 127.655 15.72 128.025 ;
      VIA 14.95 127.84 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 127.84 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 122.235 15.74 122.565 ;
      VIA 14.95 122.4 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 122.215 15.72 122.585 ;
      VIA 14.95 122.4 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 122.4 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 116.795 15.74 117.125 ;
      VIA 14.95 116.96 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 116.775 15.72 117.145 ;
      VIA 14.95 116.96 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 116.96 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 111.355 15.74 111.685 ;
      VIA 14.95 111.52 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 111.335 15.72 111.705 ;
      VIA 14.95 111.52 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 111.52 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 105.915 15.74 106.245 ;
      VIA 14.95 106.08 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 105.895 15.72 106.265 ;
      VIA 14.95 106.08 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 106.08 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 100.475 15.74 100.805 ;
      VIA 14.95 100.64 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 100.455 15.72 100.825 ;
      VIA 14.95 100.64 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 100.64 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 95.035 15.74 95.365 ;
      VIA 14.95 95.2 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 95.015 15.72 95.385 ;
      VIA 14.95 95.2 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 95.2 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 89.595 15.74 89.925 ;
      VIA 14.95 89.76 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 89.575 15.72 89.945 ;
      VIA 14.95 89.76 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 89.76 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 84.155 15.74 84.485 ;
      VIA 14.95 84.32 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 84.135 15.72 84.505 ;
      VIA 14.95 84.32 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 84.32 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 78.715 15.74 79.045 ;
      VIA 14.95 78.88 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 78.695 15.72 79.065 ;
      VIA 14.95 78.88 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 78.88 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 73.275 15.74 73.605 ;
      VIA 14.95 73.44 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 73.255 15.72 73.625 ;
      VIA 14.95 73.44 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 73.44 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 67.835 15.74 68.165 ;
      VIA 14.95 68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 67.815 15.72 68.185 ;
      VIA 14.95 68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 62.395 15.74 62.725 ;
      VIA 14.95 62.56 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 62.375 15.72 62.745 ;
      VIA 14.95 62.56 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 62.56 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 56.955 15.74 57.285 ;
      VIA 14.95 57.12 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 56.935 15.72 57.305 ;
      VIA 14.95 57.12 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 57.12 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 51.515 15.74 51.845 ;
      VIA 14.95 51.68 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 51.495 15.72 51.865 ;
      VIA 14.95 51.68 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 51.68 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 46.075 15.74 46.405 ;
      VIA 14.95 46.24 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 46.055 15.72 46.425 ;
      VIA 14.95 46.24 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 46.24 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 40.635 15.74 40.965 ;
      VIA 14.95 40.8 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 40.615 15.72 40.985 ;
      VIA 14.95 40.8 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 40.8 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 35.195 15.74 35.525 ;
      VIA 14.95 35.36 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 35.175 15.72 35.545 ;
      VIA 14.95 35.36 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 35.36 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 29.755 15.74 30.085 ;
      VIA 14.95 29.92 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 29.735 15.72 30.105 ;
      VIA 14.95 29.92 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 29.92 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 24.315 15.74 24.645 ;
      VIA 14.95 24.48 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 24.295 15.72 24.665 ;
      VIA 14.95 24.48 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 24.48 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 18.875 15.74 19.205 ;
      VIA 14.95 19.04 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 18.855 15.72 19.225 ;
      VIA 14.95 19.04 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 19.04 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 13.435 15.74 13.765 ;
      VIA 14.95 13.6 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 13.415 15.72 13.785 ;
      VIA 14.95 13.6 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 13.6 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 7.995 15.74 8.325 ;
      VIA 14.95 8.16 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 7.975 15.72 8.345 ;
      VIA 14.95 8.16 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 8.16 ibex_alu_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 2.555 15.74 2.885 ;
      VIA 14.95 2.72 ibex_alu_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 2.535 15.72 2.905 ;
      VIA 14.95 2.72 ibex_alu_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 2.72 ibex_alu_via2_3_1600_480_1_5_320_320 ;
    END
  END VSS
  PIN adder_result_ext_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 20.59 149.39 20.89 ;
    END
  END adder_result_ext_o[0]
  PIN adder_result_ext_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.16 0 92.3 0.485 ;
    END
  END adder_result_ext_o[10]
  PIN adder_result_ext_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  63.64 0 63.78 0.485 ;
    END
  END adder_result_ext_o[11]
  PIN adder_result_ext_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  54.44 0 54.58 0.485 ;
    END
  END adder_result_ext_o[12]
  PIN adder_result_ext_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 8.35 0.8 8.65 ;
    END
  END adder_result_ext_o[13]
  PIN adder_result_ext_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  53.52 0 53.66 0.485 ;
    END
  END adder_result_ext_o[14]
  PIN adder_result_ext_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.96 0 60.1 0.485 ;
    END
  END adder_result_ext_o[15]
  PIN adder_result_ext_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 19.23 0.8 19.53 ;
    END
  END adder_result_ext_o[16]
  PIN adder_result_ext_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 35.55 0.8 35.85 ;
    END
  END adder_result_ext_o[17]
  PIN adder_result_ext_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 13.79 0.8 14.09 ;
    END
  END adder_result_ext_o[18]
  PIN adder_result_ext_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 12.43 0.8 12.73 ;
    END
  END adder_result_ext_o[19]
  PIN adder_result_ext_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 99.47 149.39 99.77 ;
    END
  END adder_result_ext_o[1]
  PIN adder_result_ext_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  46.16 0 46.3 0.485 ;
    END
  END adder_result_ext_o[20]
  PIN adder_result_ext_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  26.84 0 26.98 0.485 ;
    END
  END adder_result_ext_o[21]
  PIN adder_result_ext_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  55.36 0 55.5 0.485 ;
    END
  END adder_result_ext_o[22]
  PIN adder_result_ext_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 0 73.9 0.485 ;
    END
  END adder_result_ext_o[23]
  PIN adder_result_ext_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  75.6 0 75.74 0.485 ;
    END
  END adder_result_ext_o[24]
  PIN adder_result_ext_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  95.84 0 95.98 0.485 ;
    END
  END adder_result_ext_o[25]
  PIN adder_result_ext_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.56 0 64.7 0.485 ;
    END
  END adder_result_ext_o[26]
  PIN adder_result_ext_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  101.36 0 101.5 0.485 ;
    END
  END adder_result_ext_o[27]
  PIN adder_result_ext_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  85.72 0 85.86 0.485 ;
    END
  END adder_result_ext_o[28]
  PIN adder_result_ext_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  104.12 0 104.26 0.485 ;
    END
  END adder_result_ext_o[29]
  PIN adder_result_ext_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 79.07 149.39 79.37 ;
    END
  END adder_result_ext_o[2]
  PIN adder_result_ext_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.52 0 99.66 0.485 ;
    END
  END adder_result_ext_o[30]
  PIN adder_result_ext_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 21.95 149.39 22.25 ;
    END
  END adder_result_ext_o[31]
  PIN adder_result_ext_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 92.67 149.39 92.97 ;
    END
  END adder_result_ext_o[32]
  PIN adder_result_ext_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 26.03 149.39 26.33 ;
    END
  END adder_result_ext_o[33]
  PIN adder_result_ext_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 36.91 149.39 37.21 ;
    END
  END adder_result_ext_o[3]
  PIN adder_result_ext_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 35.55 149.39 35.85 ;
    END
  END adder_result_ext_o[4]
  PIN adder_result_ext_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 83.15 149.39 83.45 ;
    END
  END adder_result_ext_o[5]
  PIN adder_result_ext_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  96.76 0 96.9 0.485 ;
    END
  END adder_result_ext_o[6]
  PIN adder_result_ext_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  79.28 0 79.42 0.485 ;
    END
  END adder_result_ext_o[7]
  PIN adder_result_ext_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 65.47 149.39 65.77 ;
    END
  END adder_result_ext_o[8]
  PIN adder_result_ext_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  69.16 0 69.3 0.485 ;
    END
  END adder_result_ext_o[9]
  PIN adder_result_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 51.87 149.39 52.17 ;
    END
  END adder_result_o[0]
  PIN adder_result_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71 0 71.14 0.485 ;
    END
  END adder_result_o[10]
  PIN adder_result_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.04 0 59.18 0.485 ;
    END
  END adder_result_o[11]
  PIN adder_result_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 83.15 0.8 83.45 ;
    END
  END adder_result_o[12]
  PIN adder_result_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 84.51 0.8 84.81 ;
    END
  END adder_result_o[13]
  PIN adder_result_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  62.72 0 62.86 0.485 ;
    END
  END adder_result_o[14]
  PIN adder_result_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 88.59 0.8 88.89 ;
    END
  END adder_result_o[15]
  PIN adder_result_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 89.95 0.8 90.25 ;
    END
  END adder_result_o[16]
  PIN adder_result_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 66.83 0.8 67.13 ;
    END
  END adder_result_o[17]
  PIN adder_result_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 30.11 0.8 30.41 ;
    END
  END adder_result_o[18]
  PIN adder_result_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 91.31 0.8 91.61 ;
    END
  END adder_result_o[19]
  PIN adder_result_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 62.75 149.39 63.05 ;
    END
  END adder_result_o[1]
  PIN adder_result_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  34.2 0 34.34 0.485 ;
    END
  END adder_result_o[20]
  PIN adder_result_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  60.88 0 61.02 0.485 ;
    END
  END adder_result_o[21]
  PIN adder_result_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  74.68 0 74.82 0.485 ;
    END
  END adder_result_o[22]
  PIN adder_result_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  77.44 0 77.58 0.485 ;
    END
  END adder_result_o[23]
  PIN adder_result_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94.92 0 95.06 0.485 ;
    END
  END adder_result_o[24]
  PIN adder_result_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  70.08 0 70.22 0.485 ;
    END
  END adder_result_o[25]
  PIN adder_result_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  97.68 0 97.82 0.485 ;
    END
  END adder_result_o[26]
  PIN adder_result_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  91.24 0 91.38 0.485 ;
    END
  END adder_result_o[27]
  PIN adder_result_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  111.48 0 111.62 0.485 ;
    END
  END adder_result_o[28]
  PIN adder_result_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  98.6 0 98.74 0.485 ;
    END
  END adder_result_o[29]
  PIN adder_result_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 45.07 149.39 45.37 ;
    END
  END adder_result_o[2]
  PIN adder_result_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 24.67 149.39 24.97 ;
    END
  END adder_result_o[30]
  PIN adder_result_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 61.39 149.39 61.69 ;
    END
  END adder_result_o[31]
  PIN adder_result_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 34.19 149.39 34.49 ;
    END
  END adder_result_o[3]
  PIN adder_result_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 47.79 149.39 48.09 ;
    END
  END adder_result_o[4]
  PIN adder_result_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  100.44 0 100.58 0.485 ;
    END
  END adder_result_o[5]
  PIN adder_result_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  80.2 0 80.34 0.485 ;
    END
  END adder_result_o[6]
  PIN adder_result_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94 0 94.14 0.485 ;
    END
  END adder_result_o[7]
  PIN adder_result_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  72.84 0 72.98 0.485 ;
    END
  END adder_result_o[8]
  PIN adder_result_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  93.08 0 93.22 0.485 ;
    END
  END adder_result_o[9]
  PIN comparison_result_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 87.23 149.39 87.53 ;
    END
  END comparison_result_o
  PIN imd_val_d_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 147.07 0.8 147.37 ;
    END
  END imd_val_d_o[0]
  PIN imd_val_d_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  15.8 148.905 15.94 149.39 ;
    END
  END imd_val_d_o[10]
  PIN imd_val_d_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.96 148.905 14.1 149.39 ;
    END
  END imd_val_d_o[11]
  PIN imd_val_d_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 136.19 0.8 136.49 ;
    END
  END imd_val_d_o[12]
  PIN imd_val_d_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 92.67 0.8 92.97 ;
    END
  END imd_val_d_o[13]
  PIN imd_val_d_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 106.27 0.8 106.57 ;
    END
  END imd_val_d_o[14]
  PIN imd_val_d_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 114.43 0.8 114.73 ;
    END
  END imd_val_d_o[15]
  PIN imd_val_d_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  17.64 148.905 17.78 149.39 ;
    END
  END imd_val_d_o[16]
  PIN imd_val_d_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 137.55 0.8 137.85 ;
    END
  END imd_val_d_o[17]
  PIN imd_val_d_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 148.905 18.7 149.39 ;
    END
  END imd_val_d_o[18]
  PIN imd_val_d_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 98.11 0.8 98.41 ;
    END
  END imd_val_d_o[19]
  PIN imd_val_d_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  14.88 148.905 15.02 149.39 ;
    END
  END imd_val_d_o[1]
  PIN imd_val_d_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  32.36 148.905 32.5 149.39 ;
    END
  END imd_val_d_o[20]
  PIN imd_val_d_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 117.15 0.8 117.45 ;
    END
  END imd_val_d_o[21]
  PIN imd_val_d_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 123.95 0.8 124.25 ;
    END
  END imd_val_d_o[22]
  PIN imd_val_d_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 138.91 0.8 139.21 ;
    END
  END imd_val_d_o[23]
  PIN imd_val_d_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  30.52 148.905 30.66 149.39 ;
    END
  END imd_val_d_o[24]
  PIN imd_val_d_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 144.35 0.8 144.65 ;
    END
  END imd_val_d_o[25]
  PIN imd_val_d_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  28.68 148.905 28.82 149.39 ;
    END
  END imd_val_d_o[26]
  PIN imd_val_d_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 134.83 0.8 135.13 ;
    END
  END imd_val_d_o[27]
  PIN imd_val_d_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  21.32 148.905 21.46 149.39 ;
    END
  END imd_val_d_o[28]
  PIN imd_val_d_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 99.47 0.8 99.77 ;
    END
  END imd_val_d_o[29]
  PIN imd_val_d_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 148.905 37.1 149.39 ;
    END
  END imd_val_d_o[2]
  PIN imd_val_d_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.04 148.905 13.18 149.39 ;
    END
  END imd_val_d_o[30]
  PIN imd_val_d_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  33.28 148.905 33.42 149.39 ;
    END
  END imd_val_d_o[31]
  PIN imd_val_d_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 145.71 0.8 146.01 ;
    END
  END imd_val_d_o[32]
  PIN imd_val_d_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 130.75 0.8 131.05 ;
    END
  END imd_val_d_o[33]
  PIN imd_val_d_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 102.19 0.8 102.49 ;
    END
  END imd_val_d_o[34]
  PIN imd_val_d_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 108.99 0.8 109.29 ;
    END
  END imd_val_d_o[35]
  PIN imd_val_d_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 132.11 0.8 132.41 ;
    END
  END imd_val_d_o[36]
  PIN imd_val_d_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 133.47 0.8 133.77 ;
    END
  END imd_val_d_o[37]
  PIN imd_val_d_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 148.905 20.54 149.39 ;
    END
  END imd_val_d_o[38]
  PIN imd_val_d_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 111.71 0.8 112.01 ;
    END
  END imd_val_d_o[39]
  PIN imd_val_d_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 148.905 27.9 149.39 ;
    END
  END imd_val_d_o[3]
  PIN imd_val_d_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 142.99 0.8 143.29 ;
    END
  END imd_val_d_o[40]
  PIN imd_val_d_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.04 148.905 36.18 149.39 ;
    END
  END imd_val_d_o[41]
  PIN imd_val_d_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  24.08 148.905 24.22 149.39 ;
    END
  END imd_val_d_o[42]
  PIN imd_val_d_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.92 148.905 26.06 149.39 ;
    END
  END imd_val_d_o[43]
  PIN imd_val_d_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  19.48 148.905 19.62 149.39 ;
    END
  END imd_val_d_o[44]
  PIN imd_val_d_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 125.31 0.8 125.61 ;
    END
  END imd_val_d_o[45]
  PIN imd_val_d_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  31.44 148.905 31.58 149.39 ;
    END
  END imd_val_d_o[46]
  PIN imd_val_d_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 95.39 0.8 95.69 ;
    END
  END imd_val_d_o[47]
  PIN imd_val_d_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 104.91 0.8 105.21 ;
    END
  END imd_val_d_o[48]
  PIN imd_val_d_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 121.23 0.8 121.53 ;
    END
  END imd_val_d_o[49]
  PIN imd_val_d_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  26.84 148.905 26.98 149.39 ;
    END
  END imd_val_d_o[4]
  PIN imd_val_d_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 113.07 0.8 113.37 ;
    END
  END imd_val_d_o[50]
  PIN imd_val_d_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 140.27 0.8 140.57 ;
    END
  END imd_val_d_o[51]
  PIN imd_val_d_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 119.87 0.8 120.17 ;
    END
  END imd_val_d_o[52]
  PIN imd_val_d_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 115.79 0.8 116.09 ;
    END
  END imd_val_d_o[53]
  PIN imd_val_d_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  8.44 148.905 8.58 149.39 ;
    END
  END imd_val_d_o[54]
  PIN imd_val_d_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 118.51 0.8 118.81 ;
    END
  END imd_val_d_o[55]
  PIN imd_val_d_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 110.35 0.8 110.65 ;
    END
  END imd_val_d_o[56]
  PIN imd_val_d_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.72 148.905 16.86 149.39 ;
    END
  END imd_val_d_o[57]
  PIN imd_val_d_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 148.905 29.74 149.39 ;
    END
  END imd_val_d_o[58]
  PIN imd_val_d_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  35.12 148.905 35.26 149.39 ;
    END
  END imd_val_d_o[59]
  PIN imd_val_d_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  23.16 148.905 23.3 149.39 ;
    END
  END imd_val_d_o[5]
  PIN imd_val_d_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 126.67 0.8 126.97 ;
    END
  END imd_val_d_o[60]
  PIN imd_val_d_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 96.75 0.8 97.05 ;
    END
  END imd_val_d_o[61]
  PIN imd_val_d_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  34.2 148.905 34.34 149.39 ;
    END
  END imd_val_d_o[62]
  PIN imd_val_d_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 107.63 0.8 107.93 ;
    END
  END imd_val_d_o[63]
  PIN imd_val_d_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 128.03 0.8 128.33 ;
    END
  END imd_val_d_o[6]
  PIN imd_val_d_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  22.24 148.905 22.38 149.39 ;
    END
  END imd_val_d_o[7]
  PIN imd_val_d_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 122.59 0.8 122.89 ;
    END
  END imd_val_d_o[8]
  PIN imd_val_d_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25 148.905 25.14 149.39 ;
    END
  END imd_val_d_o[9]
  PIN imd_val_q_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.72 0 16.86 0.485 ;
    END
  END imd_val_q_i[0]
  PIN imd_val_q_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  107.8 0 107.94 0.485 ;
    END
  END imd_val_q_i[10]
  PIN imd_val_q_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  4.76 0 4.9 0.485 ;
    END
  END imd_val_q_i[11]
  PIN imd_val_q_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.2 0 103.34 0.485 ;
    END
  END imd_val_q_i[12]
  PIN imd_val_q_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.04 0 13.18 0.485 ;
    END
  END imd_val_q_i[13]
  PIN imd_val_q_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  121.6 0 121.74 0.485 ;
    END
  END imd_val_q_i[14]
  PIN imd_val_q_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  110.56 0 110.7 0.485 ;
    END
  END imd_val_q_i[15]
  PIN imd_val_q_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  109.64 0 109.78 0.485 ;
    END
  END imd_val_q_i[16]
  PIN imd_val_q_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48 0 48.14 0.485 ;
    END
  END imd_val_q_i[17]
  PIN imd_val_q_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  106.88 0 107.02 0.485 ;
    END
  END imd_val_q_i[18]
  PIN imd_val_q_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.2 0 11.34 0.485 ;
    END
  END imd_val_q_i[19]
  PIN imd_val_q_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  5.68 0 5.82 0.485 ;
    END
  END imd_val_q_i[1]
  PIN imd_val_q_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  22.24 0 22.38 0.485 ;
    END
  END imd_val_q_i[20]
  PIN imd_val_q_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  116.08 0 116.22 0.485 ;
    END
  END imd_val_q_i[21]
  PIN imd_val_q_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  14.88 0 15.02 0.485 ;
    END
  END imd_val_q_i[22]
  PIN imd_val_q_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  28.68 0 28.82 0.485 ;
    END
  END imd_val_q_i[23]
  PIN imd_val_q_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  24.08 0 24.22 0.485 ;
    END
  END imd_val_q_i[24]
  PIN imd_val_q_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  114.24 0 114.38 0.485 ;
    END
  END imd_val_q_i[25]
  PIN imd_val_q_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 0 27.9 0.485 ;
    END
  END imd_val_q_i[26]
  PIN imd_val_q_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  19.48 0 19.62 0.485 ;
    END
  END imd_val_q_i[27]
  PIN imd_val_q_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 0 20.54 0.485 ;
    END
  END imd_val_q_i[28]
  PIN imd_val_q_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  21.32 0 21.46 0.485 ;
    END
  END imd_val_q_i[29]
  PIN imd_val_q_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.92 0 26.06 0.485 ;
    END
  END imd_val_q_i[2]
  PIN imd_val_q_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  113.32 0 113.46 0.485 ;
    END
  END imd_val_q_i[30]
  PIN imd_val_q_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 0 37.1 0.485 ;
    END
  END imd_val_q_i[31]
  PIN imd_val_q_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25 0 25.14 0.485 ;
    END
  END imd_val_q_i[32]
  PIN imd_val_q_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 0 29.74 0.485 ;
    END
  END imd_val_q_i[33]
  PIN imd_val_q_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  39.72 0 39.86 0.485 ;
    END
  END imd_val_q_i[34]
  PIN imd_val_q_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  37.88 0 38.02 0.485 ;
    END
  END imd_val_q_i[35]
  PIN imd_val_q_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  31.44 0 31.58 0.485 ;
    END
  END imd_val_q_i[36]
  PIN imd_val_q_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  30.52 0 30.66 0.485 ;
    END
  END imd_val_q_i[37]
  PIN imd_val_q_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  105.96 0 106.1 0.485 ;
    END
  END imd_val_q_i[38]
  PIN imd_val_q_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  32.36 0 32.5 0.485 ;
    END
  END imd_val_q_i[39]
  PIN imd_val_q_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  33.28 0 33.42 0.485 ;
    END
  END imd_val_q_i[3]
  PIN imd_val_q_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  117 0 117.14 0.485 ;
    END
  END imd_val_q_i[40]
  PIN imd_val_q_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.04 0 36.18 0.485 ;
    END
  END imd_val_q_i[41]
  PIN imd_val_q_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  49.84 0 49.98 0.485 ;
    END
  END imd_val_q_i[42]
  PIN imd_val_q_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  119.76 0 119.9 0.485 ;
    END
  END imd_val_q_i[43]
  PIN imd_val_q_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  117.92 0 118.06 0.485 ;
    END
  END imd_val_q_i[44]
  PIN imd_val_q_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  118.84 0 118.98 0.485 ;
    END
  END imd_val_q_i[45]
  PIN imd_val_q_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  40.64 0 40.78 0.485 ;
    END
  END imd_val_q_i[46]
  PIN imd_val_q_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  41.56 0 41.7 0.485 ;
    END
  END imd_val_q_i[47]
  PIN imd_val_q_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  42.48 0 42.62 0.485 ;
    END
  END imd_val_q_i[48]
  PIN imd_val_q_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  44.32 0 44.46 0.485 ;
    END
  END imd_val_q_i[49]
  PIN imd_val_q_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  45.24 0 45.38 0.485 ;
    END
  END imd_val_q_i[4]
  PIN imd_val_q_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.96 0 14.1 0.485 ;
    END
  END imd_val_q_i[50]
  PIN imd_val_q_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  47.08 0 47.22 0.485 ;
    END
  END imd_val_q_i[51]
  PIN imd_val_q_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  122.52 0 122.66 0.485 ;
    END
  END imd_val_q_i[52]
  PIN imd_val_q_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 0 9.5 0.485 ;
    END
  END imd_val_q_i[53]
  PIN imd_val_q_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  3.84 0 3.98 0.485 ;
    END
  END imd_val_q_i[54]
  PIN imd_val_q_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  23.16 0 23.3 0.485 ;
    END
  END imd_val_q_i[55]
  PIN imd_val_q_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  52.6 0 52.74 0.485 ;
    END
  END imd_val_q_i[56]
  PIN imd_val_q_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  6.6 0 6.74 0.485 ;
    END
  END imd_val_q_i[57]
  PIN imd_val_q_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2 0 2.14 0.485 ;
    END
  END imd_val_q_i[58]
  PIN imd_val_q_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  123.44 0 123.58 0.485 ;
    END
  END imd_val_q_i[59]
  PIN imd_val_q_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  15.8 0 15.94 0.485 ;
    END
  END imd_val_q_i[5]
  PIN imd_val_q_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  12.12 0 12.26 0.485 ;
    END
  END imd_val_q_i[60]
  PIN imd_val_q_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2.92 0 3.06 0.485 ;
    END
  END imd_val_q_i[61]
  PIN imd_val_q_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  17.64 0 17.78 0.485 ;
    END
  END imd_val_q_i[62]
  PIN imd_val_q_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  8.44 0 8.58 0.485 ;
    END
  END imd_val_q_i[63]
  PIN imd_val_q_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  10.28 0 10.42 0.485 ;
    END
  END imd_val_q_i[6]
  PIN imd_val_q_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 0 18.7 0.485 ;
    END
  END imd_val_q_i[7]
  PIN imd_val_q_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  120.68 0 120.82 0.485 ;
    END
  END imd_val_q_i[8]
  PIN imd_val_q_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.52 0 7.66 0.485 ;
    END
  END imd_val_q_i[9]
  PIN imd_val_we_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 141.63 0.8 141.93 ;
    END
  END imd_val_we_o[0]
  PIN imd_val_we_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 129.39 0.8 129.69 ;
    END
  END imd_val_we_o[1]
  PIN instr_first_cycle_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 104.91 149.39 105.21 ;
    END
  END instr_first_cycle_i
  PIN is_equal_result_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 80.43 149.39 80.73 ;
    END
  END is_equal_result_o
  PIN multdiv_operand_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 23.31 149.39 23.61 ;
    END
  END multdiv_operand_a_i[0]
  PIN multdiv_operand_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 49.15 0.8 49.45 ;
    END
  END multdiv_operand_a_i[10]
  PIN multdiv_operand_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 47.79 0.8 48.09 ;
    END
  END multdiv_operand_a_i[11]
  PIN multdiv_operand_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 45.07 0.8 45.37 ;
    END
  END multdiv_operand_a_i[12]
  PIN multdiv_operand_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 26.03 0.8 26.33 ;
    END
  END multdiv_operand_a_i[13]
  PIN multdiv_operand_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 43.71 0.8 44.01 ;
    END
  END multdiv_operand_a_i[14]
  PIN multdiv_operand_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 46.43 0.8 46.73 ;
    END
  END multdiv_operand_a_i[15]
  PIN multdiv_operand_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 9.71 0.8 10.01 ;
    END
  END multdiv_operand_a_i[16]
  PIN multdiv_operand_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 21.95 0.8 22.25 ;
    END
  END multdiv_operand_a_i[17]
  PIN multdiv_operand_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 11.07 0.8 11.37 ;
    END
  END multdiv_operand_a_i[18]
  PIN multdiv_operand_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 38.27 0.8 38.57 ;
    END
  END multdiv_operand_a_i[19]
  PIN multdiv_operand_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 40.99 149.39 41.29 ;
    END
  END multdiv_operand_a_i[1]
  PIN multdiv_operand_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 31.47 0.8 31.77 ;
    END
  END multdiv_operand_a_i[20]
  PIN multdiv_operand_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  35.12 0 35.26 0.485 ;
    END
  END multdiv_operand_a_i[21]
  PIN multdiv_operand_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48.92 0 49.06 0.485 ;
    END
  END multdiv_operand_a_i[22]
  PIN multdiv_operand_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  51.68 0 51.82 0.485 ;
    END
  END multdiv_operand_a_i[23]
  PIN multdiv_operand_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  56.28 0 56.42 0.485 ;
    END
  END multdiv_operand_a_i[24]
  PIN multdiv_operand_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.4 0 66.54 0.485 ;
    END
  END multdiv_operand_a_i[25]
  PIN multdiv_operand_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  89.4 0 89.54 0.485 ;
    END
  END multdiv_operand_a_i[26]
  PIN multdiv_operand_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  84.8 0 84.94 0.485 ;
    END
  END multdiv_operand_a_i[27]
  PIN multdiv_operand_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  105.04 0 105.18 0.485 ;
    END
  END multdiv_operand_a_i[28]
  PIN multdiv_operand_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.72 0 108.86 0.485 ;
    END
  END multdiv_operand_a_i[29]
  PIN multdiv_operand_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 64.11 149.39 64.41 ;
    END
  END multdiv_operand_a_i[2]
  PIN multdiv_operand_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 30.11 149.39 30.41 ;
    END
  END multdiv_operand_a_i[30]
  PIN multdiv_operand_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 28.75 149.39 29.05 ;
    END
  END multdiv_operand_a_i[31]
  PIN multdiv_operand_a_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 42.35 149.39 42.65 ;
    END
  END multdiv_operand_a_i[32]
  PIN multdiv_operand_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 54.59 149.39 54.89 ;
    END
  END multdiv_operand_a_i[3]
  PIN multdiv_operand_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 53.23 149.39 53.53 ;
    END
  END multdiv_operand_a_i[4]
  PIN multdiv_operand_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 38.27 149.39 38.57 ;
    END
  END multdiv_operand_a_i[5]
  PIN multdiv_operand_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 55.95 149.39 56.25 ;
    END
  END multdiv_operand_a_i[6]
  PIN multdiv_operand_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  81.12 0 81.26 0.485 ;
    END
  END multdiv_operand_a_i[7]
  PIN multdiv_operand_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  86.64 0 86.78 0.485 ;
    END
  END multdiv_operand_a_i[8]
  PIN multdiv_operand_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  67.32 0 67.46 0.485 ;
    END
  END multdiv_operand_a_i[9]
  PIN multdiv_operand_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 32.83 149.39 33.13 ;
    END
  END multdiv_operand_b_i[0]
  PIN multdiv_operand_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  58.12 0 58.26 0.485 ;
    END
  END multdiv_operand_b_i[10]
  PIN multdiv_operand_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 36.91 0.8 37.21 ;
    END
  END multdiv_operand_b_i[11]
  PIN multdiv_operand_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 34.19 0.8 34.49 ;
    END
  END multdiv_operand_b_i[12]
  PIN multdiv_operand_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 39.63 0.8 39.93 ;
    END
  END multdiv_operand_b_i[13]
  PIN multdiv_operand_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 55.95 0.8 56.25 ;
    END
  END multdiv_operand_b_i[14]
  PIN multdiv_operand_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 28.75 0.8 29.05 ;
    END
  END multdiv_operand_b_i[15]
  PIN multdiv_operand_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 16.51 0.8 16.81 ;
    END
  END multdiv_operand_b_i[16]
  PIN multdiv_operand_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 15.15 0.8 15.45 ;
    END
  END multdiv_operand_b_i[17]
  PIN multdiv_operand_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 40.99 0.8 41.29 ;
    END
  END multdiv_operand_b_i[18]
  PIN multdiv_operand_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 32.83 0.8 33.13 ;
    END
  END multdiv_operand_b_i[19]
  PIN multdiv_operand_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 60.03 149.39 60.33 ;
    END
  END multdiv_operand_b_i[1]
  PIN multdiv_operand_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 24.67 0.8 24.97 ;
    END
  END multdiv_operand_b_i[20]
  PIN multdiv_operand_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  38.8 0 38.94 0.485 ;
    END
  END multdiv_operand_b_i[21]
  PIN multdiv_operand_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  43.4 0 43.54 0.485 ;
    END
  END multdiv_operand_b_i[22]
  PIN multdiv_operand_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  50.76 0 50.9 0.485 ;
    END
  END multdiv_operand_b_i[23]
  PIN multdiv_operand_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  57.2 0 57.34 0.485 ;
    END
  END multdiv_operand_b_i[24]
  PIN multdiv_operand_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  68.24 0 68.38 0.485 ;
    END
  END multdiv_operand_b_i[25]
  PIN multdiv_operand_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.32 0 90.46 0.485 ;
    END
  END multdiv_operand_b_i[26]
  PIN multdiv_operand_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  83.88 0 84.02 0.485 ;
    END
  END multdiv_operand_b_i[27]
  PIN multdiv_operand_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  102.28 0 102.42 0.485 ;
    END
  END multdiv_operand_b_i[28]
  PIN multdiv_operand_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.4 0 112.54 0.485 ;
    END
  END multdiv_operand_b_i[29]
  PIN multdiv_operand_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 50.51 149.39 50.81 ;
    END
  END multdiv_operand_b_i[2]
  PIN multdiv_operand_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  115.16 0 115.3 0.485 ;
    END
  END multdiv_operand_b_i[30]
  PIN multdiv_operand_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 58.67 149.39 58.97 ;
    END
  END multdiv_operand_b_i[31]
  PIN multdiv_operand_b_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 57.31 149.39 57.61 ;
    END
  END multdiv_operand_b_i[32]
  PIN multdiv_operand_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 46.43 149.39 46.73 ;
    END
  END multdiv_operand_b_i[3]
  PIN multdiv_operand_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 49.15 149.39 49.45 ;
    END
  END multdiv_operand_b_i[4]
  PIN multdiv_operand_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 43.71 149.39 44.01 ;
    END
  END multdiv_operand_b_i[5]
  PIN multdiv_operand_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 39.63 149.39 39.93 ;
    END
  END multdiv_operand_b_i[6]
  PIN multdiv_operand_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.04 0 82.18 0.485 ;
    END
  END multdiv_operand_b_i[7]
  PIN multdiv_operand_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  87.56 0 87.7 0.485 ;
    END
  END multdiv_operand_b_i[8]
  PIN multdiv_operand_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  65.48 0 65.62 0.485 ;
    END
  END multdiv_operand_b_i[9]
  PIN multdiv_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  76.52 0 76.66 0.485 ;
    END
  END multdiv_sel_i
  PIN operand_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 113.07 149.39 113.37 ;
    END
  END operand_a_i[0]
  PIN operand_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 76.35 0.8 76.65 ;
    END
  END operand_a_i[10]
  PIN operand_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 74.99 0.8 75.29 ;
    END
  END operand_a_i[11]
  PIN operand_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  39.72 148.905 39.86 149.39 ;
    END
  END operand_a_i[12]
  PIN operand_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 87.23 0.8 87.53 ;
    END
  END operand_a_i[13]
  PIN operand_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 69.55 0.8 69.85 ;
    END
  END operand_a_i[14]
  PIN operand_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 103.55 0.8 103.85 ;
    END
  END operand_a_i[15]
  PIN operand_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 94.03 0.8 94.33 ;
    END
  END operand_a_i[16]
  PIN operand_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 77.71 0.8 78.01 ;
    END
  END operand_a_i[17]
  PIN operand_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 85.87 0.8 86.17 ;
    END
  END operand_a_i[18]
  PIN operand_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 100.83 0.8 101.13 ;
    END
  END operand_a_i[19]
  PIN operand_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 117.15 149.39 117.45 ;
    END
  END operand_a_i[1]
  PIN operand_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 80.43 0.8 80.73 ;
    END
  END operand_a_i[20]
  PIN operand_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 68.19 0.8 68.49 ;
    END
  END operand_a_i[21]
  PIN operand_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  49.84 148.905 49.98 149.39 ;
    END
  END operand_a_i[22]
  PIN operand_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.04 148.905 59.18 149.39 ;
    END
  END operand_a_i[23]
  PIN operand_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  77.44 148.905 77.58 149.39 ;
    END
  END operand_a_i[24]
  PIN operand_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  87.56 148.905 87.7 149.39 ;
    END
  END operand_a_i[25]
  PIN operand_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  98.6 148.905 98.74 149.39 ;
    END
  END operand_a_i[26]
  PIN operand_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.72 148.905 108.86 149.39 ;
    END
  END operand_a_i[27]
  PIN operand_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 123.95 149.39 124.25 ;
    END
  END operand_a_i[28]
  PIN operand_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 122.59 149.39 122.89 ;
    END
  END operand_a_i[29]
  PIN operand_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 125.31 149.39 125.61 ;
    END
  END operand_a_i[2]
  PIN operand_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 121.23 149.39 121.53 ;
    END
  END operand_a_i[30]
  PIN operand_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 115.79 149.39 116.09 ;
    END
  END operand_a_i[31]
  PIN operand_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 126.67 149.39 126.97 ;
    END
  END operand_a_i[3]
  PIN operand_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  106.88 148.905 107.02 149.39 ;
    END
  END operand_a_i[4]
  PIN operand_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.2 148.905 103.34 149.39 ;
    END
  END operand_a_i[5]
  PIN operand_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.32 148.905 90.46 149.39 ;
    END
  END operand_a_i[6]
  PIN operand_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  83.88 148.905 84.02 149.39 ;
    END
  END operand_a_i[7]
  PIN operand_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  65.48 148.905 65.62 149.39 ;
    END
  END operand_a_i[8]
  PIN operand_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  52.6 148.905 52.74 149.39 ;
    END
  END operand_a_i[9]
  PIN operand_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 114.43 149.39 114.73 ;
    END
  END operand_b_i[0]
  PIN operand_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 64.11 0.8 64.41 ;
    END
  END operand_b_i[10]
  PIN operand_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 57.31 0.8 57.61 ;
    END
  END operand_b_i[11]
  PIN operand_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 65.47 0.8 65.77 ;
    END
  END operand_b_i[12]
  PIN operand_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 61.39 0.8 61.69 ;
    END
  END operand_b_i[13]
  PIN operand_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 54.59 0.8 54.89 ;
    END
  END operand_b_i[14]
  PIN operand_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 27.39 0.8 27.69 ;
    END
  END operand_b_i[15]
  PIN operand_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 51.87 0.8 52.17 ;
    END
  END operand_b_i[16]
  PIN operand_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 58.67 0.8 58.97 ;
    END
  END operand_b_i[17]
  PIN operand_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 62.75 0.8 63.05 ;
    END
  END operand_b_i[18]
  PIN operand_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 60.03 0.8 60.33 ;
    END
  END operand_b_i[19]
  PIN operand_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 103.55 149.39 103.85 ;
    END
  END operand_b_i[1]
  PIN operand_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 20.59 0.8 20.89 ;
    END
  END operand_b_i[20]
  PIN operand_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 42.35 0.8 42.65 ;
    END
  END operand_b_i[21]
  PIN operand_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 50.51 0.8 50.81 ;
    END
  END operand_b_i[22]
  PIN operand_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 17.87 0.8 18.17 ;
    END
  END operand_b_i[23]
  PIN operand_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 23.31 0.8 23.61 ;
    END
  END operand_b_i[24]
  PIN operand_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  88.48 0 88.62 0.485 ;
    END
  END operand_b_i[25]
  PIN operand_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.96 0 83.1 0.485 ;
    END
  END operand_b_i[26]
  PIN operand_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 98.11 149.39 98.41 ;
    END
  END operand_b_i[27]
  PIN operand_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 31.47 149.39 31.77 ;
    END
  END operand_b_i[28]
  PIN operand_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 27.39 149.39 27.69 ;
    END
  END operand_b_i[29]
  PIN operand_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 111.71 149.39 112.01 ;
    END
  END operand_b_i[2]
  PIN operand_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 84.51 149.39 84.81 ;
    END
  END operand_b_i[30]
  PIN operand_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 77.71 149.39 78.01 ;
    END
  END operand_b_i[31]
  PIN operand_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 102.19 149.39 102.49 ;
    END
  END operand_b_i[3]
  PIN operand_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 100.83 149.39 101.13 ;
    END
  END operand_b_i[4]
  PIN operand_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 95.39 149.39 95.69 ;
    END
  END operand_b_i[5]
  PIN operand_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  78.36 0 78.5 0.485 ;
    END
  END operand_b_i[6]
  PIN operand_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 76.35 149.39 76.65 ;
    END
  END operand_b_i[7]
  PIN operand_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  61.8 0 61.94 0.485 ;
    END
  END operand_b_i[8]
  PIN operand_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 53.23 0.8 53.53 ;
    END
  END operand_b_i[9]
  PIN operator_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 118.51 149.39 118.81 ;
    END
  END operator_i[0]
  PIN operator_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 119.87 149.39 120.17 ;
    END
  END operator_i[1]
  PIN operator_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 107.63 149.39 107.93 ;
    END
  END operator_i[2]
  PIN operator_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 106.27 149.39 106.57 ;
    END
  END operator_i[3]
  PIN operator_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 110.35 149.39 110.65 ;
    END
  END operator_i[4]
  PIN operator_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 108.99 149.39 109.29 ;
    END
  END operator_i[5]
  PIN result_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 91.31 149.39 91.61 ;
    END
  END result_o[0]
  PIN result_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71.92 148.905 72.06 149.39 ;
    END
  END result_o[10]
  PIN result_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 79.07 0.8 79.37 ;
    END
  END result_o[11]
  PIN result_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  68.24 148.905 68.38 149.39 ;
    END
  END result_o[12]
  PIN result_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  61.8 148.905 61.94 149.39 ;
    END
  END result_o[13]
  PIN result_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 72.27 0.8 72.57 ;
    END
  END result_o[14]
  PIN result_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  60.88 148.905 61.02 149.39 ;
    END
  END result_o[15]
  PIN result_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.96 148.905 60.1 149.39 ;
    END
  END result_o[16]
  PIN result_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 73.63 0.8 73.93 ;
    END
  END result_o[17]
  PIN result_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  62.72 148.905 62.86 149.39 ;
    END
  END result_o[18]
  PIN result_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  67.32 148.905 67.46 149.39 ;
    END
  END result_o[19]
  PIN result_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 81.79 149.39 82.09 ;
    END
  END result_o[1]
  PIN result_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 81.79 0.8 82.09 ;
    END
  END result_o[20]
  PIN result_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 148.905 73.9 149.39 ;
    END
  END result_o[21]
  PIN result_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  72.84 148.905 72.98 149.39 ;
    END
  END result_o[22]
  PIN result_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71.92 0 72.06 0.485 ;
    END
  END result_o[23]
  PIN result_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 88.59 149.39 88.89 ;
    END
  END result_o[24]
  PIN result_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 74.99 149.39 75.29 ;
    END
  END result_o[25]
  PIN result_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 69.55 149.39 69.85 ;
    END
  END result_o[26]
  PIN result_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  88.48 148.905 88.62 149.39 ;
    END
  END result_o[27]
  PIN result_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 66.83 149.39 67.13 ;
    END
  END result_o[28]
  PIN result_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 68.19 149.39 68.49 ;
    END
  END result_o[29]
  PIN result_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 70.91 149.39 71.21 ;
    END
  END result_o[2]
  PIN result_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 85.87 149.39 86.17 ;
    END
  END result_o[30]
  PIN result_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 94.03 149.39 94.33 ;
    END
  END result_o[31]
  PIN result_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 73.63 149.39 73.93 ;
    END
  END result_o[3]
  PIN result_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  89.4 148.905 89.54 149.39 ;
    END
  END result_o[4]
  PIN result_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 96.75 149.39 97.05 ;
    END
  END result_o[5]
  PIN result_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 72.27 149.39 72.57 ;
    END
  END result_o[6]
  PIN result_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  148.59 89.95 149.39 90.25 ;
    END
  END result_o[7]
  PIN result_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 70.91 0.8 71.21 ;
    END
  END result_o[8]
  PIN result_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  74.68 148.905 74.82 149.39 ;
    END
  END result_o[9]
  OBS
    LAYER nwell ;
     RECT  0 0 149.39 149.39 ;
    LAYER pwell ;
     RECT  0 0 149.39 149.39 ;
    LAYER li1 ;
     RECT  0 0 149.39 149.39 ;
    LAYER met1 ;
     RECT  0 0 149.39 149.39 ;
    LAYER met2 ;
     RECT  0 0 149.39 149.39 ;
    LAYER met3 ;
     RECT  0 0 149.39 149.39 ;
    LAYER met4 ;
     RECT  0 0 149.39 149.39 ;
    LAYER met5 ;
     RECT  0 0 149.39 149.39 ;
  END
END ibex_alu
END LIBRARY
