module fakeram7_256x32 (ce_in,
    clk,
    we_in,
    addr_in,
    rd_out,
    wd_in);
 input ce_in;
 input clk;
 input we_in;
 input [7:0] addr_in;
 output [31:0] rd_out;
 input [31:0] wd_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;

 INVx1_ASAP7_75t_R _238_ (.A(_063_),
    .Y(_128_));
 AND2x6_ASAP7_75t_R _239_ (.A(net1),
    .B(net2),
    .Y(_129_));
 BUFx4f_ASAP7_75t_R _240_ (.A(_129_),
    .Y(_130_));
 AND2x2_ASAP7_75t_R _241_ (.A(_128_),
    .B(_130_),
    .Y(_000_));
 INVx1_ASAP7_75t_R _242_ (.A(_052_),
    .Y(_131_));
 AND2x2_ASAP7_75t_R _243_ (.A(_131_),
    .B(_130_),
    .Y(_011_));
 INVx1_ASAP7_75t_R _244_ (.A(_041_),
    .Y(_132_));
 AND2x2_ASAP7_75t_R _245_ (.A(_132_),
    .B(_130_),
    .Y(_022_));
 INVx1_ASAP7_75t_R _246_ (.A(_038_),
    .Y(_133_));
 AND2x2_ASAP7_75t_R _247_ (.A(_133_),
    .B(_130_),
    .Y(_025_));
 INVx1_ASAP7_75t_R _248_ (.A(_037_),
    .Y(_134_));
 AND2x2_ASAP7_75t_R _249_ (.A(_134_),
    .B(_130_),
    .Y(_026_));
 INVx1_ASAP7_75t_R _250_ (.A(_036_),
    .Y(_135_));
 AND2x2_ASAP7_75t_R _251_ (.A(_135_),
    .B(_130_),
    .Y(_027_));
 INVx1_ASAP7_75t_R _252_ (.A(_035_),
    .Y(_136_));
 AND2x2_ASAP7_75t_R _253_ (.A(_136_),
    .B(_130_),
    .Y(_028_));
 INVx1_ASAP7_75t_R _254_ (.A(_034_),
    .Y(_137_));
 AND2x2_ASAP7_75t_R _255_ (.A(_137_),
    .B(_130_),
    .Y(_029_));
 INVx1_ASAP7_75t_R _256_ (.A(_033_),
    .Y(_138_));
 AND2x2_ASAP7_75t_R _257_ (.A(_138_),
    .B(_130_),
    .Y(_030_));
 INVx1_ASAP7_75t_R _258_ (.A(_064_),
    .Y(_139_));
 AND2x2_ASAP7_75t_R _259_ (.A(_139_),
    .B(_130_),
    .Y(_031_));
 INVx1_ASAP7_75t_R _260_ (.A(_062_),
    .Y(_140_));
 BUFx3_ASAP7_75t_R _261_ (.A(_129_),
    .Y(_141_));
 AND2x2_ASAP7_75t_R _262_ (.A(_140_),
    .B(_141_),
    .Y(_001_));
 INVx1_ASAP7_75t_R _263_ (.A(_061_),
    .Y(_142_));
 AND2x2_ASAP7_75t_R _264_ (.A(_142_),
    .B(_141_),
    .Y(_002_));
 INVx1_ASAP7_75t_R _265_ (.A(_060_),
    .Y(_143_));
 AND2x2_ASAP7_75t_R _266_ (.A(_143_),
    .B(_141_),
    .Y(_003_));
 INVx1_ASAP7_75t_R _267_ (.A(_059_),
    .Y(_144_));
 AND2x2_ASAP7_75t_R _268_ (.A(_144_),
    .B(_141_),
    .Y(_004_));
 INVx1_ASAP7_75t_R _269_ (.A(_058_),
    .Y(_145_));
 AND2x2_ASAP7_75t_R _270_ (.A(_145_),
    .B(_141_),
    .Y(_005_));
 INVx1_ASAP7_75t_R _271_ (.A(_057_),
    .Y(_146_));
 AND2x2_ASAP7_75t_R _272_ (.A(_146_),
    .B(_141_),
    .Y(_006_));
 INVx1_ASAP7_75t_R _273_ (.A(_056_),
    .Y(_147_));
 AND2x2_ASAP7_75t_R _274_ (.A(_147_),
    .B(_141_),
    .Y(_007_));
 INVx1_ASAP7_75t_R _275_ (.A(_055_),
    .Y(_148_));
 AND2x2_ASAP7_75t_R _276_ (.A(_148_),
    .B(_141_),
    .Y(_008_));
 INVx1_ASAP7_75t_R _277_ (.A(_054_),
    .Y(_149_));
 AND2x2_ASAP7_75t_R _278_ (.A(_149_),
    .B(_141_),
    .Y(_009_));
 INVx1_ASAP7_75t_R _279_ (.A(_053_),
    .Y(_150_));
 AND2x2_ASAP7_75t_R _280_ (.A(_150_),
    .B(_141_),
    .Y(_010_));
 INVx1_ASAP7_75t_R _281_ (.A(_051_),
    .Y(_151_));
 BUFx3_ASAP7_75t_R _282_ (.A(_129_),
    .Y(_152_));
 AND2x2_ASAP7_75t_R _283_ (.A(_151_),
    .B(_152_),
    .Y(_012_));
 INVx1_ASAP7_75t_R _284_ (.A(_050_),
    .Y(_153_));
 AND2x2_ASAP7_75t_R _285_ (.A(_153_),
    .B(_152_),
    .Y(_013_));
 INVx1_ASAP7_75t_R _286_ (.A(_049_),
    .Y(_154_));
 AND2x2_ASAP7_75t_R _287_ (.A(_154_),
    .B(_152_),
    .Y(_014_));
 INVx1_ASAP7_75t_R _288_ (.A(_048_),
    .Y(_155_));
 AND2x2_ASAP7_75t_R _289_ (.A(_155_),
    .B(_152_),
    .Y(_015_));
 INVx1_ASAP7_75t_R _290_ (.A(_047_),
    .Y(_156_));
 AND2x2_ASAP7_75t_R _291_ (.A(_156_),
    .B(_152_),
    .Y(_016_));
 INVx1_ASAP7_75t_R _292_ (.A(_046_),
    .Y(_157_));
 AND2x2_ASAP7_75t_R _293_ (.A(_157_),
    .B(_152_),
    .Y(_017_));
 INVx1_ASAP7_75t_R _294_ (.A(_045_),
    .Y(_158_));
 AND2x2_ASAP7_75t_R _295_ (.A(_158_),
    .B(_152_),
    .Y(_018_));
 INVx1_ASAP7_75t_R _296_ (.A(_044_),
    .Y(_159_));
 AND2x2_ASAP7_75t_R _297_ (.A(_159_),
    .B(_152_),
    .Y(_019_));
 INVx1_ASAP7_75t_R _298_ (.A(_043_),
    .Y(_160_));
 AND2x2_ASAP7_75t_R _299_ (.A(_160_),
    .B(_152_),
    .Y(_020_));
 INVx1_ASAP7_75t_R _300_ (.A(_042_),
    .Y(_161_));
 AND2x2_ASAP7_75t_R _301_ (.A(_161_),
    .B(_152_),
    .Y(_021_));
 INVx1_ASAP7_75t_R _302_ (.A(_040_),
    .Y(_162_));
 BUFx4f_ASAP7_75t_R _303_ (.A(_129_),
    .Y(_163_));
 AND2x2_ASAP7_75t_R _304_ (.A(_162_),
    .B(_163_),
    .Y(_023_));
 INVx1_ASAP7_75t_R _305_ (.A(_039_),
    .Y(_164_));
 AND2x2_ASAP7_75t_R _306_ (.A(_164_),
    .B(_163_),
    .Y(_024_));
 INVx1_ASAP7_75t_R _307_ (.A(_032_),
    .Y(net66));
 INVx1_ASAP7_75t_R _308_ (.A(_065_),
    .Y(net35));
 INVx1_ASAP7_75t_R _309_ (.A(_066_),
    .Y(net36));
 INVx1_ASAP7_75t_R _310_ (.A(_067_),
    .Y(net37));
 INVx1_ASAP7_75t_R _311_ (.A(_068_),
    .Y(net38));
 INVx1_ASAP7_75t_R _312_ (.A(_069_),
    .Y(net39));
 INVx1_ASAP7_75t_R _313_ (.A(_070_),
    .Y(net40));
 INVx1_ASAP7_75t_R _314_ (.A(_071_),
    .Y(net41));
 INVx1_ASAP7_75t_R _315_ (.A(_072_),
    .Y(net42));
 INVx1_ASAP7_75t_R _316_ (.A(_073_),
    .Y(net43));
 INVx1_ASAP7_75t_R _317_ (.A(_074_),
    .Y(net44));
 INVx1_ASAP7_75t_R _318_ (.A(_075_),
    .Y(net45));
 INVx1_ASAP7_75t_R _319_ (.A(_076_),
    .Y(net46));
 INVx1_ASAP7_75t_R _320_ (.A(_077_),
    .Y(net47));
 INVx1_ASAP7_75t_R _321_ (.A(_078_),
    .Y(net48));
 INVx1_ASAP7_75t_R _322_ (.A(_079_),
    .Y(net49));
 INVx1_ASAP7_75t_R _323_ (.A(_080_),
    .Y(net50));
 INVx1_ASAP7_75t_R _324_ (.A(_081_),
    .Y(net51));
 INVx1_ASAP7_75t_R _325_ (.A(_082_),
    .Y(net52));
 INVx1_ASAP7_75t_R _326_ (.A(_083_),
    .Y(net53));
 INVx1_ASAP7_75t_R _327_ (.A(_084_),
    .Y(net54));
 INVx1_ASAP7_75t_R _328_ (.A(_085_),
    .Y(net55));
 INVx1_ASAP7_75t_R _329_ (.A(_086_),
    .Y(net56));
 INVx1_ASAP7_75t_R _330_ (.A(_087_),
    .Y(net57));
 INVx1_ASAP7_75t_R _331_ (.A(_088_),
    .Y(net58));
 INVx1_ASAP7_75t_R _332_ (.A(_089_),
    .Y(net59));
 INVx1_ASAP7_75t_R _333_ (.A(_090_),
    .Y(net60));
 INVx1_ASAP7_75t_R _334_ (.A(_091_),
    .Y(net61));
 INVx1_ASAP7_75t_R _335_ (.A(_092_),
    .Y(net62));
 INVx1_ASAP7_75t_R _336_ (.A(_093_),
    .Y(net63));
 INVx1_ASAP7_75t_R _337_ (.A(_094_),
    .Y(net64));
 INVx1_ASAP7_75t_R _338_ (.A(_095_),
    .Y(net65));
 BUFx12f_ASAP7_75t_R _339_ (.A(ce_in),
    .Y(_165_));
 BUFx6f_ASAP7_75t_R _340_ (.A(_165_),
    .Y(_166_));
 AND2x2_ASAP7_75t_R _341_ (.A(net3),
    .B(_166_),
    .Y(_167_));
 BUFx6f_ASAP7_75t_R _342_ (.A(_165_),
    .Y(_168_));
 NOR2x1_ASAP7_75t_R _343_ (.A(_063_),
    .B(_168_),
    .Y(_169_));
 AO211x2_ASAP7_75t_R _344_ (.A1(_128_),
    .A2(_163_),
    .B(_167_),
    .C(_169_),
    .Y(_096_));
 AND2x2_ASAP7_75t_R _345_ (.A(net4),
    .B(_166_),
    .Y(_170_));
 NOR2x1_ASAP7_75t_R _346_ (.A(_062_),
    .B(_168_),
    .Y(_171_));
 AO211x2_ASAP7_75t_R _347_ (.A1(_140_),
    .A2(_163_),
    .B(_170_),
    .C(_171_),
    .Y(_097_));
 AND2x2_ASAP7_75t_R _348_ (.A(net5),
    .B(_166_),
    .Y(_172_));
 NOR2x1_ASAP7_75t_R _349_ (.A(_061_),
    .B(_168_),
    .Y(_173_));
 AO211x2_ASAP7_75t_R _350_ (.A1(_142_),
    .A2(_163_),
    .B(_172_),
    .C(_173_),
    .Y(_098_));
 AND2x2_ASAP7_75t_R _351_ (.A(net6),
    .B(_166_),
    .Y(_174_));
 NOR2x1_ASAP7_75t_R _352_ (.A(_060_),
    .B(_168_),
    .Y(_175_));
 AO211x2_ASAP7_75t_R _353_ (.A1(_143_),
    .A2(_163_),
    .B(_174_),
    .C(_175_),
    .Y(_099_));
 AND2x2_ASAP7_75t_R _354_ (.A(net7),
    .B(_166_),
    .Y(_176_));
 NOR2x1_ASAP7_75t_R _355_ (.A(_059_),
    .B(_168_),
    .Y(_177_));
 AO211x2_ASAP7_75t_R _356_ (.A1(_144_),
    .A2(_163_),
    .B(_176_),
    .C(_177_),
    .Y(_100_));
 AND2x2_ASAP7_75t_R _357_ (.A(net8),
    .B(_166_),
    .Y(_178_));
 NOR2x1_ASAP7_75t_R _358_ (.A(_058_),
    .B(_168_),
    .Y(_179_));
 AO211x2_ASAP7_75t_R _359_ (.A1(_145_),
    .A2(_163_),
    .B(_178_),
    .C(_179_),
    .Y(_101_));
 AND2x2_ASAP7_75t_R _360_ (.A(net9),
    .B(_166_),
    .Y(_180_));
 NOR2x1_ASAP7_75t_R _361_ (.A(_057_),
    .B(_168_),
    .Y(_181_));
 AO211x2_ASAP7_75t_R _362_ (.A1(_146_),
    .A2(_163_),
    .B(_180_),
    .C(_181_),
    .Y(_102_));
 AND2x2_ASAP7_75t_R _363_ (.A(net10),
    .B(_166_),
    .Y(_182_));
 NOR2x1_ASAP7_75t_R _364_ (.A(_056_),
    .B(_168_),
    .Y(_183_));
 AO211x2_ASAP7_75t_R _365_ (.A1(_147_),
    .A2(_163_),
    .B(_182_),
    .C(_183_),
    .Y(_103_));
 BUFx6f_ASAP7_75t_R _366_ (.A(_129_),
    .Y(_184_));
 BUFx6f_ASAP7_75t_R _367_ (.A(_165_),
    .Y(_185_));
 AND2x2_ASAP7_75t_R _368_ (.A(net11),
    .B(_185_),
    .Y(_186_));
 NOR2x1_ASAP7_75t_R _369_ (.A(_055_),
    .B(_168_),
    .Y(_187_));
 AO211x2_ASAP7_75t_R _370_ (.A1(_148_),
    .A2(_184_),
    .B(_186_),
    .C(_187_),
    .Y(_104_));
 AND2x2_ASAP7_75t_R _371_ (.A(net12),
    .B(_185_),
    .Y(_188_));
 NOR2x1_ASAP7_75t_R _372_ (.A(_054_),
    .B(_168_),
    .Y(_189_));
 AO211x2_ASAP7_75t_R _373_ (.A1(_149_),
    .A2(_184_),
    .B(_188_),
    .C(_189_),
    .Y(_105_));
 AND2x2_ASAP7_75t_R _374_ (.A(net13),
    .B(_185_),
    .Y(_190_));
 BUFx6f_ASAP7_75t_R _375_ (.A(_165_),
    .Y(_191_));
 NOR2x1_ASAP7_75t_R _376_ (.A(_053_),
    .B(_191_),
    .Y(_192_));
 AO211x2_ASAP7_75t_R _377_ (.A1(_150_),
    .A2(_184_),
    .B(_190_),
    .C(_192_),
    .Y(_106_));
 AND2x2_ASAP7_75t_R _378_ (.A(net14),
    .B(_185_),
    .Y(_193_));
 NOR2x1_ASAP7_75t_R _379_ (.A(_052_),
    .B(_191_),
    .Y(_194_));
 AO211x2_ASAP7_75t_R _380_ (.A1(_131_),
    .A2(_184_),
    .B(_193_),
    .C(_194_),
    .Y(_107_));
 AND2x2_ASAP7_75t_R _381_ (.A(net15),
    .B(_185_),
    .Y(_195_));
 NOR2x1_ASAP7_75t_R _382_ (.A(_051_),
    .B(_191_),
    .Y(_196_));
 AO211x2_ASAP7_75t_R _383_ (.A1(_151_),
    .A2(_184_),
    .B(_195_),
    .C(_196_),
    .Y(_108_));
 AND2x2_ASAP7_75t_R _384_ (.A(net16),
    .B(_185_),
    .Y(_197_));
 NOR2x1_ASAP7_75t_R _385_ (.A(_050_),
    .B(_191_),
    .Y(_198_));
 AO211x2_ASAP7_75t_R _386_ (.A1(_153_),
    .A2(_184_),
    .B(_197_),
    .C(_198_),
    .Y(_109_));
 AND2x2_ASAP7_75t_R _387_ (.A(net17),
    .B(_185_),
    .Y(_199_));
 NOR2x1_ASAP7_75t_R _388_ (.A(_049_),
    .B(_191_),
    .Y(_200_));
 AO211x2_ASAP7_75t_R _389_ (.A1(_154_),
    .A2(_184_),
    .B(_199_),
    .C(_200_),
    .Y(_110_));
 AND2x2_ASAP7_75t_R _390_ (.A(net18),
    .B(_185_),
    .Y(_201_));
 NOR2x1_ASAP7_75t_R _391_ (.A(_048_),
    .B(_191_),
    .Y(_202_));
 AO211x2_ASAP7_75t_R _392_ (.A1(_155_),
    .A2(_184_),
    .B(_201_),
    .C(_202_),
    .Y(_111_));
 AND2x2_ASAP7_75t_R _393_ (.A(net19),
    .B(_185_),
    .Y(_203_));
 NOR2x1_ASAP7_75t_R _394_ (.A(_047_),
    .B(_191_),
    .Y(_204_));
 AO211x2_ASAP7_75t_R _395_ (.A1(_156_),
    .A2(_184_),
    .B(_203_),
    .C(_204_),
    .Y(_112_));
 AND2x2_ASAP7_75t_R _396_ (.A(net20),
    .B(_185_),
    .Y(_205_));
 NOR2x1_ASAP7_75t_R _397_ (.A(_046_),
    .B(_191_),
    .Y(_206_));
 AO211x2_ASAP7_75t_R _398_ (.A1(_157_),
    .A2(_184_),
    .B(_205_),
    .C(_206_),
    .Y(_113_));
 BUFx6f_ASAP7_75t_R _399_ (.A(_129_),
    .Y(_207_));
 BUFx6f_ASAP7_75t_R _400_ (.A(_165_),
    .Y(_208_));
 AND2x2_ASAP7_75t_R _401_ (.A(net21),
    .B(_208_),
    .Y(_209_));
 NOR2x1_ASAP7_75t_R _402_ (.A(_045_),
    .B(_191_),
    .Y(_210_));
 AO211x2_ASAP7_75t_R _403_ (.A1(_158_),
    .A2(_207_),
    .B(_209_),
    .C(_210_),
    .Y(_114_));
 AND2x2_ASAP7_75t_R _404_ (.A(net22),
    .B(_208_),
    .Y(_211_));
 NOR2x1_ASAP7_75t_R _405_ (.A(_044_),
    .B(_191_),
    .Y(_212_));
 AO211x2_ASAP7_75t_R _406_ (.A1(_159_),
    .A2(_207_),
    .B(_211_),
    .C(_212_),
    .Y(_115_));
 AND2x2_ASAP7_75t_R _407_ (.A(net23),
    .B(_208_),
    .Y(_213_));
 BUFx6f_ASAP7_75t_R _408_ (.A(_165_),
    .Y(_214_));
 NOR2x1_ASAP7_75t_R _409_ (.A(_043_),
    .B(_214_),
    .Y(_215_));
 AO211x2_ASAP7_75t_R _410_ (.A1(_160_),
    .A2(_207_),
    .B(_213_),
    .C(_215_),
    .Y(_116_));
 AND2x2_ASAP7_75t_R _411_ (.A(net24),
    .B(_208_),
    .Y(_216_));
 NOR2x1_ASAP7_75t_R _412_ (.A(_042_),
    .B(_214_),
    .Y(_217_));
 AO211x2_ASAP7_75t_R _413_ (.A1(_161_),
    .A2(_207_),
    .B(_216_),
    .C(_217_),
    .Y(_117_));
 AND2x2_ASAP7_75t_R _414_ (.A(net25),
    .B(_208_),
    .Y(_218_));
 NOR2x1_ASAP7_75t_R _415_ (.A(_041_),
    .B(_214_),
    .Y(_219_));
 AO211x2_ASAP7_75t_R _416_ (.A1(_132_),
    .A2(_207_),
    .B(_218_),
    .C(_219_),
    .Y(_118_));
 AND2x2_ASAP7_75t_R _417_ (.A(net26),
    .B(_208_),
    .Y(_220_));
 NOR2x1_ASAP7_75t_R _418_ (.A(_040_),
    .B(_214_),
    .Y(_221_));
 AO211x2_ASAP7_75t_R _419_ (.A1(_162_),
    .A2(_207_),
    .B(_220_),
    .C(_221_),
    .Y(_119_));
 AND2x2_ASAP7_75t_R _420_ (.A(net27),
    .B(_208_),
    .Y(_222_));
 NOR2x1_ASAP7_75t_R _421_ (.A(_039_),
    .B(_214_),
    .Y(_223_));
 AO211x2_ASAP7_75t_R _422_ (.A1(_164_),
    .A2(_207_),
    .B(_222_),
    .C(_223_),
    .Y(_120_));
 AND2x2_ASAP7_75t_R _423_ (.A(net28),
    .B(_208_),
    .Y(_224_));
 NOR2x1_ASAP7_75t_R _424_ (.A(_038_),
    .B(_214_),
    .Y(_225_));
 AO211x2_ASAP7_75t_R _425_ (.A1(_133_),
    .A2(_207_),
    .B(_224_),
    .C(_225_),
    .Y(_121_));
 AND2x2_ASAP7_75t_R _426_ (.A(net29),
    .B(_208_),
    .Y(_226_));
 NOR2x1_ASAP7_75t_R _427_ (.A(_037_),
    .B(_214_),
    .Y(_227_));
 AO211x2_ASAP7_75t_R _428_ (.A1(_134_),
    .A2(_207_),
    .B(_226_),
    .C(_227_),
    .Y(_122_));
 AND2x2_ASAP7_75t_R _429_ (.A(net30),
    .B(_208_),
    .Y(_228_));
 NOR2x1_ASAP7_75t_R _430_ (.A(_036_),
    .B(_214_),
    .Y(_229_));
 AO211x2_ASAP7_75t_R _431_ (.A1(_135_),
    .A2(_207_),
    .B(_228_),
    .C(_229_),
    .Y(_123_));
 AND2x2_ASAP7_75t_R _432_ (.A(net31),
    .B(_165_),
    .Y(_230_));
 NOR2x1_ASAP7_75t_R _433_ (.A(_035_),
    .B(_214_),
    .Y(_231_));
 AO211x2_ASAP7_75t_R _434_ (.A1(_136_),
    .A2(_129_),
    .B(_230_),
    .C(_231_),
    .Y(_124_));
 AND2x2_ASAP7_75t_R _435_ (.A(net32),
    .B(_165_),
    .Y(_232_));
 NOR2x1_ASAP7_75t_R _436_ (.A(_034_),
    .B(_214_),
    .Y(_233_));
 AO211x2_ASAP7_75t_R _437_ (.A1(_137_),
    .A2(_129_),
    .B(_232_),
    .C(_233_),
    .Y(_125_));
 AND2x2_ASAP7_75t_R _438_ (.A(net33),
    .B(_165_),
    .Y(_234_));
 NOR2x1_ASAP7_75t_R _439_ (.A(_033_),
    .B(_166_),
    .Y(_235_));
 AO211x2_ASAP7_75t_R _440_ (.A1(_138_),
    .A2(_129_),
    .B(_234_),
    .C(_235_),
    .Y(_126_));
 AND2x2_ASAP7_75t_R _441_ (.A(net34),
    .B(_165_),
    .Y(_236_));
 NOR2x1_ASAP7_75t_R _442_ (.A(_064_),
    .B(_166_),
    .Y(_237_));
 AO211x2_ASAP7_75t_R _443_ (.A1(_139_),
    .A2(_129_),
    .B(_236_),
    .C(_237_),
    .Y(_127_));
 DFFHQNx2_ASAP7_75t_R \mem[3][0]$_DFFE_PP_  (.CLK(clknet_3_3_0_clk),
    .D(_096_),
    .QN(_063_));
 DFFHQNx2_ASAP7_75t_R \mem[3][10]$_DFFE_PP_  (.CLK(clknet_3_2_0_clk),
    .D(_097_),
    .QN(_062_));
 DFFHQNx2_ASAP7_75t_R \mem[3][11]$_DFFE_PP_  (.CLK(clknet_3_0_0_clk),
    .D(_098_),
    .QN(_061_));
 DFFHQNx2_ASAP7_75t_R \mem[3][12]$_DFFE_PP_  (.CLK(clknet_3_2_0_clk),
    .D(_099_),
    .QN(_060_));
 DFFHQNx2_ASAP7_75t_R \mem[3][13]$_DFFE_PP_  (.CLK(clknet_3_2_0_clk),
    .D(_100_),
    .QN(_059_));
 DFFHQNx2_ASAP7_75t_R \mem[3][14]$_DFFE_PP_  (.CLK(clknet_3_0_0_clk),
    .D(_101_),
    .QN(_058_));
 DFFHQNx2_ASAP7_75t_R \mem[3][15]$_DFFE_PP_  (.CLK(clknet_3_2_0_clk),
    .D(_102_),
    .QN(_057_));
 DFFHQNx2_ASAP7_75t_R \mem[3][16]$_DFFE_PP_  (.CLK(clknet_3_0_0_clk),
    .D(_103_),
    .QN(_056_));
 DFFHQNx2_ASAP7_75t_R \mem[3][17]$_DFFE_PP_  (.CLK(clknet_3_1_0_clk),
    .D(_104_),
    .QN(_055_));
 DFFHQNx2_ASAP7_75t_R \mem[3][18]$_DFFE_PP_  (.CLK(clknet_3_3_0_clk),
    .D(_105_),
    .QN(_054_));
 DFFHQNx2_ASAP7_75t_R \mem[3][19]$_DFFE_PP_  (.CLK(clknet_3_3_0_clk),
    .D(_106_),
    .QN(_053_));
 DFFHQNx2_ASAP7_75t_R \mem[3][1]$_DFFE_PP_  (.CLK(clknet_3_3_0_clk),
    .D(_107_),
    .QN(_052_));
 DFFHQNx2_ASAP7_75t_R \mem[3][20]$_DFFE_PP_  (.CLK(clknet_3_6_0_clk),
    .D(_108_),
    .QN(_051_));
 DFFHQNx2_ASAP7_75t_R \mem[3][21]$_DFFE_PP_  (.CLK(clknet_3_4_0_clk),
    .D(_109_),
    .QN(_050_));
 DFFHQNx2_ASAP7_75t_R \mem[3][22]$_DFFE_PP_  (.CLK(clknet_3_6_0_clk),
    .D(_110_),
    .QN(_049_));
 DFFHQNx2_ASAP7_75t_R \mem[3][23]$_DFFE_PP_  (.CLK(clknet_3_6_0_clk),
    .D(_111_),
    .QN(_048_));
 DFFHQNx2_ASAP7_75t_R \mem[3][24]$_DFFE_PP_  (.CLK(clknet_3_4_0_clk),
    .D(_112_),
    .QN(_047_));
 DFFHQNx2_ASAP7_75t_R \mem[3][25]$_DFFE_PP_  (.CLK(clknet_3_6_0_clk),
    .D(_113_),
    .QN(_046_));
 DFFHQNx2_ASAP7_75t_R \mem[3][26]$_DFFE_PP_  (.CLK(clknet_3_7_0_clk),
    .D(_114_),
    .QN(_045_));
 DFFHQNx2_ASAP7_75t_R \mem[3][27]$_DFFE_PP_  (.CLK(clknet_3_5_0_clk),
    .D(_115_),
    .QN(_044_));
 DFFHQNx2_ASAP7_75t_R \mem[3][28]$_DFFE_PP_  (.CLK(clknet_3_5_0_clk),
    .D(_116_),
    .QN(_043_));
 DFFHQNx2_ASAP7_75t_R \mem[3][29]$_DFFE_PP_  (.CLK(clknet_3_7_0_clk),
    .D(_117_),
    .QN(_042_));
 DFFHQNx2_ASAP7_75t_R \mem[3][2]$_DFFE_PP_  (.CLK(clknet_3_7_0_clk),
    .D(_118_),
    .QN(_041_));
 DFFHQNx2_ASAP7_75t_R \mem[3][30]$_DFFE_PP_  (.CLK(clknet_3_7_0_clk),
    .D(_119_),
    .QN(_040_));
 DFFHQNx2_ASAP7_75t_R \mem[3][31]$_DFFE_PP_  (.CLK(clknet_3_6_0_clk),
    .D(_120_),
    .QN(_039_));
 DFFHQNx2_ASAP7_75t_R \mem[3][3]$_DFFE_PP_  (.CLK(clknet_3_7_0_clk),
    .D(_121_),
    .QN(_038_));
 DFFHQNx2_ASAP7_75t_R \mem[3][4]$_DFFE_PP_  (.CLK(clknet_3_5_0_clk),
    .D(_122_),
    .QN(_037_));
 DFFHQNx2_ASAP7_75t_R \mem[3][5]$_DFFE_PP_  (.CLK(clknet_3_7_0_clk),
    .D(_123_),
    .QN(_036_));
 DFFHQNx2_ASAP7_75t_R \mem[3][6]$_DFFE_PP_  (.CLK(clknet_3_4_0_clk),
    .D(_124_),
    .QN(_035_));
 DFFHQNx2_ASAP7_75t_R \mem[3][7]$_DFFE_PP_  (.CLK(clknet_3_6_0_clk),
    .D(_125_),
    .QN(_034_));
 DFFHQNx2_ASAP7_75t_R \mem[3][8]$_DFFE_PP_  (.CLK(clknet_3_1_0_clk),
    .D(_126_),
    .QN(_033_));
 DFFHQNx2_ASAP7_75t_R \mem[3][9]$_DFFE_PP_  (.CLK(clknet_3_1_0_clk),
    .D(_127_),
    .QN(_064_));
 DFFHQNx3_ASAP7_75t_R \rd_out[0]$_DFF_P_  (.CLK(clknet_3_3_0_clk),
    .D(_000_),
    .QN(_065_));
 DFFHQNx3_ASAP7_75t_R \rd_out[10]$_DFF_P_  (.CLK(clknet_3_2_0_clk),
    .D(_001_),
    .QN(_066_));
 DFFHQNx3_ASAP7_75t_R \rd_out[11]$_DFF_P_  (.CLK(clknet_3_0_0_clk),
    .D(_002_),
    .QN(_067_));
 DFFHQNx3_ASAP7_75t_R \rd_out[12]$_DFF_P_  (.CLK(clknet_3_2_0_clk),
    .D(_003_),
    .QN(_068_));
 DFFHQNx3_ASAP7_75t_R \rd_out[13]$_DFF_P_  (.CLK(clknet_3_2_0_clk),
    .D(_004_),
    .QN(_069_));
 DFFHQNx3_ASAP7_75t_R \rd_out[14]$_DFF_P_  (.CLK(clknet_3_0_0_clk),
    .D(_005_),
    .QN(_070_));
 DFFHQNx3_ASAP7_75t_R \rd_out[15]$_DFF_P_  (.CLK(clknet_3_0_0_clk),
    .D(_006_),
    .QN(_071_));
 DFFHQNx3_ASAP7_75t_R \rd_out[16]$_DFF_P_  (.CLK(clknet_3_0_0_clk),
    .D(_007_),
    .QN(_072_));
 DFFHQNx3_ASAP7_75t_R \rd_out[17]$_DFF_P_  (.CLK(clknet_3_1_0_clk),
    .D(_008_),
    .QN(_073_));
 DFFHQNx3_ASAP7_75t_R \rd_out[18]$_DFF_P_  (.CLK(clknet_3_3_0_clk),
    .D(_009_),
    .QN(_074_));
 DFFHQNx3_ASAP7_75t_R \rd_out[19]$_DFF_P_  (.CLK(clknet_3_3_0_clk),
    .D(_010_),
    .QN(_075_));
 DFFHQNx3_ASAP7_75t_R \rd_out[1]$_DFF_P_  (.CLK(clknet_3_1_0_clk),
    .D(_011_),
    .QN(_076_));
 DFFHQNx3_ASAP7_75t_R \rd_out[20]$_DFF_P_  (.CLK(clknet_3_4_0_clk),
    .D(_012_),
    .QN(_077_));
 DFFHQNx3_ASAP7_75t_R \rd_out[21]$_DFF_P_  (.CLK(clknet_3_4_0_clk),
    .D(_013_),
    .QN(_078_));
 DFFHQNx3_ASAP7_75t_R \rd_out[22]$_DFF_P_  (.CLK(clknet_3_6_0_clk),
    .D(_014_),
    .QN(_079_));
 DFFHQNx3_ASAP7_75t_R \rd_out[23]$_DFF_P_  (.CLK(clknet_3_6_0_clk),
    .D(_015_),
    .QN(_080_));
 DFFHQNx3_ASAP7_75t_R \rd_out[24]$_DFF_P_  (.CLK(clknet_3_4_0_clk),
    .D(_016_),
    .QN(_081_));
 DFFHQNx3_ASAP7_75t_R \rd_out[25]$_DFF_P_  (.CLK(clknet_3_6_0_clk),
    .D(_017_),
    .QN(_082_));
 DFFHQNx3_ASAP7_75t_R \rd_out[26]$_DFF_P_  (.CLK(clknet_3_7_0_clk),
    .D(_018_),
    .QN(_083_));
 DFFHQNx3_ASAP7_75t_R \rd_out[27]$_DFF_P_  (.CLK(clknet_3_5_0_clk),
    .D(_019_),
    .QN(_084_));
 DFFHQNx3_ASAP7_75t_R \rd_out[28]$_DFF_P_  (.CLK(clknet_3_5_0_clk),
    .D(_020_),
    .QN(_085_));
 DFFHQNx3_ASAP7_75t_R \rd_out[29]$_DFF_P_  (.CLK(clknet_3_5_0_clk),
    .D(_021_),
    .QN(_086_));
 DFFHQNx3_ASAP7_75t_R \rd_out[2]$_DFF_P_  (.CLK(clknet_3_7_0_clk),
    .D(_022_),
    .QN(_087_));
 DFFHQNx3_ASAP7_75t_R \rd_out[30]$_DFF_P_  (.CLK(clknet_3_6_0_clk),
    .D(_023_),
    .QN(_088_));
 DFFHQNx3_ASAP7_75t_R \rd_out[31]$_DFF_P_  (.CLK(clknet_3_4_0_clk),
    .D(_024_),
    .QN(_089_));
 DFFHQNx3_ASAP7_75t_R \rd_out[3]$_DFF_P_  (.CLK(clknet_3_7_0_clk),
    .D(_025_),
    .QN(_090_));
 DFFHQNx3_ASAP7_75t_R \rd_out[4]$_DFF_P_  (.CLK(clknet_3_5_0_clk),
    .D(_026_),
    .QN(_091_));
 DFFHQNx3_ASAP7_75t_R \rd_out[5]$_DFF_P_  (.CLK(clknet_3_7_0_clk),
    .D(_027_),
    .QN(_092_));
 DFFHQNx3_ASAP7_75t_R \rd_out[6]$_DFF_P_  (.CLK(clknet_3_1_0_clk),
    .D(_028_),
    .QN(_093_));
 DFFHQNx3_ASAP7_75t_R \rd_out[7]$_DFF_P_  (.CLK(clknet_3_1_0_clk),
    .D(_029_),
    .QN(_094_));
 DFFHQNx3_ASAP7_75t_R \rd_out[8]$_DFF_P_  (.CLK(clknet_3_3_0_clk),
    .D(_030_),
    .QN(_095_));
 DFFHQNx3_ASAP7_75t_R \rd_out[9]$_DFF_P_  (.CLK(clknet_3_1_0_clk),
    .D(_031_),
    .QN(_032_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Left_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Left_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Left_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Left_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Left_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Left_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Left_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Left_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Left_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Left_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Left_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Left_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Left_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Left_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Left_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_185 ();
 BUFx2_ASAP7_75t_R input1 (.A(addr_in[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_R input2 (.A(addr_in[1]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input3 (.A(wd_in[0]),
    .Y(net3));
 BUFx2_ASAP7_75t_R input4 (.A(wd_in[10]),
    .Y(net4));
 BUFx2_ASAP7_75t_R input5 (.A(wd_in[11]),
    .Y(net5));
 BUFx2_ASAP7_75t_R input6 (.A(wd_in[12]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input7 (.A(wd_in[13]),
    .Y(net7));
 BUFx2_ASAP7_75t_R input8 (.A(wd_in[14]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input9 (.A(wd_in[15]),
    .Y(net9));
 BUFx2_ASAP7_75t_R input10 (.A(wd_in[16]),
    .Y(net10));
 BUFx2_ASAP7_75t_R input11 (.A(wd_in[17]),
    .Y(net11));
 BUFx2_ASAP7_75t_R input12 (.A(wd_in[18]),
    .Y(net12));
 BUFx2_ASAP7_75t_R input13 (.A(wd_in[19]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input14 (.A(wd_in[1]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input15 (.A(wd_in[20]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input16 (.A(wd_in[21]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input17 (.A(wd_in[22]),
    .Y(net17));
 BUFx2_ASAP7_75t_R input18 (.A(wd_in[23]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input19 (.A(wd_in[24]),
    .Y(net19));
 BUFx2_ASAP7_75t_R input20 (.A(wd_in[25]),
    .Y(net20));
 BUFx2_ASAP7_75t_R input21 (.A(wd_in[26]),
    .Y(net21));
 BUFx2_ASAP7_75t_R input22 (.A(wd_in[27]),
    .Y(net22));
 BUFx2_ASAP7_75t_R input23 (.A(wd_in[28]),
    .Y(net23));
 BUFx2_ASAP7_75t_R input24 (.A(wd_in[29]),
    .Y(net24));
 BUFx2_ASAP7_75t_R input25 (.A(wd_in[2]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input26 (.A(wd_in[30]),
    .Y(net26));
 BUFx2_ASAP7_75t_R input27 (.A(wd_in[31]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input28 (.A(wd_in[3]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input29 (.A(wd_in[4]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input30 (.A(wd_in[5]),
    .Y(net30));
 BUFx2_ASAP7_75t_R input31 (.A(wd_in[6]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input32 (.A(wd_in[7]),
    .Y(net32));
 BUFx2_ASAP7_75t_R input33 (.A(wd_in[8]),
    .Y(net33));
 BUFx2_ASAP7_75t_R input34 (.A(wd_in[9]),
    .Y(net34));
 BUFx2_ASAP7_75t_R output35 (.A(net35),
    .Y(rd_out[0]));
 BUFx2_ASAP7_75t_R output36 (.A(net36),
    .Y(rd_out[10]));
 BUFx2_ASAP7_75t_R output37 (.A(net37),
    .Y(rd_out[11]));
 BUFx2_ASAP7_75t_R output38 (.A(net38),
    .Y(rd_out[12]));
 BUFx2_ASAP7_75t_R output39 (.A(net39),
    .Y(rd_out[13]));
 BUFx2_ASAP7_75t_R output40 (.A(net40),
    .Y(rd_out[14]));
 BUFx2_ASAP7_75t_R output41 (.A(net41),
    .Y(rd_out[15]));
 BUFx2_ASAP7_75t_R output42 (.A(net42),
    .Y(rd_out[16]));
 BUFx2_ASAP7_75t_R output43 (.A(net43),
    .Y(rd_out[17]));
 BUFx2_ASAP7_75t_R output44 (.A(net44),
    .Y(rd_out[18]));
 BUFx2_ASAP7_75t_R output45 (.A(net45),
    .Y(rd_out[19]));
 BUFx2_ASAP7_75t_R output46 (.A(net46),
    .Y(rd_out[1]));
 BUFx2_ASAP7_75t_R output47 (.A(net47),
    .Y(rd_out[20]));
 BUFx2_ASAP7_75t_R output48 (.A(net48),
    .Y(rd_out[21]));
 BUFx2_ASAP7_75t_R output49 (.A(net49),
    .Y(rd_out[22]));
 BUFx2_ASAP7_75t_R output50 (.A(net50),
    .Y(rd_out[23]));
 BUFx2_ASAP7_75t_R output51 (.A(net51),
    .Y(rd_out[24]));
 BUFx2_ASAP7_75t_R output52 (.A(net52),
    .Y(rd_out[25]));
 BUFx2_ASAP7_75t_R output53 (.A(net53),
    .Y(rd_out[26]));
 BUFx2_ASAP7_75t_R output54 (.A(net54),
    .Y(rd_out[27]));
 BUFx2_ASAP7_75t_R output55 (.A(net55),
    .Y(rd_out[28]));
 BUFx2_ASAP7_75t_R output56 (.A(net56),
    .Y(rd_out[29]));
 BUFx2_ASAP7_75t_R output57 (.A(net57),
    .Y(rd_out[2]));
 BUFx2_ASAP7_75t_R output58 (.A(net58),
    .Y(rd_out[30]));
 BUFx2_ASAP7_75t_R output59 (.A(net59),
    .Y(rd_out[31]));
 BUFx2_ASAP7_75t_R output60 (.A(net60),
    .Y(rd_out[3]));
 BUFx2_ASAP7_75t_R output61 (.A(net61),
    .Y(rd_out[4]));
 BUFx2_ASAP7_75t_R output62 (.A(net62),
    .Y(rd_out[5]));
 BUFx2_ASAP7_75t_R output63 (.A(net63),
    .Y(rd_out[6]));
 BUFx2_ASAP7_75t_R output64 (.A(net64),
    .Y(rd_out[7]));
 BUFx2_ASAP7_75t_R output65 (.A(net65),
    .Y(rd_out[8]));
 BUFx2_ASAP7_75t_R output66 (.A(net66),
    .Y(rd_out[9]));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_0_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_1_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_2_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_3_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_4_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_5_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_6_0_clk));
 BUFx10_ASAP7_75t_R clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .Y(clknet_3_7_0_clk));
 BUFx12_ASAP7_75t_R clkload0 (.A(clknet_3_0_0_clk));
 BUFx4f_ASAP7_75t_R clkload1 (.A(clknet_3_1_0_clk));
 BUFx12_ASAP7_75t_R clkload2 (.A(clknet_3_2_0_clk));
 BUFx4f_ASAP7_75t_R clkload3 (.A(clknet_3_3_0_clk));
 BUFx12_ASAP7_75t_R clkload4 (.A(clknet_3_4_0_clk));
 BUFx12_ASAP7_75t_R clkload5 (.A(clknet_3_5_0_clk));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx4_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx4_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx4_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx4_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx4_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx4_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx4_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx4_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx4_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx4_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx4_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx1_ASAP7_75t_R FILLER_12_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_50 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx6_ASAP7_75t_R FILLER_14_2 ();
 FILLER_ASAP7_75t_R FILLER_14_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_18 ();
 FILLER_ASAP7_75t_R FILLER_14_44 ();
 FILLER_ASAP7_75t_R FILLER_14_54 ();
 DECAPx1_ASAP7_75t_R FILLER_15_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_30 ();
 DECAPx2_ASAP7_75t_R FILLER_17_2 ();
 FILLER_ASAP7_75t_R FILLER_17_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_10 ();
 DECAPx1_ASAP7_75t_R FILLER_17_17 ();
 FILLER_ASAP7_75t_R FILLER_17_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_55 ();
 FILLER_ASAP7_75t_R FILLER_18_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_4 ();
 FILLER_ASAP7_75t_R FILLER_18_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_28 ();
 FILLER_ASAP7_75t_R FILLER_19_2 ();
 FILLER_ASAP7_75t_R FILLER_19_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_25 ();
 FILLER_ASAP7_75t_R FILLER_20_2 ();
 FILLER_ASAP7_75t_R FILLER_20_10 ();
 FILLER_ASAP7_75t_R FILLER_20_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_55 ();
 DECAPx1_ASAP7_75t_R FILLER_21_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_32 ();
 FILLER_ASAP7_75t_R FILLER_22_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_2 ();
 FILLER_ASAP7_75t_R FILLER_27_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_27 ();
 FILLER_ASAP7_75t_R FILLER_31_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_36 ();
 FILLER_ASAP7_75t_R FILLER_36_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_25 ();
 FILLER_ASAP7_75t_R FILLER_36_54 ();
 FILLER_ASAP7_75t_R FILLER_37_2 ();
 FILLER_ASAP7_75t_R FILLER_37_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_32 ();
 FILLER_ASAP7_75t_R FILLER_38_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_2 ();
 FILLER_ASAP7_75t_R FILLER_40_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_4 ();
 FILLER_ASAP7_75t_R FILLER_40_8 ();
 FILLER_ASAP7_75t_R FILLER_40_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_47 ();
 DECAPx1_ASAP7_75t_R FILLER_40_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_55 ();
 DECAPx4_ASAP7_75t_R FILLER_41_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_12 ();
 DECAPx4_ASAP7_75t_R FILLER_42_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_33 ();
 DECAPx2_ASAP7_75t_R FILLER_43_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_2 ();
 DECAPx4_ASAP7_75t_R FILLER_44_9 ();
 FILLER_ASAP7_75t_R FILLER_44_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_21 ();
 FILLER_ASAP7_75t_R FILLER_44_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_55 ();
 DECAPx1_ASAP7_75t_R FILLER_45_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_55 ();
 FILLER_ASAP7_75t_R FILLER_46_27 ();
 FILLER_ASAP7_75t_R FILLER_46_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_50 ();
 FILLER_ASAP7_75t_R FILLER_47_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_55 ();
 DECAPx2_ASAP7_75t_R FILLER_49_24 ();
 FILLER_ASAP7_75t_R FILLER_49_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_55 ();
 DECAPx4_ASAP7_75t_R FILLER_50_2 ();
 FILLER_ASAP7_75t_R FILLER_50_12 ();
 FILLER_ASAP7_75t_R FILLER_50_26 ();
 FILLER_ASAP7_75t_R FILLER_50_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_33 ();
 DECAPx1_ASAP7_75t_R FILLER_51_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_6 ();
 DECAPx2_ASAP7_75t_R FILLER_51_20 ();
 FILLER_ASAP7_75t_R FILLER_51_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_28 ();
 FILLER_ASAP7_75t_R FILLER_52_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_4 ();
 FILLER_ASAP7_75t_R FILLER_52_54 ();
 FILLER_ASAP7_75t_R FILLER_53_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_43 ();
 FILLER_ASAP7_75t_R FILLER_53_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_31 ();
 FILLER_ASAP7_75t_R FILLER_54_35 ();
 FILLER_ASAP7_75t_R FILLER_54_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_50 ();
 FILLER_ASAP7_75t_R FILLER_55_2 ();
 FILLER_ASAP7_75t_R FILLER_56_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_24 ();
 FILLER_ASAP7_75t_R FILLER_57_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_55 ();
 FILLER_ASAP7_75t_R FILLER_58_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_35 ();
 DECAPx1_ASAP7_75t_R FILLER_59_47 ();
 FILLER_ASAP7_75t_R FILLER_60_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_2 ();
 FILLER_ASAP7_75t_R FILLER_61_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_2 ();
 FILLER_ASAP7_75t_R FILLER_63_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_55 ();
 FILLER_ASAP7_75t_R FILLER_64_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_4 ();
 FILLER_ASAP7_75t_R FILLER_65_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_4 ();
 FILLER_ASAP7_75t_R FILLER_65_26 ();
 FILLER_ASAP7_75t_R FILLER_66_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_11 ();
 FILLER_ASAP7_75t_R FILLER_67_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_2 ();
 FILLER_ASAP7_75t_R FILLER_68_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_2 ();
 FILLER_ASAP7_75t_R FILLER_69_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_2 ();
 DECAPx4_ASAP7_75t_R FILLER_79_6 ();
 DECAPx10_ASAP7_75t_R FILLER_80_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_42 ();
 DECAPx10_ASAP7_75t_R FILLER_81_2 ();
 DECAPx4_ASAP7_75t_R FILLER_81_24 ();
 FILLER_ASAP7_75t_R FILLER_81_34 ();
 DECAPx10_ASAP7_75t_R FILLER_82_2 ();
 DECAPx10_ASAP7_75t_R FILLER_82_24 ();
 DECAPx2_ASAP7_75t_R FILLER_82_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_55 ();
 DECAPx10_ASAP7_75t_R FILLER_83_2 ();
 DECAPx10_ASAP7_75t_R FILLER_83_24 ();
 DECAPx4_ASAP7_75t_R FILLER_83_46 ();
 DECAPx10_ASAP7_75t_R FILLER_84_2 ();
 DECAPx10_ASAP7_75t_R FILLER_84_24 ();
 DECAPx4_ASAP7_75t_R FILLER_84_46 ();
 DECAPx10_ASAP7_75t_R FILLER_85_2 ();
 DECAPx10_ASAP7_75t_R FILLER_85_24 ();
 DECAPx4_ASAP7_75t_R FILLER_85_46 ();
 DECAPx10_ASAP7_75t_R FILLER_86_2 ();
 DECAPx10_ASAP7_75t_R FILLER_86_24 ();
 DECAPx4_ASAP7_75t_R FILLER_86_46 ();
 DECAPx10_ASAP7_75t_R FILLER_87_2 ();
 DECAPx10_ASAP7_75t_R FILLER_87_24 ();
 DECAPx4_ASAP7_75t_R FILLER_87_46 ();
 DECAPx10_ASAP7_75t_R FILLER_88_2 ();
 DECAPx10_ASAP7_75t_R FILLER_88_24 ();
 DECAPx4_ASAP7_75t_R FILLER_88_46 ();
 DECAPx10_ASAP7_75t_R FILLER_89_2 ();
 DECAPx10_ASAP7_75t_R FILLER_89_24 ();
 DECAPx4_ASAP7_75t_R FILLER_89_46 ();
 DECAPx10_ASAP7_75t_R FILLER_90_2 ();
 DECAPx10_ASAP7_75t_R FILLER_90_24 ();
 DECAPx4_ASAP7_75t_R FILLER_90_46 ();
 DECAPx10_ASAP7_75t_R FILLER_91_2 ();
 DECAPx10_ASAP7_75t_R FILLER_91_24 ();
 DECAPx4_ASAP7_75t_R FILLER_91_46 ();
 DECAPx10_ASAP7_75t_R FILLER_92_2 ();
 DECAPx10_ASAP7_75t_R FILLER_92_24 ();
 DECAPx4_ASAP7_75t_R FILLER_92_46 ();
endmodule
