module ibex_id_stage (branch_decision_i,
    clk_i,
    csr_access_o,
    csr_mstatus_mie_i,
    csr_mstatus_tw_i,
    csr_op_en_o,
    csr_restore_dret_id_o,
    csr_restore_mret_id_o,
    csr_save_cause_o,
    csr_save_id_o,
    csr_save_if_o,
    csr_save_wb_o,
    ctrl_busy_o,
    data_ind_timing_i,
    debug_csr_save_o,
    debug_ebreakm_i,
    debug_ebreaku_i,
    debug_mode_o,
    debug_req_i,
    debug_single_step_i,
    div_en_ex_o,
    div_sel_ex_o,
    en_wb_o,
    ex_valid_i,
    icache_inval_o,
    id_in_ready_o,
    illegal_c_insn_i,
    illegal_csr_insn_i,
    illegal_insn_o,
    instr_bp_taken_i,
    instr_fetch_err_i,
    instr_fetch_err_plus2_i,
    instr_first_cycle_id_o,
    instr_id_done_o,
    instr_is_compressed_i,
    instr_perf_count_id_o,
    instr_req_o,
    instr_valid_clear_o,
    instr_valid_i,
    irq_nm_i,
    irq_pending_i,
    lsu_addr_incr_req_i,
    lsu_load_err_i,
    lsu_req_done_i,
    lsu_req_o,
    lsu_resp_valid_i,
    lsu_sign_ext_o,
    lsu_store_err_i,
    lsu_we_o,
    mult_en_ex_o,
    mult_sel_ex_o,
    multdiv_ready_id_o,
    nmi_mode_o,
    nt_branch_mispredict_o,
    outstanding_load_wb_i,
    outstanding_store_wb_i,
    pc_set_o,
    pc_set_spec_o,
    perf_branch_o,
    perf_div_wait_o,
    perf_dside_wait_o,
    perf_jump_o,
    perf_mul_wait_o,
    perf_tbranch_o,
    ready_wb_i,
    rf_rd_a_wb_match_o,
    rf_rd_b_wb_match_o,
    rf_ren_a_o,
    rf_ren_b_o,
    rf_we_id_o,
    rf_write_wb_i,
    rst_ni,
    trigger_match_i,
    alu_operand_a_ex_o,
    alu_operand_b_ex_o,
    alu_operator_ex_o,
    bt_a_operand_o,
    bt_b_operand_o,
    csr_mtval_o,
    csr_op_o,
    csr_rdata_i,
    debug_cause_o,
    exc_cause_o,
    exc_pc_mux_o,
    imd_val_d_ex_i,
    imd_val_q_ex_o,
    imd_val_we_ex_i,
    instr_rdata_alu_i,
    instr_rdata_c_i,
    instr_rdata_i,
    instr_type_wb_o,
    irqs_i,
    lsu_addr_last_i,
    lsu_type_o,
    lsu_wdata_o,
    multdiv_operand_a_ex_o,
    multdiv_operand_b_ex_o,
    multdiv_operator_ex_o,
    multdiv_signed_mode_ex_o,
    pc_id_i,
    pc_mux_o,
    priv_mode_i,
    result_ex_i,
    rf_raddr_a_o,
    rf_raddr_b_o,
    rf_rdata_a_i,
    rf_rdata_b_i,
    rf_waddr_id_o,
    rf_waddr_wb_i,
    rf_wdata_fwd_wb_i,
    rf_wdata_id_o);
 input branch_decision_i;
 input clk_i;
 output csr_access_o;
 input csr_mstatus_mie_i;
 input csr_mstatus_tw_i;
 output csr_op_en_o;
 output csr_restore_dret_id_o;
 output csr_restore_mret_id_o;
 output csr_save_cause_o;
 output csr_save_id_o;
 output csr_save_if_o;
 output csr_save_wb_o;
 output ctrl_busy_o;
 input data_ind_timing_i;
 output debug_csr_save_o;
 input debug_ebreakm_i;
 input debug_ebreaku_i;
 output debug_mode_o;
 input debug_req_i;
 input debug_single_step_i;
 output div_en_ex_o;
 output div_sel_ex_o;
 output en_wb_o;
 input ex_valid_i;
 output icache_inval_o;
 output id_in_ready_o;
 input illegal_c_insn_i;
 input illegal_csr_insn_i;
 output illegal_insn_o;
 input instr_bp_taken_i;
 input instr_fetch_err_i;
 input instr_fetch_err_plus2_i;
 output instr_first_cycle_id_o;
 output instr_id_done_o;
 input instr_is_compressed_i;
 output instr_perf_count_id_o;
 output instr_req_o;
 output instr_valid_clear_o;
 input instr_valid_i;
 input irq_nm_i;
 input irq_pending_i;
 input lsu_addr_incr_req_i;
 input lsu_load_err_i;
 input lsu_req_done_i;
 output lsu_req_o;
 input lsu_resp_valid_i;
 output lsu_sign_ext_o;
 input lsu_store_err_i;
 output lsu_we_o;
 output mult_en_ex_o;
 output mult_sel_ex_o;
 output multdiv_ready_id_o;
 output nmi_mode_o;
 output nt_branch_mispredict_o;
 input outstanding_load_wb_i;
 input outstanding_store_wb_i;
 output pc_set_o;
 output pc_set_spec_o;
 output perf_branch_o;
 output perf_div_wait_o;
 output perf_dside_wait_o;
 output perf_jump_o;
 output perf_mul_wait_o;
 output perf_tbranch_o;
 input ready_wb_i;
 output rf_rd_a_wb_match_o;
 output rf_rd_b_wb_match_o;
 output rf_ren_a_o;
 output rf_ren_b_o;
 output rf_we_id_o;
 input rf_write_wb_i;
 input rst_ni;
 input trigger_match_i;
 output [31:0] alu_operand_a_ex_o;
 output [31:0] alu_operand_b_ex_o;
 output [5:0] alu_operator_ex_o;
 output [31:0] bt_a_operand_o;
 output [31:0] bt_b_operand_o;
 output [31:0] csr_mtval_o;
 output [1:0] csr_op_o;
 input [31:0] csr_rdata_i;
 output [2:0] debug_cause_o;
 output [5:0] exc_cause_o;
 output [1:0] exc_pc_mux_o;
 input [67:0] imd_val_d_ex_i;
 output [67:0] imd_val_q_ex_o;
 input [1:0] imd_val_we_ex_i;
 input [31:0] instr_rdata_alu_i;
 input [15:0] instr_rdata_c_i;
 input [31:0] instr_rdata_i;
 output [1:0] instr_type_wb_o;
 input [17:0] irqs_i;
 input [31:0] lsu_addr_last_i;
 output [1:0] lsu_type_o;
 output [31:0] lsu_wdata_o;
 output [31:0] multdiv_operand_a_ex_o;
 output [31:0] multdiv_operand_b_ex_o;
 output [1:0] multdiv_operator_ex_o;
 output [1:0] multdiv_signed_mode_ex_o;
 input [31:0] pc_id_i;
 output [2:0] pc_mux_o;
 input [1:0] priv_mode_i;
 input [31:0] result_ex_i;
 output [4:0] rf_raddr_a_o;
 output [4:0] rf_raddr_b_o;
 input [31:0] rf_rdata_a_i;
 input [31:0] rf_rdata_b_i;
 output [4:0] rf_waddr_id_o;
 input [4:0] rf_waddr_wb_i;
 input [31:0] rf_wdata_fwd_wb_i;
 output [31:0] rf_wdata_id_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire clknet_0_clk_i;
 wire net802;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire branch_set;
 wire branch_set_d;
 wire \controller_i.ctrl_fsm_cs[0] ;
 wire \controller_i.ctrl_fsm_cs[1] ;
 wire \controller_i.ctrl_fsm_cs[2] ;
 wire \controller_i.ctrl_fsm_cs[3] ;
 wire \controller_i.exc_req_d ;
 wire \controller_i.exc_req_q ;
 wire \controller_i.illegal_insn_d ;
 wire \controller_i.illegal_insn_q ;
 wire \controller_i.load_err_q ;
 wire \controller_i.store_err_q ;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire id_fsm_q;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire clknet_3_0_0_clk_i;
 wire clknet_3_1_0_clk_i;
 wire clknet_3_2_0_clk_i;
 wire clknet_3_3_0_clk_i;
 wire clknet_3_4_0_clk_i;
 wire clknet_3_5_0_clk_i;
 wire clknet_3_6_0_clk_i;
 wire clknet_3_7_0_clk_i;

 sky130_fd_sc_hd__clkbuf_4 _0867_ (.A(id_fsm_q),
    .X(_0607_));
 sky130_fd_sc_hd__clkbuf_16 _0868_ (.A(instr_valid_i),
    .X(_0608_));
 sky130_fd_sc_hd__nand2b_4 _0869_ (.A_N(_0607_),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__clkinv_4 _0870_ (.A(_0609_),
    .Y(net558));
 sky130_fd_sc_hd__buf_6 _0871_ (.A(net116),
    .X(_0610_));
 sky130_fd_sc_hd__clkbuf_4 _0872_ (.A(instr_rdata_alu_i[5]),
    .X(_0611_));
 sky130_fd_sc_hd__clkbuf_4 _0873_ (.A(instr_rdata_alu_i[2]),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_4 _0874_ (.A(instr_rdata_alu_i[3]),
    .X(_0613_));
 sky130_fd_sc_hd__nor4bb_2 _0875_ (.A(_0612_),
    .B(_0613_),
    .C_N(net114),
    .D_N(net117),
    .Y(_0614_));
 sky130_fd_sc_hd__clkbuf_4 _0876_ (.A(net126),
    .X(_0615_));
 sky130_fd_sc_hd__clkbuf_4 _0877_ (.A(net125),
    .X(_0616_));
 sky130_fd_sc_hd__nor2b_4 _0878_ (.A(_0615_),
    .B_N(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand3_4 _0879_ (.A(_0611_),
    .B(_0614_),
    .C(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__or4_4 _0880_ (.A(net120),
    .B(net122),
    .C(net121),
    .D(net124),
    .X(_0619_));
 sky130_fd_sc_hd__nor3_4 _0881_ (.A(net119),
    .B(net123),
    .C(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nand2_4 _0882_ (.A(net118),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__nor3_4 _0883_ (.A(_0610_),
    .B(_0618_),
    .C(_0621_),
    .Y(net601));
 sky130_fd_sc_hd__inv_6 _0884_ (.A(net116),
    .Y(_0622_));
 sky130_fd_sc_hd__nor3_4 _0885_ (.A(_0622_),
    .B(_0618_),
    .C(_0621_),
    .Y(net477));
 sky130_fd_sc_hd__clkbuf_4 _0886_ (.A(instr_rdata_i[12]),
    .X(_0623_));
 sky130_fd_sc_hd__or3_4 _0887_ (.A(net146),
    .B(_0623_),
    .C(net147),
    .X(_0624_));
 sky130_fd_sc_hd__buf_4 _0888_ (.A(instr_rdata_i[2]),
    .X(_0625_));
 sky130_fd_sc_hd__nand4bb_4 _0889_ (.A_N(net165),
    .B_N(_0625_),
    .C(net143),
    .D(net153),
    .Y(_0626_));
 sky130_fd_sc_hd__buf_4 _0890_ (.A(instr_rdata_i[6]),
    .X(_0627_));
 sky130_fd_sc_hd__buf_4 _0891_ (.A(net166),
    .X(_0628_));
 sky130_fd_sc_hd__nand3_4 _0892_ (.A(_0627_),
    .B(_0628_),
    .C(net167),
    .Y(_0629_));
 sky130_fd_sc_hd__nor2_4 _0893_ (.A(_0626_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_4 _0894_ (.A(_0624_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__buf_4 _0895_ (.A(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__buf_6 _0896_ (.A(net147),
    .X(_0633_));
 sky130_fd_sc_hd__nor2_2 _0897_ (.A(net146),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__buf_4 _0898_ (.A(_0627_),
    .X(_0635_));
 sky130_fd_sc_hd__buf_4 _0899_ (.A(net167),
    .X(_0636_));
 sky130_fd_sc_hd__nor3_1 _0900_ (.A(_0633_),
    .B(net165),
    .C(_0625_),
    .Y(_0637_));
 sky130_fd_sc_hd__nor3b_4 _0901_ (.A(_0627_),
    .B(net167),
    .C_N(net165),
    .Y(_0638_));
 sky130_fd_sc_hd__a32oi_2 _0902_ (.A1(_0635_),
    .A2(_0636_),
    .A3(_0637_),
    .B1(_0638_),
    .B2(_0625_),
    .Y(_0639_));
 sky130_fd_sc_hd__nor3_1 _0903_ (.A(_0628_),
    .B(_0634_),
    .C(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__buf_8 _0904_ (.A(net164),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _0905_ (.A(net159),
    .B(net160),
    .C(net161),
    .D(net162),
    .X(_0642_));
 sky130_fd_sc_hd__nor2_1 _0906_ (.A(_0641_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__clkinv_2 _0907_ (.A(_0633_),
    .Y(_0644_));
 sky130_fd_sc_hd__buf_6 _0908_ (.A(net163),
    .X(_0645_));
 sky130_fd_sc_hd__buf_16 _0909_ (.A(instr_rdata_i[25]),
    .X(_0646_));
 sky130_fd_sc_hd__a21oi_1 _0910_ (.A1(_0644_),
    .A2(_0645_),
    .B1(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2b_4 _0911_ (.A_N(_0627_),
    .B(net166),
    .Y(_0648_));
 sky130_fd_sc_hd__nand2b_1 _0912_ (.A_N(net146),
    .B(_0623_),
    .Y(_0649_));
 sky130_fd_sc_hd__or4_1 _0913_ (.A(_0636_),
    .B(_0626_),
    .C(_0648_),
    .D(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a21oi_1 _0914_ (.A1(_0643_),
    .A2(_0647_),
    .B1(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__nand2b_1 _0915_ (.A_N(_0628_),
    .B(_0625_),
    .Y(_0652_));
 sky130_fd_sc_hd__a21oi_1 _0916_ (.A1(_0635_),
    .A2(_0636_),
    .B1(_0638_),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_1 _0917_ (.A(net165),
    .Y(_0654_));
 sky130_fd_sc_hd__nor2b_1 _0918_ (.A(_0636_),
    .B_N(_0627_),
    .Y(_0655_));
 sky130_fd_sc_hd__o21ai_1 _0919_ (.A1(_0625_),
    .A2(_0655_),
    .B1(_0648_),
    .Y(_0656_));
 sky130_fd_sc_hd__a2bb2oi_4 _0920_ (.A1_N(_0652_),
    .A2_N(_0653_),
    .B1(_0654_),
    .B2(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nor3_4 _0921_ (.A(_0640_),
    .B(_0651_),
    .C(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__buf_8 _0922_ (.A(net146),
    .X(_0659_));
 sky130_fd_sc_hd__buf_6 _0923_ (.A(_0623_),
    .X(_0660_));
 sky130_fd_sc_hd__or2_2 _0924_ (.A(_0626_),
    .B(_0629_),
    .X(_0661_));
 sky130_fd_sc_hd__nor3_4 _0925_ (.A(_0659_),
    .B(_0660_),
    .C(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__nor2_1 _0926_ (.A(net150),
    .B(net152),
    .Y(_0663_));
 sky130_fd_sc_hd__nor3_1 _0927_ (.A(net149),
    .B(net148),
    .C(net151),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _0928_ (.A(_0663_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__or4_1 _0929_ (.A(net147),
    .B(net169),
    .C(net168),
    .D(net144),
    .X(_0666_));
 sky130_fd_sc_hd__or4_2 _0930_ (.A(net170),
    .B(net145),
    .C(_0665_),
    .D(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__and4bb_4 _0931_ (.A_N(net165),
    .B_N(_0625_),
    .C(net143),
    .D(net153),
    .X(_0668_));
 sky130_fd_sc_hd__nor2_2 _0932_ (.A(_0627_),
    .B(_0628_),
    .Y(_0669_));
 sky130_fd_sc_hd__o2111ai_2 _0933_ (.A1(_0623_),
    .A2(_0633_),
    .B1(_0668_),
    .C1(_0669_),
    .D1(_0659_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2b_2 _0934_ (.A(_0628_),
    .B_N(_0636_),
    .Y(_0671_));
 sky130_fd_sc_hd__xnor2_1 _0935_ (.A(_0625_),
    .B(_0627_),
    .Y(_0672_));
 sky130_fd_sc_hd__and4b_1 _0936_ (.A_N(net165),
    .B(net153),
    .C(net143),
    .D(net147),
    .X(_0673_));
 sky130_fd_sc_hd__nand3_1 _0937_ (.A(_0671_),
    .B(_0672_),
    .C(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _0938_ (.A(net143),
    .B(net153),
    .Y(_0675_));
 sky130_fd_sc_hd__nor2_1 _0939_ (.A(net42),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__nor2_1 _0940_ (.A(net146),
    .B(_0623_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand4b_2 _0941_ (.A_N(_0628_),
    .B(_0636_),
    .C(_0625_),
    .D(_0627_),
    .Y(_0678_));
 sky130_fd_sc_hd__or3_1 _0942_ (.A(net165),
    .B(_0677_),
    .C(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__nand4_4 _0943_ (.A(_0670_),
    .B(_0674_),
    .C(_0676_),
    .D(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__xor2_1 _0944_ (.A(_0623_),
    .B(net147),
    .X(_0681_));
 sky130_fd_sc_hd__o31ai_1 _0945_ (.A1(net146),
    .A2(_0646_),
    .A3(_0681_),
    .B1(_0645_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_2 _0946_ (.A(_0636_),
    .B(_0668_),
    .Y(_0683_));
 sky130_fd_sc_hd__a211oi_2 _0947_ (.A1(_0643_),
    .A2(_0682_),
    .B1(_0683_),
    .C1(_0648_),
    .Y(_0684_));
 sky130_fd_sc_hd__a211oi_4 _0948_ (.A1(_0662_),
    .A2(_0667_),
    .B1(_0680_),
    .C1(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__nor4b_2 _0949_ (.A(net154),
    .B(net157),
    .C(net156),
    .D_N(net155),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2_2 _0950_ (.A(_0645_),
    .B(_0641_),
    .Y(_0687_));
 sky130_fd_sc_hd__and4_2 _0951_ (.A(net161),
    .B(net162),
    .C(_0686_),
    .D(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__buf_6 _0952_ (.A(net154),
    .X(_0689_));
 sky130_fd_sc_hd__nor4_2 _0953_ (.A(net155),
    .B(net157),
    .C(_0645_),
    .D(net164),
    .Y(_0690_));
 sky130_fd_sc_hd__nor2b_1 _0954_ (.A(net162),
    .B_N(net161),
    .Y(_0691_));
 sky130_fd_sc_hd__and4_1 _0955_ (.A(_0689_),
    .B(net156),
    .C(_0690_),
    .D(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__nor4_4 _0956_ (.A(net158),
    .B(_0646_),
    .C(net159),
    .D(net160),
    .Y(_0693_));
 sky130_fd_sc_hd__o21a_1 _0957_ (.A1(_0688_),
    .A2(_0692_),
    .B1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__and4b_1 _0958_ (.A_N(net159),
    .B(net160),
    .C(_0645_),
    .D(_0646_),
    .X(_0695_));
 sky130_fd_sc_hd__and4b_1 _0959_ (.A_N(_0641_),
    .B(net162),
    .C(net161),
    .D(net158),
    .X(_0696_));
 sky130_fd_sc_hd__nand3_4 _0960_ (.A(_0686_),
    .B(_0695_),
    .C(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__nor3_2 _0961_ (.A(net155),
    .B(net163),
    .C(net164),
    .Y(_0698_));
 sky130_fd_sc_hd__nor4_2 _0962_ (.A(net157),
    .B(net156),
    .C(net161),
    .D(net162),
    .Y(_0699_));
 sky130_fd_sc_hd__nand3_4 _0963_ (.A(_0693_),
    .B(_0698_),
    .C(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand4b_4 _0964_ (.A_N(_0694_),
    .B(_0697_),
    .C(_0700_),
    .D(_0662_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand3_4 _0965_ (.A(_0658_),
    .B(_0685_),
    .C(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__nor2_2 _0966_ (.A(_0632_),
    .B(_0702_),
    .Y(net429));
 sky130_fd_sc_hd__o21a_2 _0967_ (.A1(net43),
    .A2(_0702_),
    .B1(_0608_),
    .X(net489));
 sky130_fd_sc_hd__buf_6 _0968_ (.A(\controller_i.ctrl_fsm_cs[0] ),
    .X(_0703_));
 sky130_fd_sc_hd__buf_4 _0969_ (.A(\controller_i.ctrl_fsm_cs[3] ),
    .X(_0704_));
 sky130_fd_sc_hd__nor2b_2 _0970_ (.A(_0704_),
    .B_N(\controller_i.ctrl_fsm_cs[1] ),
    .Y(_0705_));
 sky130_fd_sc_hd__nand2_2 _0971_ (.A(\controller_i.ctrl_fsm_cs[2] ),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__nor2_8 _0972_ (.A(_0703_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__or4_1 _0973_ (.A(net158),
    .B(_0646_),
    .C(net159),
    .D(net160),
    .X(_0708_));
 sky130_fd_sc_hd__a21oi_1 _0974_ (.A1(net3),
    .A2(_0692_),
    .B1(_0688_),
    .Y(_0709_));
 sky130_fd_sc_hd__and2_0 _0975_ (.A(net258),
    .B(net259),
    .X(_0710_));
 sky130_fd_sc_hd__buf_6 _0976_ (.A(net475),
    .X(_0711_));
 sky130_fd_sc_hd__o32ai_2 _0977_ (.A1(_0708_),
    .A2(_0709_),
    .A3(_0710_),
    .B1(_0697_),
    .B2(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__clkinv_4 _0978_ (.A(_0608_),
    .Y(_0713_));
 sky130_fd_sc_hd__nor4_4 _0979_ (.A(_0713_),
    .B(_0624_),
    .C(_0626_),
    .D(_0629_),
    .Y(_0714_));
 sky130_fd_sc_hd__buf_4 _0980_ (.A(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__a21oi_1 _0981_ (.A1(_0712_),
    .A2(_0715_),
    .B1(net489),
    .Y(_0716_));
 sky130_fd_sc_hd__nor2_1 _0982_ (.A(_0707_),
    .B(_0716_),
    .Y(\controller_i.illegal_insn_d ));
 sky130_fd_sc_hd__buf_6 _0983_ (.A(instr_fetch_err_i),
    .X(_0717_));
 sky130_fd_sc_hd__nor3_2 _0984_ (.A(_0717_),
    .B(net43),
    .C(_0702_),
    .Y(_0718_));
 sky130_fd_sc_hd__and3_1 _0985_ (.A(_0693_),
    .B(_0698_),
    .C(_0699_),
    .X(_0719_));
 sky130_fd_sc_hd__buf_2 _0986_ (.A(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__o21ai_0 _0987_ (.A1(_0720_),
    .A2(_0712_),
    .B1(_0715_),
    .Y(_0721_));
 sky130_fd_sc_hd__clkinv_4 _0988_ (.A(\controller_i.ctrl_fsm_cs[0] ),
    .Y(_0722_));
 sky130_fd_sc_hd__and2_2 _0989_ (.A(\controller_i.ctrl_fsm_cs[2] ),
    .B(_0705_),
    .X(_0723_));
 sky130_fd_sc_hd__nand2_2 _0990_ (.A(_0722_),
    .B(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__nand2_1 _0991_ (.A(_0608_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__a21oi_1 _0992_ (.A1(_0718_),
    .A2(_0721_),
    .B1(_0725_),
    .Y(\controller_i.exc_req_d ));
 sky130_fd_sc_hd__clkinv_2 _0993_ (.A(\controller_i.ctrl_fsm_cs[2] ),
    .Y(_0726_));
 sky130_fd_sc_hd__or3_1 _0994_ (.A(\controller_i.ctrl_fsm_cs[1] ),
    .B(\controller_i.ctrl_fsm_cs[3] ),
    .C(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__clkbuf_4 _0995_ (.A(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__a21oi_1 _0996_ (.A1(net172),
    .A2(net2),
    .B1(net171),
    .Y(_0729_));
 sky130_fd_sc_hd__nor3_4 _0997_ (.A(_0711_),
    .B(net671),
    .C(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__a211oi_2 _0998_ (.A1(net40),
    .A2(_0608_),
    .B1(net358),
    .C1(net39),
    .Y(_0731_));
 sky130_fd_sc_hd__nor2_2 _0999_ (.A(_0711_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__nor2_1 _1000_ (.A(_0730_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(_0697_),
    .B(_0700_),
    .Y(_0734_));
 sky130_fd_sc_hd__nor2_1 _1002_ (.A(_0694_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor3_4 _1003_ (.A(_0659_),
    .B(_0660_),
    .C(_0633_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand3_4 _1004_ (.A(_0608_),
    .B(_0736_),
    .C(_0630_),
    .Y(_0737_));
 sky130_fd_sc_hd__nor2_4 _1005_ (.A(net223),
    .B(net225),
    .Y(_0738_));
 sky130_fd_sc_hd__o21ai_2 _1006_ (.A1(_0735_),
    .A2(_0737_),
    .B1(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2b_1 _1007_ (.A(_0694_),
    .B_N(_0697_),
    .Y(_0740_));
 sky130_fd_sc_hd__o211ai_2 _1008_ (.A1(_0740_),
    .A2(_0737_),
    .B1(_0725_),
    .C1(_0738_),
    .Y(_0741_));
 sky130_fd_sc_hd__o41a_2 _1009_ (.A1(_0717_),
    .A2(net43),
    .A3(_0702_),
    .A4(_0739_),
    .B1(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__and3_2 _1010_ (.A(_0658_),
    .B(_0685_),
    .C(_0701_),
    .X(_0743_));
 sky130_fd_sc_hd__inv_1 _1011_ (.A(_0611_),
    .Y(_0744_));
 sky130_fd_sc_hd__nand4bb_4 _1012_ (.A_N(_0612_),
    .B_N(_0613_),
    .C(net114),
    .D(net117),
    .Y(_0745_));
 sky130_fd_sc_hd__nor2_4 _1013_ (.A(_0744_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand4_4 _1014_ (.A(net118),
    .B(_0617_),
    .C(_0620_),
    .D(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__or2_4 _1015_ (.A(_0675_),
    .B(_0652_),
    .X(_0748_));
 sky130_fd_sc_hd__a32oi_4 _1016_ (.A1(_0623_),
    .A2(_0634_),
    .A3(_0638_),
    .B1(_0635_),
    .B2(_0636_),
    .Y(_0749_));
 sky130_fd_sc_hd__nand3_4 _1017_ (.A(_0635_),
    .B(_0668_),
    .C(_0671_),
    .Y(_0750_));
 sky130_fd_sc_hd__o21a_1 _1018_ (.A1(_0748_),
    .A2(_0749_),
    .B1(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__inv_1 _1019_ (.A(net41),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_8 _1020_ (.A(_0668_),
    .B(_0669_),
    .Y(_0753_));
 sky130_fd_sc_hd__o41ai_1 _1021_ (.A1(_0635_),
    .A2(_0628_),
    .A3(net224),
    .A4(_0626_),
    .B1(net260),
    .Y(_0754_));
 sky130_fd_sc_hd__a22oi_2 _1022_ (.A1(_0752_),
    .A2(_0753_),
    .B1(_0754_),
    .B2(_0607_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand3b_2 _1023_ (.A_N(_0615_),
    .B(_0611_),
    .C(_0616_),
    .Y(_0756_));
 sky130_fd_sc_hd__or3b_1 _1024_ (.A(net119),
    .B(net123),
    .C_N(net118),
    .X(_0757_));
 sky130_fd_sc_hd__nor4_4 _1025_ (.A(_0745_),
    .B(_0756_),
    .C(_0619_),
    .D(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__nor2_2 _1026_ (.A(_0607_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__or4_4 _1027_ (.A(_0722_),
    .B(_0713_),
    .C(_0717_),
    .D(_0728_),
    .X(_0760_));
 sky130_fd_sc_hd__a2111oi_2 _1028_ (.A1(_0747_),
    .A2(_0751_),
    .B1(_0755_),
    .C1(_0759_),
    .D1(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__nor4_4 _1029_ (.A(_0722_),
    .B(_0713_),
    .C(_0717_),
    .D(_0728_),
    .Y(_0762_));
 sky130_fd_sc_hd__nor2_1 _1030_ (.A(net1),
    .B(net36),
    .Y(_0763_));
 sky130_fd_sc_hd__o22ai_4 _1031_ (.A1(_0748_),
    .A2(_0749_),
    .B1(_0750_),
    .B2(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__a21oi_1 _1032_ (.A1(net224),
    .A2(_0607_),
    .B1(_0713_),
    .Y(_0765_));
 sky130_fd_sc_hd__nor3_2 _1033_ (.A(_0635_),
    .B(_0628_),
    .C(_0626_),
    .Y(_0766_));
 sky130_fd_sc_hd__a32o_1 _1034_ (.A1(_0762_),
    .A2(_0759_),
    .A3(_0764_),
    .B1(_0765_),
    .B2(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__nor2_4 _1035_ (.A(_0761_),
    .B(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__nor2_8 _1036_ (.A(_0736_),
    .B(_0661_),
    .Y(_0769_));
 sky130_fd_sc_hd__nor4_1 _1037_ (.A(net157),
    .B(net156),
    .C(_0861_),
    .D(_0862_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand3_1 _1038_ (.A(_0695_),
    .B(_0696_),
    .C(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__and4b_1 _1039_ (.A_N(_0689_),
    .B(net161),
    .C(net162),
    .D(_0862_),
    .X(_0772_));
 sky130_fd_sc_hd__nand3_1 _1040_ (.A(_0693_),
    .B(_0690_),
    .C(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(_0771_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__and3_1 _1042_ (.A(_0769_),
    .B(_0762_),
    .C(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__and3_1 _1043_ (.A(_0743_),
    .B(_0768_),
    .C(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__nor2_2 _1044_ (.A(_0722_),
    .B(_0728_),
    .Y(_0777_));
 sky130_fd_sc_hd__o21ai_0 _1045_ (.A1(_0742_),
    .A2(_0776_),
    .B1(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nor2_4 _1046_ (.A(_0702_),
    .B(_0768_),
    .Y(_0779_));
 sky130_fd_sc_hd__and2_1 _1047_ (.A(_0726_),
    .B(_0705_),
    .X(_0780_));
 sky130_fd_sc_hd__nor3_1 _1048_ (.A(_0707_),
    .B(_0779_),
    .C(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__o211a_2 _1049_ (.A1(_0728_),
    .A2(_0733_),
    .B1(_0778_),
    .C1(_0781_),
    .X(net488));
 sky130_fd_sc_hd__nor3_2 _1050_ (.A(\controller_i.store_err_q ),
    .B(\controller_i.exc_req_q ),
    .C(\controller_i.load_err_q ),
    .Y(_0782_));
 sky130_fd_sc_hd__nand2_2 _1051_ (.A(_0707_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__nand3_1 _1052_ (.A(_0693_),
    .B(_0688_),
    .C(_0715_),
    .Y(_0784_));
 sky130_fd_sc_hd__nor2_4 _1053_ (.A(_0783_),
    .B(_0784_),
    .Y(net466));
 sky130_fd_sc_hd__nand3_4 _1054_ (.A(_0660_),
    .B(_0634_),
    .C(_0638_),
    .Y(_0785_));
 sky130_fd_sc_hd__nor3_4 _1055_ (.A(_0609_),
    .B(_0748_),
    .C(_0785_),
    .Y(net487));
 sky130_fd_sc_hd__nor2_1 _1056_ (.A(net258),
    .B(net259),
    .Y(_0786_));
 sky130_fd_sc_hd__a22o_2 _1057_ (.A1(net37),
    .A2(_0710_),
    .B1(_0786_),
    .B2(net38),
    .X(_0787_));
 sky130_fd_sc_hd__nor2_4 _1058_ (.A(\controller_i.ctrl_fsm_cs[1] ),
    .B(\controller_i.ctrl_fsm_cs[2] ),
    .Y(_0788_));
 sky130_fd_sc_hd__nor2_1 _1059_ (.A(_0722_),
    .B(_0711_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand4_4 _1060_ (.A(_0704_),
    .B(_0787_),
    .C(_0788_),
    .D(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(_0790_),
    .Y(net468));
 sky130_fd_sc_hd__nand3_1 _1062_ (.A(_0659_),
    .B(_0663_),
    .C(_0664_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand3_1 _1063_ (.A(_0660_),
    .B(_0630_),
    .C(_0791_),
    .Y(_0859_));
 sky130_fd_sc_hd__inv_1 _1064_ (.A(_0859_),
    .Y(net463));
 sky130_fd_sc_hd__nand3_1 _1065_ (.A(_0659_),
    .B(_0630_),
    .C(_0665_),
    .Y(_0860_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(_0860_),
    .Y(net464));
 sky130_fd_sc_hd__o41ai_4 _1067_ (.A1(_0717_),
    .A2(net43),
    .A3(_0702_),
    .A4(_0739_),
    .B1(_0741_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand3_1 _1068_ (.A(_0769_),
    .B(_0762_),
    .C(_0774_),
    .Y(_0793_));
 sky130_fd_sc_hd__a21o_1 _1069_ (.A1(_0768_),
    .A2(_0793_),
    .B1(_0702_),
    .X(_0794_));
 sky130_fd_sc_hd__nor2_1 _1070_ (.A(_0717_),
    .B(net43),
    .Y(_0795_));
 sky130_fd_sc_hd__a41oi_2 _1071_ (.A1(_0658_),
    .A2(_0685_),
    .A3(_0701_),
    .A4(_0795_),
    .B1(_0713_),
    .Y(_0796_));
 sky130_fd_sc_hd__o211ai_2 _1072_ (.A1(_0735_),
    .A2(_0737_),
    .B1(_0738_),
    .C1(_0703_),
    .Y(_0797_));
 sky130_fd_sc_hd__a311oi_2 _1073_ (.A1(_0743_),
    .A2(_0768_),
    .A3(_0775_),
    .B1(_0796_),
    .C1(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_0 _1074_ (.A1(\controller_i.ctrl_fsm_cs[1] ),
    .A2(_0732_),
    .B1(\controller_i.ctrl_fsm_cs[2] ),
    .Y(_0799_));
 sky130_fd_sc_hd__nor2_1 _1075_ (.A(\controller_i.ctrl_fsm_cs[0] ),
    .B(_0704_),
    .Y(_0800_));
 sky130_fd_sc_hd__or4_1 _1076_ (.A(net171),
    .B(net39),
    .C(_0711_),
    .D(net40),
    .X(_0801_));
 sky130_fd_sc_hd__nor2_2 _1077_ (.A(net172),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__nor2_1 _1078_ (.A(\controller_i.ctrl_fsm_cs[2] ),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_1 _1079_ (.A(\controller_i.ctrl_fsm_cs[1] ),
    .B(\controller_i.ctrl_fsm_cs[0] ),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_4 _1080_ (.A(_0704_),
    .B(_0788_),
    .Y(_0805_));
 sky130_fd_sc_hd__o31ai_1 _1081_ (.A1(_0704_),
    .A2(_0803_),
    .A3(_0804_),
    .B1(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__or3_4 _1082_ (.A(\controller_i.store_err_q ),
    .B(\controller_i.exc_req_q ),
    .C(\controller_i.load_err_q ),
    .X(_0807_));
 sky130_fd_sc_hd__a31oi_4 _1083_ (.A1(_0693_),
    .A2(_0688_),
    .A3(_0714_),
    .B1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__and3_1 _1084_ (.A(_0693_),
    .B(_0692_),
    .C(_0714_),
    .X(_0809_));
 sky130_fd_sc_hd__nor4b_1 _1085_ (.A(net155),
    .B(_0645_),
    .C(_0641_),
    .D_N(_0689_),
    .Y(_0810_));
 sky130_fd_sc_hd__a21oi_4 _1086_ (.A1(_0608_),
    .A2(_0717_),
    .B1(\controller_i.illegal_insn_q ),
    .Y(_0811_));
 sky130_fd_sc_hd__and4_1 _1087_ (.A(_0693_),
    .B(_0810_),
    .C(_0699_),
    .D(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__or2_2 _1088_ (.A(_0711_),
    .B(_0731_),
    .X(_0813_));
 sky130_fd_sc_hd__a31oi_2 _1089_ (.A1(_0715_),
    .A2(_0787_),
    .A3(_0812_),
    .B1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a211oi_1 _1090_ (.A1(_0808_),
    .A2(_0809_),
    .B1(_0724_),
    .C1(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__a211oi_2 _1091_ (.A1(_0799_),
    .A2(_0800_),
    .B1(_0806_),
    .C1(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__o21ai_0 _1092_ (.A1(_0722_),
    .A2(net260),
    .B1(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__a311oi_1 _1093_ (.A1(_0730_),
    .A2(_0792_),
    .A3(_0794_),
    .B1(_0798_),
    .C1(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__a21oi_2 _1094_ (.A1(_0768_),
    .A2(_0793_),
    .B1(_0702_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(_0732_),
    .B(_0816_),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_1 _1096_ (.A(_0816_),
    .Y(_0821_));
 sky130_fd_sc_hd__o32ai_1 _1097_ (.A1(_0742_),
    .A2(_0819_),
    .A3(_0820_),
    .B1(_0821_),
    .B2(_0777_),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_1 _1098_ (.A(_0730_),
    .Y(_0823_));
 sky130_fd_sc_hd__nor3_1 _1099_ (.A(_0703_),
    .B(_0728_),
    .C(_0732_),
    .Y(_0824_));
 sky130_fd_sc_hd__o311a_1 _1100_ (.A1(_0707_),
    .A2(_0779_),
    .A3(_0780_),
    .B1(_0823_),
    .C1(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__nor3_1 _1101_ (.A(_0818_),
    .B(_0822_),
    .C(_0825_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_1 _1102_ (.A(net260),
    .Y(_0826_));
 sky130_fd_sc_hd__a41oi_1 _1103_ (.A1(net260),
    .A2(_0743_),
    .A3(_0768_),
    .A4(_0775_),
    .B1(\controller_i.ctrl_fsm_cs[1] ),
    .Y(_0827_));
 sky130_fd_sc_hd__o21ai_0 _1104_ (.A1(_0826_),
    .A2(_0792_),
    .B1(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__o21ai_2 _1105_ (.A1(_0697_),
    .A2(_0737_),
    .B1(_0808_),
    .Y(_0829_));
 sky130_fd_sc_hd__nor3_1 _1106_ (.A(_0724_),
    .B(_0814_),
    .C(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__o21ai_4 _1107_ (.A1(_0722_),
    .A2(_0802_),
    .B1(_0780_),
    .Y(net470));
 sky130_fd_sc_hd__o41ai_1 _1108_ (.A1(_0703_),
    .A2(_0728_),
    .A3(_0823_),
    .A4(_0732_),
    .B1(net470),
    .Y(_0831_));
 sky130_fd_sc_hd__a21oi_2 _1109_ (.A1(_0809_),
    .A2(_0830_),
    .B1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__o31ai_1 _1110_ (.A1(_0823_),
    .A2(_0742_),
    .A3(_0819_),
    .B1(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__o31ai_2 _1111_ (.A1(_0813_),
    .A2(_0742_),
    .A3(_0819_),
    .B1(_0777_),
    .Y(_0834_));
 sky130_fd_sc_hd__a2bb2oi_1 _1112_ (.A1_N(_0828_),
    .A2_N(_0833_),
    .B1(_0832_),
    .B2(_0834_),
    .Y(_0001_));
 sky130_fd_sc_hd__nand4_1 _1113_ (.A(_0689_),
    .B(_0720_),
    .C(_0715_),
    .D(_0811_),
    .Y(_0835_));
 sky130_fd_sc_hd__nor2_1 _1114_ (.A(_0711_),
    .B(_0787_),
    .Y(_0836_));
 sky130_fd_sc_hd__or3_2 _1115_ (.A(_0782_),
    .B(_0835_),
    .C(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__and3_1 _1116_ (.A(\controller_i.ctrl_fsm_cs[2] ),
    .B(_0813_),
    .C(_0800_),
    .X(_0838_));
 sky130_fd_sc_hd__a21oi_1 _1117_ (.A1(_0704_),
    .A2(_0726_),
    .B1(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__o21ai_0 _1118_ (.A1(_0705_),
    .A2(_0788_),
    .B1(_0703_),
    .Y(_0840_));
 sky130_fd_sc_hd__o21ai_0 _1119_ (.A1(\controller_i.ctrl_fsm_cs[1] ),
    .A2(_0839_),
    .B1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__a21oi_1 _1120_ (.A1(_0815_),
    .A2(_0837_),
    .B1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__a32oi_1 _1121_ (.A1(_0703_),
    .A2(_0780_),
    .A3(_0802_),
    .B1(_0834_),
    .B2(_0842_),
    .Y(_0002_));
 sky130_fd_sc_hd__a21oi_1 _1122_ (.A1(_0792_),
    .A2(_0794_),
    .B1(_0722_),
    .Y(_0843_));
 sky130_fd_sc_hd__nand4_1 _1123_ (.A(_0689_),
    .B(_0720_),
    .C(_0715_),
    .D(_0811_),
    .Y(_0844_));
 sky130_fd_sc_hd__nor3_1 _1124_ (.A(_0782_),
    .B(_0844_),
    .C(_0836_),
    .Y(_0845_));
 sky130_fd_sc_hd__o21ai_0 _1125_ (.A1(_0814_),
    .A2(_0845_),
    .B1(_0707_),
    .Y(_0846_));
 sky130_fd_sc_hd__o31ai_1 _1126_ (.A1(_0728_),
    .A2(_0813_),
    .A3(_0843_),
    .B1(_0846_),
    .Y(_0003_));
 sky130_fd_sc_hd__clkinvlp_4 _1127_ (.A(_0711_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor3_4 _1128_ (.A(_0697_),
    .B(_0737_),
    .C(_0783_),
    .Y(net465));
 sky130_fd_sc_hd__or3_2 _1129_ (.A(net39),
    .B(net40),
    .C(net358),
    .X(_0848_));
 sky130_fd_sc_hd__o211ai_4 _1130_ (.A1(_0703_),
    .A2(_0848_),
    .B1(_0788_),
    .C1(_0704_),
    .Y(_0849_));
 sky130_fd_sc_hd__o21ai_1 _1131_ (.A1(_0847_),
    .A2(net465),
    .B1(_0849_),
    .Y(_0004_));
 sky130_fd_sc_hd__a31oi_1 _1132_ (.A1(net171),
    .A2(_0723_),
    .A3(_0789_),
    .B1(net671),
    .Y(_0850_));
 sky130_fd_sc_hd__nor2_1 _1133_ (.A(net466),
    .B(_0850_),
    .Y(_0005_));
 sky130_fd_sc_hd__nand4_4 _1134_ (.A(_0658_),
    .B(_0766_),
    .C(_0685_),
    .D(_0701_),
    .Y(_0851_));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(net224),
    .A1(net41),
    .S(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_4 _1136_ (.A(_0702_),
    .B(_0760_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _1137_ (.A(net41),
    .B(_0758_),
    .Y(_0854_));
 sky130_fd_sc_hd__o21ai_0 _1138_ (.A1(_0758_),
    .A2(_0764_),
    .B1(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_1 _1139_ (.A(_0753_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21oi_1 _1140_ (.A1(_0853_),
    .A2(_0856_),
    .B1(_0607_),
    .Y(_0857_));
 sky130_fd_sc_hd__a41oi_1 _1141_ (.A1(net260),
    .A2(_0607_),
    .A3(_0762_),
    .A4(_0852_),
    .B1(_0857_),
    .Y(_0006_));
 sky130_fd_sc_hd__buf_4 _1142_ (.A(imd_val_we_ex_i[1]),
    .X(_0858_));
 sky130_fd_sc_hd__buf_4 _1143_ (.A(_0858_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1144_ (.A0(net490),
    .A1(net44),
    .S(_0075_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _1145_ (.A0(net491),
    .A1(net45),
    .S(_0075_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _1146_ (.A0(net492),
    .A1(net46),
    .S(_0075_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _1147_ (.A0(net493),
    .A1(net47),
    .S(_0075_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _1148_ (.A0(net494),
    .A1(net48),
    .S(_0075_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _1149_ (.A0(net495),
    .A1(net49),
    .S(_0075_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _1150_ (.A0(net496),
    .A1(net50),
    .S(_0075_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _1151_ (.A0(net497),
    .A1(net51),
    .S(_0075_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _1152_ (.A0(net498),
    .A1(net52),
    .S(_0075_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _1153_ (.A0(net499),
    .A1(net53),
    .S(_0075_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_4 _1154_ (.A(_0858_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1155_ (.A0(net500),
    .A1(net54),
    .S(_0076_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _1156_ (.A0(net501),
    .A1(net55),
    .S(_0076_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _1157_ (.A0(net502),
    .A1(net56),
    .S(_0076_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(net503),
    .A1(net57),
    .S(_0076_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1159_ (.A0(net504),
    .A1(net58),
    .S(_0076_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1160_ (.A0(net505),
    .A1(net59),
    .S(_0076_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1161_ (.A0(net506),
    .A1(net60),
    .S(_0076_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1162_ (.A0(net507),
    .A1(net61),
    .S(_0076_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(net508),
    .A1(net62),
    .S(_0076_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1164_ (.A0(net509),
    .A1(net63),
    .S(_0076_),
    .X(_0026_));
 sky130_fd_sc_hd__buf_4 _1165_ (.A(_0858_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1166_ (.A0(net510),
    .A1(net64),
    .S(_0077_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1167_ (.A0(net511),
    .A1(net65),
    .S(_0077_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(net512),
    .A1(net66),
    .S(_0077_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1169_ (.A0(net513),
    .A1(net67),
    .S(_0077_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1170_ (.A0(net514),
    .A1(net68),
    .S(_0077_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1171_ (.A0(net515),
    .A1(net69),
    .S(_0077_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1172_ (.A0(net516),
    .A1(net70),
    .S(_0077_),
    .X(_0033_));
 sky130_fd_sc_hd__buf_2 _1173_ (.A(imd_val_we_ex_i[0]),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_8 _1174_ (.A(_0078_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(net517),
    .A1(net71),
    .S(_0079_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1176_ (.A0(net518),
    .A1(net72),
    .S(_0079_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1177_ (.A0(net519),
    .A1(net73),
    .S(_0079_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(net520),
    .A1(net74),
    .S(_0079_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _1179_ (.A0(net521),
    .A1(net75),
    .S(_0079_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _1180_ (.A0(net522),
    .A1(net76),
    .S(_0079_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1181_ (.A0(net523),
    .A1(net77),
    .S(_0077_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(net524),
    .A1(net78),
    .S(_0079_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1183_ (.A0(net525),
    .A1(net79),
    .S(_0079_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(net526),
    .A1(net80),
    .S(_0079_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1185_ (.A0(net527),
    .A1(net81),
    .S(_0079_),
    .X(_0044_));
 sky130_fd_sc_hd__buf_4 _1186_ (.A(_0078_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1187_ (.A0(net528),
    .A1(net82),
    .S(_0080_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1188_ (.A0(net529),
    .A1(net83),
    .S(_0080_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1189_ (.A0(net530),
    .A1(net84),
    .S(_0080_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(net531),
    .A1(net85),
    .S(_0080_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1191_ (.A0(net532),
    .A1(net86),
    .S(_0080_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1192_ (.A0(net533),
    .A1(net87),
    .S(_0080_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1193_ (.A0(net534),
    .A1(net88),
    .S(_0077_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1194_ (.A0(net535),
    .A1(net89),
    .S(_0080_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(net536),
    .A1(net90),
    .S(_0080_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1196_ (.A0(net537),
    .A1(net91),
    .S(_0080_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1197_ (.A0(net538),
    .A1(net92),
    .S(_0080_),
    .X(_0055_));
 sky130_fd_sc_hd__buf_4 _1198_ (.A(_0078_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1199_ (.A0(net539),
    .A1(net93),
    .S(_0081_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(net540),
    .A1(net94),
    .S(_0081_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1201_ (.A0(net541),
    .A1(net95),
    .S(_0081_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1202_ (.A0(net542),
    .A1(net96),
    .S(_0081_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1203_ (.A0(net543),
    .A1(net97),
    .S(_0081_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1204_ (.A0(net544),
    .A1(net98),
    .S(_0081_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1205_ (.A0(net545),
    .A1(net99),
    .S(_0077_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1206_ (.A0(net546),
    .A1(net100),
    .S(_0081_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1207_ (.A0(net547),
    .A1(net101),
    .S(_0081_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1208_ (.A0(net548),
    .A1(net102),
    .S(_0081_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1209_ (.A0(net549),
    .A1(net103),
    .S(_0081_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1210_ (.A0(net550),
    .A1(net104),
    .S(_0078_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1211_ (.A0(net551),
    .A1(net105),
    .S(_0078_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1212_ (.A0(net552),
    .A1(net106),
    .S(_0078_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(net553),
    .A1(net107),
    .S(_0078_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1214_ (.A0(net554),
    .A1(net108),
    .S(_0858_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1215_ (.A0(net555),
    .A1(net109),
    .S(_0858_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1216_ (.A0(net556),
    .A1(net110),
    .S(_0858_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1217_ (.A0(net557),
    .A1(net111),
    .S(_0858_),
    .X(_0074_));
 sky130_fd_sc_hd__nand2_4 _1218_ (.A(net114),
    .B(net117),
    .Y(_0082_));
 sky130_fd_sc_hd__nand2_1 _1219_ (.A(_0611_),
    .B(_0615_),
    .Y(_0083_));
 sky130_fd_sc_hd__nor2_1 _1220_ (.A(_0613_),
    .B(_0609_),
    .Y(_0084_));
 sky130_fd_sc_hd__nor3_2 _1221_ (.A(_0082_),
    .B(_0083_),
    .C(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_1 _1222_ (.A(_0612_),
    .Y(_0086_));
 sky130_fd_sc_hd__a21oi_1 _1223_ (.A1(_0086_),
    .A2(_0613_),
    .B1(_0616_),
    .Y(_0087_));
 sky130_fd_sc_hd__nand2_1 _1224_ (.A(_0085_),
    .B(_0087_),
    .Y(_0088_));
 sky130_fd_sc_hd__nand2b_1 _1225_ (.A_N(net125),
    .B(_0612_),
    .Y(_0089_));
 sky130_fd_sc_hd__or3b_2 _1226_ (.A(_0611_),
    .B(net126),
    .C_N(_0613_),
    .X(_0090_));
 sky130_fd_sc_hd__a21o_1 _1227_ (.A1(_0744_),
    .A2(net126),
    .B1(_0612_),
    .X(_0091_));
 sky130_fd_sc_hd__o21a_1 _1228_ (.A1(_0616_),
    .A2(_0083_),
    .B1(_0091_),
    .X(_0092_));
 sky130_fd_sc_hd__o22ai_1 _1229_ (.A1(_0089_),
    .A2(_0090_),
    .B1(_0092_),
    .B2(_0613_),
    .Y(_0093_));
 sky130_fd_sc_hd__or3_2 _1230_ (.A(_0082_),
    .B(_0089_),
    .C(_0090_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_4 _1231_ (.A(instr_rdata_alu_i[12]),
    .X(_0095_));
 sky130_fd_sc_hd__nor2_1 _1232_ (.A(net115),
    .B(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__nor2_1 _1233_ (.A(_0094_),
    .B(_0096_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_2 _1234_ (.A(_0611_),
    .B(_0614_),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_2 _1235_ (.A(_0616_),
    .B(_0615_),
    .Y(_0099_));
 sky130_fd_sc_hd__o21ai_1 _1236_ (.A1(_0098_),
    .A2(_0099_),
    .B1(_0094_),
    .Y(_0100_));
 sky130_fd_sc_hd__o21ai_0 _1237_ (.A1(net116),
    .A2(_0097_),
    .B1(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__and4b_2 _1238_ (.A_N(_0082_),
    .B(_0088_),
    .C(_0093_),
    .D(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__clkinv_2 _1239_ (.A(net115),
    .Y(_0103_));
 sky130_fd_sc_hd__o21ai_2 _1240_ (.A1(_0103_),
    .A2(_0094_),
    .B1(_0622_),
    .Y(_0104_));
 sky130_fd_sc_hd__a21oi_4 _1241_ (.A1(_0100_),
    .A2(_0104_),
    .B1(net190),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2_8 _1242_ (.A(_0102_),
    .B(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__buf_16 _1243_ (.A(net190),
    .X(_0107_));
 sky130_fd_sc_hd__buf_6 _1244_ (.A(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__nor2_4 _1245_ (.A(_0086_),
    .B(_0616_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand2_1 _1246_ (.A(_0083_),
    .B(_0090_),
    .Y(_0110_));
 sky130_fd_sc_hd__nor2_1 _1247_ (.A(_0611_),
    .B(_0615_),
    .Y(_0111_));
 sky130_fd_sc_hd__nand2_1 _1248_ (.A(_0616_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__a21oi_1 _1249_ (.A1(_0091_),
    .A2(_0112_),
    .B1(_0613_),
    .Y(_0113_));
 sky130_fd_sc_hd__a21oi_2 _1250_ (.A1(_0109_),
    .A2(_0110_),
    .B1(_0113_),
    .Y(_0114_));
 sky130_fd_sc_hd__nor4b_4 _1251_ (.A(_0082_),
    .B(_0102_),
    .C(_0114_),
    .D_N(_0105_),
    .Y(_0115_));
 sky130_fd_sc_hd__buf_6 _1252_ (.A(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__nor4b_4 _1253_ (.A(_0107_),
    .B(_0098_),
    .C(_0099_),
    .D_N(_0104_),
    .Y(_0117_));
 sky130_fd_sc_hd__a222oi_1 _1254_ (.A1(_0108_),
    .A2(net191),
    .B1(_0116_),
    .B2(net226),
    .C1(_0117_),
    .C2(net148),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_1 _1255_ (.A(net293),
    .B(_0106_),
    .Y(_0119_));
 sky130_fd_sc_hd__a21oi_4 _1256_ (.A1(_0106_),
    .A2(_0118_),
    .B1(_0119_),
    .Y(net359));
 sky130_fd_sc_hd__clkbuf_4 _1257_ (.A(_0107_),
    .X(_0120_));
 sky130_fd_sc_hd__and2_0 _1258_ (.A(_0102_),
    .B(_0105_),
    .X(_0121_));
 sky130_fd_sc_hd__buf_6 _1259_ (.A(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_4 _1260_ (.A(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__buf_4 _1261_ (.A(_0115_),
    .X(_0124_));
 sky130_fd_sc_hd__a222oi_1 _1262_ (.A1(_0120_),
    .A2(net192),
    .B1(net294),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net227),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_1 _1263_ (.A(_0125_),
    .Y(net360));
 sky130_fd_sc_hd__a222oi_1 _1264_ (.A1(_0120_),
    .A2(net193),
    .B1(net295),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net228),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_1 _1265_ (.A(_0126_),
    .Y(net361));
 sky130_fd_sc_hd__a222oi_1 _1266_ (.A1(_0120_),
    .A2(net194),
    .B1(net296),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net229),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_1 _1267_ (.A(_0127_),
    .Y(net362));
 sky130_fd_sc_hd__a222oi_1 _1268_ (.A1(_0120_),
    .A2(net195),
    .B1(net297),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net230),
    .Y(_0128_));
 sky130_fd_sc_hd__clkinv_4 _1269_ (.A(_0128_),
    .Y(net363));
 sky130_fd_sc_hd__a222oi_1 _1270_ (.A1(_0120_),
    .A2(net196),
    .B1(net298),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net231),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1271_ (.A(_0129_),
    .Y(net364));
 sky130_fd_sc_hd__a222oi_1 _1272_ (.A1(_0120_),
    .A2(net197),
    .B1(net299),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net232),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_1 _1273_ (.A(_0130_),
    .Y(net365));
 sky130_fd_sc_hd__a222oi_1 _1274_ (.A1(_0120_),
    .A2(net198),
    .B1(net300),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net233),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_1 _1275_ (.A(_0131_),
    .Y(net366));
 sky130_fd_sc_hd__a222oi_1 _1276_ (.A1(_0120_),
    .A2(net199),
    .B1(net301),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net234),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_1 _1277_ (.A(_0132_),
    .Y(net367));
 sky130_fd_sc_hd__a222oi_1 _1278_ (.A1(_0120_),
    .A2(net200),
    .B1(net302),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net235),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_1 _1279_ (.A(_0133_),
    .Y(net368));
 sky130_fd_sc_hd__a222oi_1 _1280_ (.A1(_0120_),
    .A2(net201),
    .B1(net303),
    .B2(_0123_),
    .C1(_0124_),
    .C2(net236),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_1 _1281_ (.A(_0134_),
    .Y(net369));
 sky130_fd_sc_hd__a222oi_1 _1282_ (.A1(_0108_),
    .A2(net202),
    .B1(net237),
    .B2(_0116_),
    .C1(_0117_),
    .C2(net149),
    .Y(_0135_));
 sky130_fd_sc_hd__nor2_1 _1283_ (.A(net304),
    .B(_0106_),
    .Y(_0136_));
 sky130_fd_sc_hd__a21oi_4 _1284_ (.A1(_0106_),
    .A2(_0135_),
    .B1(_0136_),
    .Y(net370));
 sky130_fd_sc_hd__clkbuf_4 _1285_ (.A(_0107_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_4 _1286_ (.A(_0122_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_4 _1287_ (.A(_0115_),
    .X(_0139_));
 sky130_fd_sc_hd__a222oi_1 _1288_ (.A1(_0137_),
    .A2(net203),
    .B1(net305),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net238),
    .Y(_0140_));
 sky130_fd_sc_hd__clkinvlp_4 _1289_ (.A(_0140_),
    .Y(net371));
 sky130_fd_sc_hd__a222oi_1 _1290_ (.A1(_0137_),
    .A2(net204),
    .B1(net306),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net239),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_1 _1291_ (.A(_0141_),
    .Y(net372));
 sky130_fd_sc_hd__a222oi_1 _1292_ (.A1(_0137_),
    .A2(net205),
    .B1(net307),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net240),
    .Y(_0142_));
 sky130_fd_sc_hd__clkinv_4 _1293_ (.A(_0142_),
    .Y(net373));
 sky130_fd_sc_hd__a222oi_1 _1294_ (.A1(_0137_),
    .A2(net206),
    .B1(net308),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net241),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1295_ (.A(_0143_),
    .Y(net374));
 sky130_fd_sc_hd__a222oi_1 _1296_ (.A1(_0137_),
    .A2(net207),
    .B1(net309),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net242),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_1 _1297_ (.A(_0144_),
    .Y(net375));
 sky130_fd_sc_hd__a222oi_1 _1298_ (.A1(_0137_),
    .A2(net208),
    .B1(net310),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net243),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_1 _1299_ (.A(_0145_),
    .Y(net376));
 sky130_fd_sc_hd__a222oi_1 _1300_ (.A1(_0137_),
    .A2(net209),
    .B1(net311),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net244),
    .Y(_0146_));
 sky130_fd_sc_hd__clkinv_2 _1301_ (.A(_0146_),
    .Y(net377));
 sky130_fd_sc_hd__a222oi_1 _1302_ (.A1(_0137_),
    .A2(net210),
    .B1(net312),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net245),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1303_ (.A(_0147_),
    .Y(net378));
 sky130_fd_sc_hd__a222oi_1 _1304_ (.A1(_0137_),
    .A2(net211),
    .B1(net313),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net246),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1305_ (.A(_0148_),
    .Y(net379));
 sky130_fd_sc_hd__a222oi_1 _1306_ (.A1(_0137_),
    .A2(net212),
    .B1(net314),
    .B2(_0138_),
    .C1(_0139_),
    .C2(net247),
    .Y(_0149_));
 sky130_fd_sc_hd__clkinv_2 _1307_ (.A(_0149_),
    .Y(net380));
 sky130_fd_sc_hd__a222oi_1 _1308_ (.A1(_0107_),
    .A2(net213),
    .B1(net248),
    .B2(_0116_),
    .C1(_0117_),
    .C2(net150),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _1309_ (.A(net315),
    .B(_0106_),
    .Y(_0151_));
 sky130_fd_sc_hd__a21oi_4 _1310_ (.A1(_0106_),
    .A2(_0150_),
    .B1(_0151_),
    .Y(net381));
 sky130_fd_sc_hd__a222oi_1 _1311_ (.A1(_0108_),
    .A2(net214),
    .B1(net316),
    .B2(_0122_),
    .C1(_0116_),
    .C2(net249),
    .Y(_0152_));
 sky130_fd_sc_hd__clkinv_2 _1312_ (.A(_0152_),
    .Y(net382));
 sky130_fd_sc_hd__a222oi_1 _1313_ (.A1(_0108_),
    .A2(net215),
    .B1(net317),
    .B2(_0122_),
    .C1(_0116_),
    .C2(net250),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_4 _1314_ (.A(_0153_),
    .Y(net383));
 sky130_fd_sc_hd__a222oi_1 _1315_ (.A1(_0107_),
    .A2(net216),
    .B1(net251),
    .B2(_0115_),
    .C1(_0117_),
    .C2(net151),
    .Y(_0154_));
 sky130_fd_sc_hd__nor2_1 _1316_ (.A(net318),
    .B(_0106_),
    .Y(_0155_));
 sky130_fd_sc_hd__a21oi_4 _1317_ (.A1(_0106_),
    .A2(_0154_),
    .B1(_0155_),
    .Y(net384));
 sky130_fd_sc_hd__a222oi_1 _1318_ (.A1(_0107_),
    .A2(net217),
    .B1(net252),
    .B2(_0115_),
    .C1(_0117_),
    .C2(net152),
    .Y(_0156_));
 sky130_fd_sc_hd__nor2_1 _1319_ (.A(net319),
    .B(_0106_),
    .Y(_0157_));
 sky130_fd_sc_hd__a21oi_2 _1320_ (.A1(_0106_),
    .A2(_0156_),
    .B1(_0157_),
    .Y(net385));
 sky130_fd_sc_hd__a222oi_1 _1321_ (.A1(_0108_),
    .A2(net218),
    .B1(net320),
    .B2(_0122_),
    .C1(_0116_),
    .C2(net253),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_1 _1322_ (.A(_0158_),
    .Y(net386));
 sky130_fd_sc_hd__a222oi_1 _1323_ (.A1(_0108_),
    .A2(net219),
    .B1(net321),
    .B2(_0122_),
    .C1(_0116_),
    .C2(net254),
    .Y(_0159_));
 sky130_fd_sc_hd__clkinvlp_4 _1324_ (.A(_0159_),
    .Y(net387));
 sky130_fd_sc_hd__a222oi_1 _1325_ (.A1(_0108_),
    .A2(net220),
    .B1(net322),
    .B2(_0122_),
    .C1(_0116_),
    .C2(net255),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_1 _1326_ (.A(_0160_),
    .Y(net388));
 sky130_fd_sc_hd__a222oi_1 _1327_ (.A1(_0108_),
    .A2(net221),
    .B1(net323),
    .B2(_0122_),
    .C1(_0116_),
    .C2(net256),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_1 _1328_ (.A(_0161_),
    .Y(net389));
 sky130_fd_sc_hd__a222oi_1 _1329_ (.A1(_0108_),
    .A2(net222),
    .B1(net324),
    .B2(_0122_),
    .C1(_0116_),
    .C2(net257),
    .Y(_0162_));
 sky130_fd_sc_hd__clkinv_4 _1330_ (.A(_0162_),
    .Y(net390));
 sky130_fd_sc_hd__nor2b_2 _1331_ (.A(net125),
    .B_N(_0615_),
    .Y(_0163_));
 sky130_fd_sc_hd__a31oi_4 _1332_ (.A1(_0609_),
    .A2(_0746_),
    .A3(_0163_),
    .B1(net190),
    .Y(_0164_));
 sky130_fd_sc_hd__or3_1 _1333_ (.A(_0616_),
    .B(_0615_),
    .C(net116),
    .X(_0165_));
 sky130_fd_sc_hd__and4_1 _1334_ (.A(_0746_),
    .B(_0099_),
    .C(_0164_),
    .D(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__buf_8 _1335_ (.A(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__buf_6 _1336_ (.A(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__nor2_1 _1337_ (.A(_0613_),
    .B(_0082_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand3_4 _1338_ (.A(_0612_),
    .B(_0169_),
    .C(_0617_),
    .Y(_0170_));
 sky130_fd_sc_hd__nor2_1 _1339_ (.A(_0612_),
    .B(_0613_),
    .Y(_0171_));
 sky130_fd_sc_hd__nor2_1 _1340_ (.A(_0615_),
    .B(net116),
    .Y(_0172_));
 sky130_fd_sc_hd__a32o_1 _1341_ (.A1(_0612_),
    .A2(_0615_),
    .A3(_0609_),
    .B1(_0171_),
    .B2(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__nor3_2 _1342_ (.A(_0616_),
    .B(_0744_),
    .C(_0082_),
    .Y(_0174_));
 sky130_fd_sc_hd__or3b_1 _1343_ (.A(net115),
    .B(net116),
    .C_N(_0095_),
    .X(_0175_));
 sky130_fd_sc_hd__nor4_4 _1344_ (.A(_0082_),
    .B(_0089_),
    .C(_0090_),
    .D(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__a21oi_1 _1345_ (.A1(_0173_),
    .A2(_0174_),
    .B1(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__a21oi_4 _1346_ (.A1(_0170_),
    .A2(_0177_),
    .B1(net190),
    .Y(_0178_));
 sky130_fd_sc_hd__mux2i_2 _1347_ (.A0(_0689_),
    .A1(net168),
    .S(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__a211o_4 _1348_ (.A1(_0085_),
    .A2(_0109_),
    .B1(_0176_),
    .C1(net190),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_4 _1349_ (.A(_0164_),
    .B(_0170_),
    .Y(_0181_));
 sky130_fd_sc_hd__clkbuf_4 _1350_ (.A(_0167_),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(net325),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__o41ai_4 _1352_ (.A1(_0168_),
    .A2(_0179_),
    .A3(_0180_),
    .A4(_0181_),
    .B1(_0183_),
    .Y(net391));
 sky130_fd_sc_hd__clkbuf_8 _1353_ (.A(_0167_),
    .X(_0184_));
 sky130_fd_sc_hd__nor2_1 _1354_ (.A(_0178_),
    .B(_0181_),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_1 _1355_ (.A(net190),
    .Y(_0186_));
 sky130_fd_sc_hd__a21o_2 _1356_ (.A1(_0173_),
    .A2(_0174_),
    .B1(_0176_),
    .X(_0187_));
 sky130_fd_sc_hd__nand3_1 _1357_ (.A(_0186_),
    .B(_0170_),
    .C(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__a21oi_4 _1358_ (.A1(_0164_),
    .A2(_0188_),
    .B1(_0180_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _1359_ (.A(_0185_),
    .B(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__nor3_4 _1360_ (.A(_0107_),
    .B(_0167_),
    .C(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__a22o_2 _1361_ (.A1(net326),
    .A2(_0184_),
    .B1(_0191_),
    .B2(_0645_),
    .X(net392));
 sky130_fd_sc_hd__buf_6 _1362_ (.A(_0167_),
    .X(_0192_));
 sky130_fd_sc_hd__a211oi_4 _1363_ (.A1(_0085_),
    .A2(_0109_),
    .B1(_0176_),
    .C1(_0107_),
    .Y(_0193_));
 sky130_fd_sc_hd__and2_1 _1364_ (.A(_0164_),
    .B(_0170_),
    .X(_0194_));
 sky130_fd_sc_hd__nand3_1 _1365_ (.A(net168),
    .B(_0193_),
    .C(_0181_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand3_1 _1366_ (.A(_0689_),
    .B(_0180_),
    .C(_0194_),
    .Y(_0196_));
 sky130_fd_sc_hd__a21oi_1 _1367_ (.A1(_0195_),
    .A2(_0196_),
    .B1(_0178_),
    .Y(_0197_));
 sky130_fd_sc_hd__a31oi_2 _1368_ (.A1(_0641_),
    .A2(_0193_),
    .A3(_0194_),
    .B1(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(net327),
    .B(_0182_),
    .Y(_0199_));
 sky130_fd_sc_hd__o21ai_4 _1370_ (.A1(_0192_),
    .A2(_0198_),
    .B1(_0199_),
    .Y(net393));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(_0180_),
    .B(_0194_),
    .Y(_0200_));
 sky130_fd_sc_hd__and2_1 _1372_ (.A(_0178_),
    .B(_0181_),
    .X(_0201_));
 sky130_fd_sc_hd__o21bai_4 _1373_ (.A1(_0178_),
    .A2(_0200_),
    .B1_N(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _1374_ (.A(_0641_),
    .B(_0193_),
    .Y(_0203_));
 sky130_fd_sc_hd__nor2_2 _1375_ (.A(_0203_),
    .B(_0201_),
    .Y(_0204_));
 sky130_fd_sc_hd__a21oi_1 _1376_ (.A1(_0660_),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__nand2_1 _1377_ (.A(net328),
    .B(_0182_),
    .Y(_0206_));
 sky130_fd_sc_hd__o21ai_2 _1378_ (.A1(_0192_),
    .A2(_0205_),
    .B1(_0206_),
    .Y(net394));
 sky130_fd_sc_hd__a21oi_1 _1379_ (.A1(_0659_),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _1380_ (.A(net329),
    .B(_0182_),
    .Y(_0208_));
 sky130_fd_sc_hd__o21ai_2 _1381_ (.A1(_0192_),
    .A2(_0207_),
    .B1(_0208_),
    .Y(net395));
 sky130_fd_sc_hd__a21oi_1 _1382_ (.A1(_0633_),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0209_));
 sky130_fd_sc_hd__nand2_1 _1383_ (.A(net330),
    .B(_0182_),
    .Y(_0210_));
 sky130_fd_sc_hd__o21ai_1 _1384_ (.A1(_0192_),
    .A2(_0209_),
    .B1(_0210_),
    .Y(net396));
 sky130_fd_sc_hd__a21oi_1 _1385_ (.A1(net148),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _1386_ (.A(net331),
    .B(_0182_),
    .Y(_0212_));
 sky130_fd_sc_hd__o21ai_2 _1387_ (.A1(_0192_),
    .A2(_0211_),
    .B1(_0212_),
    .Y(net397));
 sky130_fd_sc_hd__a21oi_1 _1388_ (.A1(net149),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0213_));
 sky130_fd_sc_hd__nand2_1 _1389_ (.A(net332),
    .B(_0182_),
    .Y(_0214_));
 sky130_fd_sc_hd__o21ai_1 _1390_ (.A1(_0192_),
    .A2(_0213_),
    .B1(_0214_),
    .Y(net398));
 sky130_fd_sc_hd__a21oi_1 _1391_ (.A1(net150),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0215_));
 sky130_fd_sc_hd__nand2_1 _1392_ (.A(net333),
    .B(_0182_),
    .Y(_0216_));
 sky130_fd_sc_hd__o21ai_4 _1393_ (.A1(_0192_),
    .A2(_0215_),
    .B1(_0216_),
    .Y(net399));
 sky130_fd_sc_hd__a21oi_1 _1394_ (.A1(net151),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _1395_ (.A(net334),
    .B(_0182_),
    .Y(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1396_ (.A1(_0192_),
    .A2(_0217_),
    .B1(_0218_),
    .Y(net400));
 sky130_fd_sc_hd__a21oi_1 _1397_ (.A1(net152),
    .A2(_0202_),
    .B1(_0204_),
    .Y(_0219_));
 sky130_fd_sc_hd__clkbuf_4 _1398_ (.A(_0167_),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _1399_ (.A(net335),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__o21ai_1 _1400_ (.A1(_0192_),
    .A2(_0219_),
    .B1(_0221_),
    .Y(net401));
 sky130_fd_sc_hd__nand2b_1 _1401_ (.A_N(_0178_),
    .B(net155),
    .Y(_0222_));
 sky130_fd_sc_hd__buf_6 _1402_ (.A(net113),
    .X(_0223_));
 sky130_fd_sc_hd__nand3_1 _1403_ (.A(_0223_),
    .B(_0178_),
    .C(_0180_),
    .Y(_0224_));
 sky130_fd_sc_hd__a21oi_1 _1404_ (.A1(_0222_),
    .A2(_0224_),
    .B1(_0181_),
    .Y(_0225_));
 sky130_fd_sc_hd__a21oi_2 _1405_ (.A1(net169),
    .A2(_0189_),
    .B1(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _1406_ (.A(net336),
    .B(_0220_),
    .Y(_0227_));
 sky130_fd_sc_hd__o21ai_1 _1407_ (.A1(_0192_),
    .A2(_0226_),
    .B1(_0227_),
    .Y(net402));
 sky130_fd_sc_hd__clkbuf_4 _1408_ (.A(_0201_),
    .X(_0228_));
 sky130_fd_sc_hd__o21a_2 _1409_ (.A1(_0185_),
    .A2(_0189_),
    .B1(_0641_),
    .X(_0229_));
 sky130_fd_sc_hd__a21oi_1 _1410_ (.A1(_0689_),
    .A2(_0228_),
    .B1(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _1411_ (.A(net337),
    .B(_0220_),
    .Y(_0231_));
 sky130_fd_sc_hd__o21ai_2 _1412_ (.A1(_0184_),
    .A2(_0230_),
    .B1(_0231_),
    .Y(net403));
 sky130_fd_sc_hd__a21oi_1 _1413_ (.A1(net155),
    .A2(_0228_),
    .B1(_0229_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _1414_ (.A(net338),
    .B(_0220_),
    .Y(_0233_));
 sky130_fd_sc_hd__o21ai_2 _1415_ (.A1(_0184_),
    .A2(_0232_),
    .B1(_0233_),
    .Y(net404));
 sky130_fd_sc_hd__a21oi_1 _1416_ (.A1(net156),
    .A2(_0228_),
    .B1(_0229_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _1417_ (.A(net339),
    .B(_0220_),
    .Y(_0235_));
 sky130_fd_sc_hd__o21ai_2 _1418_ (.A1(_0184_),
    .A2(_0234_),
    .B1(_0235_),
    .Y(net405));
 sky130_fd_sc_hd__a21oi_1 _1419_ (.A1(net157),
    .A2(_0228_),
    .B1(_0229_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _1420_ (.A(net340),
    .B(_0220_),
    .Y(_0237_));
 sky130_fd_sc_hd__o21ai_4 _1421_ (.A1(_0184_),
    .A2(_0236_),
    .B1(_0237_),
    .Y(net406));
 sky130_fd_sc_hd__a21oi_1 _1422_ (.A1(net158),
    .A2(_0228_),
    .B1(_0229_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _1423_ (.A(net341),
    .B(_0220_),
    .Y(_0239_));
 sky130_fd_sc_hd__o21ai_2 _1424_ (.A1(_0184_),
    .A2(_0238_),
    .B1(_0239_),
    .Y(net407));
 sky130_fd_sc_hd__nor3b_4 _1425_ (.A(_0107_),
    .B(_0167_),
    .C_N(_0229_),
    .Y(_0240_));
 sky130_fd_sc_hd__a221o_1 _1426_ (.A1(net342),
    .A2(_0168_),
    .B1(_0228_),
    .B2(_0646_),
    .C1(_0240_),
    .X(net408));
 sky130_fd_sc_hd__a221o_1 _1427_ (.A1(net343),
    .A2(_0168_),
    .B1(_0228_),
    .B2(net159),
    .C1(_0240_),
    .X(net409));
 sky130_fd_sc_hd__a221o_2 _1428_ (.A1(net344),
    .A2(_0168_),
    .B1(_0228_),
    .B2(net160),
    .C1(_0240_),
    .X(net410));
 sky130_fd_sc_hd__a221o_2 _1429_ (.A1(net345),
    .A2(_0168_),
    .B1(_0228_),
    .B2(net161),
    .C1(_0240_),
    .X(net411));
 sky130_fd_sc_hd__a221o_2 _1430_ (.A1(net346),
    .A2(_0167_),
    .B1(_0228_),
    .B2(net162),
    .C1(_0240_),
    .X(net412));
 sky130_fd_sc_hd__inv_1 _1431_ (.A(net347),
    .Y(_0241_));
 sky130_fd_sc_hd__nand2b_1 _1432_ (.A_N(_0178_),
    .B(net156),
    .Y(_0242_));
 sky130_fd_sc_hd__nand3b_1 _1433_ (.A_N(_0223_),
    .B(_0178_),
    .C(_0180_),
    .Y(_0243_));
 sky130_fd_sc_hd__a21oi_1 _1434_ (.A1(_0242_),
    .A2(_0243_),
    .B1(_0181_),
    .Y(_0244_));
 sky130_fd_sc_hd__a2111oi_1 _1435_ (.A1(net170),
    .A2(_0189_),
    .B1(_0244_),
    .C1(_0108_),
    .D1(_0168_),
    .Y(_0245_));
 sky130_fd_sc_hd__a21oi_2 _1436_ (.A1(_0241_),
    .A2(_0182_),
    .B1(_0245_),
    .Y(net413));
 sky130_fd_sc_hd__a221o_1 _1437_ (.A1(net348),
    .A2(_0167_),
    .B1(_0201_),
    .B2(_0645_),
    .C1(_0240_),
    .X(net414));
 sky130_fd_sc_hd__nand2_1 _1438_ (.A(_0178_),
    .B(_0180_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand3_1 _1439_ (.A(_0641_),
    .B(_0186_),
    .C(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_1 _1440_ (.A(net349),
    .B(_0220_),
    .Y(_0248_));
 sky130_fd_sc_hd__o21ai_1 _1441_ (.A1(_0184_),
    .A2(_0247_),
    .B1(_0248_),
    .Y(net415));
 sky130_fd_sc_hd__a22oi_1 _1442_ (.A1(net157),
    .A2(_0185_),
    .B1(_0189_),
    .B2(net144),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _1443_ (.A(net350),
    .B(_0220_),
    .Y(_0250_));
 sky130_fd_sc_hd__o21ai_2 _1444_ (.A1(_0184_),
    .A2(_0249_),
    .B1(_0250_),
    .Y(net416));
 sky130_fd_sc_hd__a22oi_1 _1445_ (.A1(net158),
    .A2(_0185_),
    .B1(_0189_),
    .B2(net145),
    .Y(_0251_));
 sky130_fd_sc_hd__nand2_1 _1446_ (.A(net351),
    .B(_0220_),
    .Y(_0252_));
 sky130_fd_sc_hd__o21ai_1 _1447_ (.A1(_0184_),
    .A2(_0251_),
    .B1(_0252_),
    .Y(net417));
 sky130_fd_sc_hd__a22o_1 _1448_ (.A1(net352),
    .A2(_0184_),
    .B1(_0191_),
    .B2(_0646_),
    .X(net418));
 sky130_fd_sc_hd__a22o_4 _1449_ (.A1(net353),
    .A2(_0168_),
    .B1(_0191_),
    .B2(net159),
    .X(net419));
 sky130_fd_sc_hd__a22o_2 _1450_ (.A1(net354),
    .A2(_0168_),
    .B1(_0191_),
    .B2(net160),
    .X(net420));
 sky130_fd_sc_hd__a22o_1 _1451_ (.A1(net355),
    .A2(_0168_),
    .B1(_0191_),
    .B2(net161),
    .X(net421));
 sky130_fd_sc_hd__a22o_1 _1452_ (.A1(net356),
    .A2(_0168_),
    .B1(_0191_),
    .B2(net162),
    .X(net422));
 sky130_fd_sc_hd__buf_4 _1453_ (.A(net115),
    .X(_0253_));
 sky130_fd_sc_hd__nor2_1 _1454_ (.A(_0095_),
    .B(net118),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _1455_ (.A(_0095_),
    .Y(_0255_));
 sky130_fd_sc_hd__nor3_1 _1456_ (.A(net118),
    .B(net119),
    .C(_0619_),
    .Y(_0256_));
 sky130_fd_sc_hd__and2_1 _1457_ (.A(net123),
    .B(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__nand3_1 _1458_ (.A(_0255_),
    .B(_0622_),
    .C(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__nand4b_1 _1459_ (.A_N(net118),
    .B(_0620_),
    .C(_0095_),
    .D(_0610_),
    .Y(_0259_));
 sky130_fd_sc_hd__a21oi_1 _1460_ (.A1(_0258_),
    .A2(_0259_),
    .B1(_0253_),
    .Y(_0260_));
 sky130_fd_sc_hd__a31oi_2 _1461_ (.A1(_0253_),
    .A2(_0620_),
    .A3(_0254_),
    .B1(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__or3_1 _1462_ (.A(_0745_),
    .B(_0619_),
    .C(_0112_),
    .X(_0262_));
 sky130_fd_sc_hd__nand3_4 _1463_ (.A(net558),
    .B(_0746_),
    .C(_0163_),
    .Y(_0263_));
 sky130_fd_sc_hd__o31a_1 _1464_ (.A1(_0255_),
    .A2(net123),
    .A3(_0262_),
    .B1(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_2 _1465_ (.A(_0745_),
    .B(_0112_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor2_1 _1466_ (.A(_0253_),
    .B(_0263_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21oi_1 _1467_ (.A1(_0253_),
    .A2(_0265_),
    .B1(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__o32a_2 _1468_ (.A1(_0253_),
    .A2(_0622_),
    .A3(_0264_),
    .B1(_0267_),
    .B2(_0095_),
    .X(_0268_));
 sky130_fd_sc_hd__o31ai_4 _1469_ (.A1(net119),
    .A2(_0618_),
    .A3(_0261_),
    .B1(_0268_),
    .Y(net423));
 sky130_fd_sc_hd__nand2_1 _1470_ (.A(_0255_),
    .B(_0610_),
    .Y(_0269_));
 sky130_fd_sc_hd__a21oi_1 _1471_ (.A1(_0253_),
    .A2(_0269_),
    .B1(_0096_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(_0095_),
    .B(_0622_),
    .Y(_0271_));
 sky130_fd_sc_hd__and2_1 _1473_ (.A(_0269_),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2b_1 _1474_ (.A_N(_0272_),
    .B(_0265_),
    .Y(_0273_));
 sky130_fd_sc_hd__nor2_2 _1475_ (.A(_0745_),
    .B(_0756_),
    .Y(_0274_));
 sky130_fd_sc_hd__and3_1 _1476_ (.A(_0103_),
    .B(net123),
    .C(_0256_),
    .X(_0275_));
 sky130_fd_sc_hd__o21ai_1 _1477_ (.A1(_0620_),
    .A2(_0275_),
    .B1(_0272_),
    .Y(_0276_));
 sky130_fd_sc_hd__a22oi_1 _1478_ (.A1(_0611_),
    .A2(_0171_),
    .B1(_0110_),
    .B2(_0612_),
    .Y(_0277_));
 sky130_fd_sc_hd__o32a_1 _1479_ (.A1(_0613_),
    .A2(_0615_),
    .A3(_0109_),
    .B1(_0277_),
    .B2(_0616_),
    .X(_0278_));
 sky130_fd_sc_hd__nand4_1 _1480_ (.A(_0103_),
    .B(_0095_),
    .C(_0619_),
    .D(_0265_),
    .Y(_0279_));
 sky130_fd_sc_hd__nor2_2 _1481_ (.A(net115),
    .B(net116),
    .Y(_0280_));
 sky130_fd_sc_hd__a21oi_1 _1482_ (.A1(_0094_),
    .A2(_0279_),
    .B1(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__or3_2 _1483_ (.A(_0082_),
    .B(_0278_),
    .C(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__a31oi_4 _1484_ (.A1(_0274_),
    .A2(_0621_),
    .A3(_0276_),
    .B1(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__o211ai_4 _1485_ (.A1(_0263_),
    .A2(_0270_),
    .B1(_0273_),
    .C1(_0283_),
    .Y(net424));
 sky130_fd_sc_hd__and3_1 _1486_ (.A(net558),
    .B(_0746_),
    .C(_0163_),
    .X(_0284_));
 sky130_fd_sc_hd__a21oi_1 _1487_ (.A1(net115),
    .A2(_0284_),
    .B1(_0269_),
    .Y(_0285_));
 sky130_fd_sc_hd__nor2_2 _1488_ (.A(_0284_),
    .B(_0265_),
    .Y(_0286_));
 sky130_fd_sc_hd__a21oi_1 _1489_ (.A1(_0284_),
    .A2(_0271_),
    .B1(net115),
    .Y(_0287_));
 sky130_fd_sc_hd__nor3_1 _1490_ (.A(_0285_),
    .B(_0286_),
    .C(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _1491_ (.A(_0274_),
    .B(_0621_),
    .Y(_0289_));
 sky130_fd_sc_hd__a22oi_1 _1492_ (.A1(_0610_),
    .A2(_0620_),
    .B1(_0257_),
    .B2(_0280_),
    .Y(_0290_));
 sky130_fd_sc_hd__a31oi_1 _1493_ (.A1(_0095_),
    .A2(_0610_),
    .A3(_0257_),
    .B1(_0620_),
    .Y(_0291_));
 sky130_fd_sc_hd__o22ai_1 _1494_ (.A1(_0095_),
    .A2(_0290_),
    .B1(_0291_),
    .B2(_0253_),
    .Y(_0292_));
 sky130_fd_sc_hd__nor2_1 _1495_ (.A(_0289_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__or3_4 _1496_ (.A(_0282_),
    .B(_0288_),
    .C(_0293_),
    .X(net425));
 sky130_fd_sc_hd__nand2_1 _1497_ (.A(_0622_),
    .B(net123),
    .Y(_0294_));
 sky130_fd_sc_hd__a21oi_1 _1498_ (.A1(_0610_),
    .A2(_0262_),
    .B1(_0286_),
    .Y(_0295_));
 sky130_fd_sc_hd__a31oi_2 _1499_ (.A1(_0274_),
    .A2(_0256_),
    .A3(_0294_),
    .B1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__nor3_4 _1500_ (.A(_0253_),
    .B(_0255_),
    .C(_0296_),
    .Y(net426));
 sky130_fd_sc_hd__a21oi_4 _1501_ (.A1(_0253_),
    .A2(_0622_),
    .B1(_0263_),
    .Y(net427));
 sky130_fd_sc_hd__o21ai_0 _1502_ (.A1(_0610_),
    .A2(net118),
    .B1(_0620_),
    .Y(_0297_));
 sky130_fd_sc_hd__a21oi_1 _1503_ (.A1(_0257_),
    .A2(_0272_),
    .B1(_0620_),
    .Y(_0298_));
 sky130_fd_sc_hd__a21oi_1 _1504_ (.A1(_0253_),
    .A2(_0297_),
    .B1(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__nor2_1 _1505_ (.A(_0618_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__nor2_1 _1506_ (.A(_0282_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__o31ai_4 _1507_ (.A1(_0103_),
    .A2(_0610_),
    .A3(_0286_),
    .B1(_0301_),
    .Y(net428));
 sky130_fd_sc_hd__nand3_4 _1508_ (.A(_0753_),
    .B(_0759_),
    .C(_0853_),
    .Y(_0302_));
 sky130_fd_sc_hd__nor3_1 _1509_ (.A(_0750_),
    .B(_0763_),
    .C(_0302_),
    .Y(branch_set_d));
 sky130_fd_sc_hd__nand2_8 _1510_ (.A(_0707_),
    .B(_0807_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_4 _1511_ (.A(_0608_),
    .B(_0717_),
    .Y(_0304_));
 sky130_fd_sc_hd__nor2_1 _1512_ (.A(net226),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21ai_1 _1513_ (.A1(\controller_i.store_err_q ),
    .A2(\controller_i.load_err_q ),
    .B1(_0811_),
    .Y(_0306_));
 sky130_fd_sc_hd__a21oi_4 _1514_ (.A1(_0720_),
    .A2(_0715_),
    .B1(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__buf_6 _1515_ (.A(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(net143),
    .A1(net127),
    .S(_0223_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_8 _1517_ (.A(\controller_i.illegal_insn_q ),
    .X(_0310_));
 sky130_fd_sc_hd__buf_8 _1518_ (.A(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _1519_ (.A(_0608_),
    .B(_0717_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_8 _1520_ (.A(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__a221oi_1 _1521_ (.A1(net191),
    .A2(_0308_),
    .B1(_0309_),
    .B2(_0311_),
    .C1(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__nor3_2 _1522_ (.A(_0303_),
    .B(_0305_),
    .C(_0314_),
    .Y(net430));
 sky130_fd_sc_hd__buf_8 _1523_ (.A(_0312_),
    .X(_0315_));
 sky130_fd_sc_hd__buf_4 _1524_ (.A(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__inv_1 _1525_ (.A(net254),
    .Y(_0317_));
 sky130_fd_sc_hd__nand4_4 _1526_ (.A(net112),
    .B(net237),
    .C(net248),
    .D(net251),
    .Y(_0318_));
 sky130_fd_sc_hd__nand2_1 _1527_ (.A(net252),
    .B(net253),
    .Y(_0319_));
 sky130_fd_sc_hd__nor3_4 _1528_ (.A(_0317_),
    .B(_0318_),
    .C(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__nand4_1 _1529_ (.A(net255),
    .B(net256),
    .C(net257),
    .D(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__xor2_1 _1530_ (.A(net227),
    .B(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1531_ (.A0(net144),
    .A1(net128),
    .S(_0223_),
    .X(_0323_));
 sky130_fd_sc_hd__a221oi_1 _1532_ (.A1(net192),
    .A2(_0308_),
    .B1(_0323_),
    .B2(_0311_),
    .C1(_0313_),
    .Y(_0324_));
 sky130_fd_sc_hd__buf_4 _1533_ (.A(_0303_),
    .X(_0325_));
 sky130_fd_sc_hd__a211oi_2 _1534_ (.A1(_0316_),
    .A2(_0322_),
    .B1(_0324_),
    .C1(_0325_),
    .Y(net431));
 sky130_fd_sc_hd__nand4_4 _1535_ (.A(net112),
    .B(net251),
    .C(_0863_),
    .D(net252),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_1 _1536_ (.A(net253),
    .B(net254),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_4 _1537_ (.A(_0326_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__and4_2 _1538_ (.A(net255),
    .B(net256),
    .C(net257),
    .D(net227),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_2 _1539_ (.A(_0328_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xor2_1 _1540_ (.A(net228),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__buf_6 _1541_ (.A(net113),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(net145),
    .A1(net129),
    .S(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__a221oi_1 _1543_ (.A1(net193),
    .A2(_0308_),
    .B1(_0333_),
    .B2(_0311_),
    .C1(_0313_),
    .Y(_0334_));
 sky130_fd_sc_hd__a211oi_1 _1544_ (.A1(_0316_),
    .A2(_0331_),
    .B1(_0334_),
    .C1(_0325_),
    .Y(net432));
 sky130_fd_sc_hd__nand3_1 _1545_ (.A(net228),
    .B(_0320_),
    .C(_0329_),
    .Y(_0335_));
 sky130_fd_sc_hd__xor2_1 _1546_ (.A(net229),
    .B(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _1547_ (.A0(_0660_),
    .A1(net130),
    .S(_0332_),
    .X(_0337_));
 sky130_fd_sc_hd__a221oi_1 _1548_ (.A1(net194),
    .A2(_0308_),
    .B1(_0337_),
    .B2(_0311_),
    .C1(_0313_),
    .Y(_0338_));
 sky130_fd_sc_hd__a211oi_1 _1549_ (.A1(_0316_),
    .A2(_0336_),
    .B1(_0338_),
    .C1(_0325_),
    .Y(net433));
 sky130_fd_sc_hd__nand2_1 _1550_ (.A(net228),
    .B(net229),
    .Y(_0339_));
 sky130_fd_sc_hd__nor2_1 _1551_ (.A(_0330_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__xnor2_1 _1552_ (.A(net230),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__mux2_1 _1553_ (.A0(_0659_),
    .A1(net131),
    .S(_0332_),
    .X(_0342_));
 sky130_fd_sc_hd__a221oi_1 _1554_ (.A1(net195),
    .A2(_0308_),
    .B1(_0342_),
    .B2(_0311_),
    .C1(_0313_),
    .Y(_0343_));
 sky130_fd_sc_hd__a211oi_1 _1555_ (.A1(_0316_),
    .A2(_0341_),
    .B1(_0343_),
    .C1(_0325_),
    .Y(net434));
 sky130_fd_sc_hd__nand2_2 _1556_ (.A(_0320_),
    .B(_0329_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand3_1 _1557_ (.A(net228),
    .B(net229),
    .C(net230),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_1 _1558_ (.A(_0344_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__xnor2_1 _1559_ (.A(net231),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _1560_ (.A(_0223_),
    .B(net132),
    .Y(_0348_));
 sky130_fd_sc_hd__o21ai_2 _1561_ (.A1(_0644_),
    .A2(_0223_),
    .B1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__a221oi_2 _1562_ (.A1(net196),
    .A2(_0308_),
    .B1(_0349_),
    .B2(_0311_),
    .C1(_0313_),
    .Y(_0350_));
 sky130_fd_sc_hd__a211oi_4 _1563_ (.A1(_0316_),
    .A2(_0347_),
    .B1(_0350_),
    .C1(_0325_),
    .Y(net435));
 sky130_fd_sc_hd__and4_1 _1564_ (.A(net228),
    .B(net229),
    .C(net230),
    .D(net231),
    .X(_0351_));
 sky130_fd_sc_hd__nand3_1 _1565_ (.A(_0328_),
    .B(_0329_),
    .C(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__xor2_1 _1566_ (.A(net232),
    .B(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(net148),
    .A1(net133),
    .S(_0332_),
    .X(_0354_));
 sky130_fd_sc_hd__a221oi_1 _1568_ (.A1(net197),
    .A2(_0308_),
    .B1(_0354_),
    .B2(_0311_),
    .C1(_0313_),
    .Y(_0355_));
 sky130_fd_sc_hd__a211oi_1 _1569_ (.A1(_0316_),
    .A2(_0353_),
    .B1(_0355_),
    .C1(_0325_),
    .Y(net436));
 sky130_fd_sc_hd__nand2_1 _1570_ (.A(net232),
    .B(_0351_),
    .Y(_0356_));
 sky130_fd_sc_hd__nor2_1 _1571_ (.A(_0344_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__xnor2_1 _1572_ (.A(net233),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2b_1 _1573_ (.A(net113),
    .B_N(_0310_),
    .Y(_0359_));
 sky130_fd_sc_hd__buf_4 _1574_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_4 _1575_ (.A(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__a221oi_1 _1576_ (.A1(net198),
    .A2(_0308_),
    .B1(_0361_),
    .B2(net149),
    .C1(_0313_),
    .Y(_0362_));
 sky130_fd_sc_hd__a211oi_2 _1577_ (.A1(_0316_),
    .A2(_0358_),
    .B1(_0362_),
    .C1(_0325_),
    .Y(net437));
 sky130_fd_sc_hd__nand3_1 _1578_ (.A(net232),
    .B(net233),
    .C(_0351_),
    .Y(_0363_));
 sky130_fd_sc_hd__nor2_1 _1579_ (.A(_0330_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__xnor2_1 _1580_ (.A(net234),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2b_1 _1581_ (.A(_0310_),
    .B_N(net199),
    .Y(_0366_));
 sky130_fd_sc_hd__buf_4 _1582_ (.A(_0315_),
    .X(_0367_));
 sky130_fd_sc_hd__a221oi_1 _1583_ (.A1(net150),
    .A2(_0360_),
    .B1(_0366_),
    .B2(_0308_),
    .C1(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__a211oi_2 _1584_ (.A1(_0316_),
    .A2(_0365_),
    .B1(_0368_),
    .C1(_0325_),
    .Y(net438));
 sky130_fd_sc_hd__nand4_1 _1585_ (.A(net232),
    .B(net233),
    .C(net234),
    .D(_0351_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _1586_ (.A(_0344_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__xnor2_1 _1587_ (.A(net235),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__buf_4 _1588_ (.A(_0307_),
    .X(_0372_));
 sky130_fd_sc_hd__a221oi_1 _1589_ (.A1(net200),
    .A2(_0372_),
    .B1(_0361_),
    .B2(net151),
    .C1(_0367_),
    .Y(_0373_));
 sky130_fd_sc_hd__a211oi_2 _1590_ (.A1(_0316_),
    .A2(_0371_),
    .B1(_0373_),
    .C1(_0325_),
    .Y(net439));
 sky130_fd_sc_hd__inv_1 _1591_ (.A(net235),
    .Y(_0374_));
 sky130_fd_sc_hd__or2_2 _1592_ (.A(_0374_),
    .B(_0369_),
    .X(_0375_));
 sky130_fd_sc_hd__nor2_4 _1593_ (.A(_0330_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__xnor2_1 _1594_ (.A(net236),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__a221oi_1 _1595_ (.A1(net201),
    .A2(_0372_),
    .B1(_0361_),
    .B2(net152),
    .C1(_0367_),
    .Y(_0378_));
 sky130_fd_sc_hd__a211oi_2 _1596_ (.A1(_0316_),
    .A2(_0377_),
    .B1(_0378_),
    .C1(_0325_),
    .Y(net440));
 sky130_fd_sc_hd__buf_6 _1597_ (.A(_0315_),
    .X(_0379_));
 sky130_fd_sc_hd__xnor2_1 _1598_ (.A(net112),
    .B(net237),
    .Y(_0380_));
 sky130_fd_sc_hd__mux2_1 _1599_ (.A0(net153),
    .A1(net134),
    .S(_0332_),
    .X(_0381_));
 sky130_fd_sc_hd__a221oi_2 _1600_ (.A1(net202),
    .A2(_0372_),
    .B1(_0381_),
    .B2(_0311_),
    .C1(_0367_),
    .Y(_0382_));
 sky130_fd_sc_hd__buf_6 _1601_ (.A(_0303_),
    .X(_0383_));
 sky130_fd_sc_hd__a211oi_2 _1602_ (.A1(_0379_),
    .A2(_0380_),
    .B1(_0382_),
    .C1(_0383_),
    .Y(net441));
 sky130_fd_sc_hd__nor2_4 _1603_ (.A(_0344_),
    .B(_0375_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_1 _1604_ (.A(net236),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__xor2_1 _1605_ (.A(net238),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a221oi_1 _1606_ (.A1(net203),
    .A2(_0372_),
    .B1(_0361_),
    .B2(_0689_),
    .C1(_0367_),
    .Y(_0387_));
 sky130_fd_sc_hd__a211oi_1 _1607_ (.A1(_0379_),
    .A2(_0386_),
    .B1(_0387_),
    .C1(_0383_),
    .Y(net442));
 sky130_fd_sc_hd__nand3_1 _1608_ (.A(net236),
    .B(net238),
    .C(_0376_),
    .Y(_0388_));
 sky130_fd_sc_hd__xor2_1 _1609_ (.A(net239),
    .B(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__a221oi_2 _1610_ (.A1(net204),
    .A2(_0372_),
    .B1(_0361_),
    .B2(net155),
    .C1(_0367_),
    .Y(_0390_));
 sky130_fd_sc_hd__a211oi_4 _1611_ (.A1(_0379_),
    .A2(_0389_),
    .B1(_0390_),
    .C1(_0383_),
    .Y(net443));
 sky130_fd_sc_hd__nand4_1 _1612_ (.A(net236),
    .B(net238),
    .C(net239),
    .D(_0384_),
    .Y(_0391_));
 sky130_fd_sc_hd__xor2_1 _1613_ (.A(net240),
    .B(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__a221oi_1 _1614_ (.A1(net205),
    .A2(_0372_),
    .B1(_0361_),
    .B2(net156),
    .C1(_0367_),
    .Y(_0393_));
 sky130_fd_sc_hd__a211oi_2 _1615_ (.A1(_0379_),
    .A2(_0392_),
    .B1(_0393_),
    .C1(_0383_),
    .Y(net444));
 sky130_fd_sc_hd__and4_2 _1616_ (.A(net236),
    .B(net238),
    .C(net239),
    .D(net240),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _1617_ (.A(_0376_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__xor2_1 _1618_ (.A(net241),
    .B(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__a221oi_2 _1619_ (.A1(net206),
    .A2(_0372_),
    .B1(_0361_),
    .B2(net157),
    .C1(_0367_),
    .Y(_0397_));
 sky130_fd_sc_hd__a211oi_2 _1620_ (.A1(_0379_),
    .A2(_0396_),
    .B1(_0397_),
    .C1(_0383_),
    .Y(net445));
 sky130_fd_sc_hd__nand3_1 _1621_ (.A(net241),
    .B(_0384_),
    .C(_0394_),
    .Y(_0398_));
 sky130_fd_sc_hd__xor2_1 _1622_ (.A(net242),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__a221oi_1 _1623_ (.A1(net207),
    .A2(_0372_),
    .B1(_0361_),
    .B2(net158),
    .C1(_0367_),
    .Y(_0400_));
 sky130_fd_sc_hd__a211oi_1 _1624_ (.A1(_0379_),
    .A2(_0399_),
    .B1(_0400_),
    .C1(_0383_),
    .Y(net446));
 sky130_fd_sc_hd__nand4_1 _1625_ (.A(net241),
    .B(net242),
    .C(_0376_),
    .D(_0394_),
    .Y(_0401_));
 sky130_fd_sc_hd__xor2_2 _1626_ (.A(net243),
    .B(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__a221oi_2 _1627_ (.A1(net208),
    .A2(_0372_),
    .B1(_0361_),
    .B2(_0646_),
    .C1(_0367_),
    .Y(_0403_));
 sky130_fd_sc_hd__a211oi_4 _1628_ (.A1(_0379_),
    .A2(_0402_),
    .B1(_0403_),
    .C1(_0383_),
    .Y(net447));
 sky130_fd_sc_hd__nand2_1 _1629_ (.A(_0384_),
    .B(_0394_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand3_1 _1630_ (.A(net241),
    .B(net242),
    .C(net243),
    .Y(_0405_));
 sky130_fd_sc_hd__nor2_1 _1631_ (.A(_0404_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__xnor2_1 _1632_ (.A(net244),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__buf_6 _1633_ (.A(_0315_),
    .X(_0408_));
 sky130_fd_sc_hd__a221oi_1 _1634_ (.A1(net209),
    .A2(_0372_),
    .B1(_0361_),
    .B2(net159),
    .C1(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__a211oi_1 _1635_ (.A1(_0379_),
    .A2(_0407_),
    .B1(_0409_),
    .C1(_0383_),
    .Y(net448));
 sky130_fd_sc_hd__nand4_1 _1636_ (.A(net241),
    .B(net242),
    .C(net243),
    .D(net244),
    .Y(_0410_));
 sky130_fd_sc_hd__nor2_1 _1637_ (.A(_0395_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__xnor2_1 _1638_ (.A(net245),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__buf_8 _1639_ (.A(_0307_),
    .X(_0413_));
 sky130_fd_sc_hd__a221oi_1 _1640_ (.A1(net210),
    .A2(_0413_),
    .B1(_0360_),
    .B2(net160),
    .C1(_0408_),
    .Y(_0414_));
 sky130_fd_sc_hd__a211oi_2 _1641_ (.A1(_0379_),
    .A2(_0412_),
    .B1(_0414_),
    .C1(_0383_),
    .Y(net449));
 sky130_fd_sc_hd__inv_1 _1642_ (.A(net245),
    .Y(_0415_));
 sky130_fd_sc_hd__nor3_1 _1643_ (.A(_0415_),
    .B(_0404_),
    .C(_0410_),
    .Y(_0416_));
 sky130_fd_sc_hd__xnor2_1 _1644_ (.A(net246),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__a221oi_2 _1645_ (.A1(net211),
    .A2(_0413_),
    .B1(_0360_),
    .B2(net161),
    .C1(_0408_),
    .Y(_0418_));
 sky130_fd_sc_hd__a211oi_4 _1646_ (.A1(_0379_),
    .A2(_0417_),
    .B1(_0418_),
    .C1(_0383_),
    .Y(net450));
 sky130_fd_sc_hd__clkbuf_16 _1647_ (.A(_0315_),
    .X(_0419_));
 sky130_fd_sc_hd__nor2_1 _1648_ (.A(_0415_),
    .B(_0410_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand4_1 _1649_ (.A(net246),
    .B(_0376_),
    .C(_0394_),
    .D(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__xor2_1 _1650_ (.A(net247),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__a221oi_4 _1651_ (.A1(net212),
    .A2(_0413_),
    .B1(_0360_),
    .B2(net162),
    .C1(_0408_),
    .Y(_0423_));
 sky130_fd_sc_hd__clkbuf_16 _1652_ (.A(_0303_),
    .X(_0424_));
 sky130_fd_sc_hd__a211oi_4 _1653_ (.A1(_0419_),
    .A2(_0422_),
    .B1(_0423_),
    .C1(_0424_),
    .Y(net451));
 sky130_fd_sc_hd__mux2i_2 _1654_ (.A0(net248),
    .A1(_0864_),
    .S(net112),
    .Y(_0425_));
 sky130_fd_sc_hd__mux2_1 _1655_ (.A0(_0625_),
    .A1(net135),
    .S(_0332_),
    .X(_0426_));
 sky130_fd_sc_hd__a221oi_2 _1656_ (.A1(net213),
    .A2(_0413_),
    .B1(_0426_),
    .B2(_0311_),
    .C1(_0408_),
    .Y(_0427_));
 sky130_fd_sc_hd__a211oi_4 _1657_ (.A1(_0419_),
    .A2(_0425_),
    .B1(_0427_),
    .C1(_0424_),
    .Y(net452));
 sky130_fd_sc_hd__nand3_1 _1658_ (.A(net246),
    .B(net247),
    .C(_0420_),
    .Y(_0428_));
 sky130_fd_sc_hd__nor2_1 _1659_ (.A(_0404_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__xnor2_1 _1660_ (.A(net249),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__a221oi_4 _1661_ (.A1(net214),
    .A2(_0413_),
    .B1(_0360_),
    .B2(_0645_),
    .C1(_0408_),
    .Y(_0431_));
 sky130_fd_sc_hd__a211oi_4 _1662_ (.A1(_0419_),
    .A2(_0430_),
    .B1(_0431_),
    .C1(_0424_),
    .Y(net453));
 sky130_fd_sc_hd__inv_1 _1663_ (.A(net249),
    .Y(_0432_));
 sky130_fd_sc_hd__nor3_1 _1664_ (.A(_0432_),
    .B(_0395_),
    .C(_0428_),
    .Y(_0433_));
 sky130_fd_sc_hd__xnor2_1 _1665_ (.A(net250),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__a221oi_2 _1666_ (.A1(net215),
    .A2(_0413_),
    .B1(_0360_),
    .B2(_0641_),
    .C1(_0408_),
    .Y(_0435_));
 sky130_fd_sc_hd__a211oi_4 _1667_ (.A1(_0419_),
    .A2(_0434_),
    .B1(_0435_),
    .C1(_0424_),
    .Y(net454));
 sky130_fd_sc_hd__nand2_1 _1668_ (.A(net112),
    .B(_0863_),
    .Y(_0436_));
 sky130_fd_sc_hd__xor2_2 _1669_ (.A(net251),
    .B(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__nand2_1 _1670_ (.A(_0223_),
    .B(net136),
    .Y(_0438_));
 sky130_fd_sc_hd__o21ai_2 _1671_ (.A1(_0654_),
    .A2(_0223_),
    .B1(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a221oi_4 _1672_ (.A1(net216),
    .A2(_0413_),
    .B1(_0439_),
    .B2(_0310_),
    .C1(_0408_),
    .Y(_0440_));
 sky130_fd_sc_hd__a211oi_4 _1673_ (.A1(_0419_),
    .A2(_0437_),
    .B1(_0440_),
    .C1(_0424_),
    .Y(net455));
 sky130_fd_sc_hd__xor2_1 _1674_ (.A(net252),
    .B(_0318_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(_0628_),
    .A1(net137),
    .S(_0332_),
    .X(_0442_));
 sky130_fd_sc_hd__a221oi_2 _1676_ (.A1(net217),
    .A2(_0413_),
    .B1(_0442_),
    .B2(_0310_),
    .C1(_0408_),
    .Y(_0443_));
 sky130_fd_sc_hd__a211oi_4 _1677_ (.A1(_0419_),
    .A2(_0441_),
    .B1(_0443_),
    .C1(_0424_),
    .Y(net456));
 sky130_fd_sc_hd__xor2_1 _1678_ (.A(net253),
    .B(_0326_),
    .X(_0444_));
 sky130_fd_sc_hd__clkinvlp_4 _1679_ (.A(_0636_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _1680_ (.A(_0223_),
    .B(net138),
    .Y(_0446_));
 sky130_fd_sc_hd__o21ai_0 _1681_ (.A1(_0445_),
    .A2(_0223_),
    .B1(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__a221oi_2 _1682_ (.A1(net218),
    .A2(_0413_),
    .B1(_0447_),
    .B2(_0310_),
    .C1(_0408_),
    .Y(_0448_));
 sky130_fd_sc_hd__a211oi_4 _1683_ (.A1(_0419_),
    .A2(_0444_),
    .B1(_0448_),
    .C1(_0424_),
    .Y(net457));
 sky130_fd_sc_hd__nor2_1 _1684_ (.A(_0318_),
    .B(_0319_),
    .Y(_0449_));
 sky130_fd_sc_hd__xnor2_1 _1685_ (.A(net254),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(_0635_),
    .A1(net139),
    .S(_0332_),
    .X(_0451_));
 sky130_fd_sc_hd__a221oi_2 _1687_ (.A1(net219),
    .A2(_0413_),
    .B1(_0451_),
    .B2(_0310_),
    .C1(_0315_),
    .Y(_0452_));
 sky130_fd_sc_hd__a211oi_4 _1688_ (.A1(_0419_),
    .A2(_0450_),
    .B1(_0452_),
    .C1(_0424_),
    .Y(net458));
 sky130_fd_sc_hd__xnor2_1 _1689_ (.A(net255),
    .B(_0328_),
    .Y(_0453_));
 sky130_fd_sc_hd__mux2_2 _1690_ (.A0(net168),
    .A1(net140),
    .S(_0332_),
    .X(_0454_));
 sky130_fd_sc_hd__a221oi_4 _1691_ (.A1(net220),
    .A2(_0307_),
    .B1(_0454_),
    .B2(_0310_),
    .C1(_0315_),
    .Y(_0455_));
 sky130_fd_sc_hd__a211oi_4 _1692_ (.A1(_0419_),
    .A2(_0453_),
    .B1(_0455_),
    .C1(_0424_),
    .Y(net459));
 sky130_fd_sc_hd__nand2_1 _1693_ (.A(net255),
    .B(_0320_),
    .Y(_0456_));
 sky130_fd_sc_hd__xor2_1 _1694_ (.A(net256),
    .B(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_2 _1695_ (.A0(net169),
    .A1(net141),
    .S(_0332_),
    .X(_0458_));
 sky130_fd_sc_hd__a221oi_4 _1696_ (.A1(net221),
    .A2(_0307_),
    .B1(_0458_),
    .B2(_0310_),
    .C1(_0315_),
    .Y(_0459_));
 sky130_fd_sc_hd__a211oi_4 _1697_ (.A1(_0419_),
    .A2(_0457_),
    .B1(_0459_),
    .C1(_0424_),
    .Y(net460));
 sky130_fd_sc_hd__nand3_1 _1698_ (.A(net255),
    .B(net256),
    .C(_0328_),
    .Y(_0460_));
 sky130_fd_sc_hd__xor2_1 _1699_ (.A(net257),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _1700_ (.A0(net170),
    .A1(net142),
    .S(net113),
    .X(_0462_));
 sky130_fd_sc_hd__a221oi_2 _1701_ (.A1(net222),
    .A2(_0307_),
    .B1(_0462_),
    .B2(_0310_),
    .C1(_0315_),
    .Y(_0463_));
 sky130_fd_sc_hd__a211oi_4 _1702_ (.A1(_0313_),
    .A2(_0461_),
    .B1(_0463_),
    .C1(_0303_),
    .Y(net461));
 sky130_fd_sc_hd__nand2_4 _1703_ (.A(_0743_),
    .B(_0762_),
    .Y(_0464_));
 sky130_fd_sc_hd__nor3_2 _1704_ (.A(_0631_),
    .B(_0779_),
    .C(_0464_),
    .Y(net462));
 sky130_fd_sc_hd__nor2_2 _1705_ (.A(_0844_),
    .B(_0836_),
    .Y(_0465_));
 sky130_fd_sc_hd__nand3_4 _1706_ (.A(_0703_),
    .B(_0723_),
    .C(_0730_),
    .Y(_0466_));
 sky130_fd_sc_hd__nor2_2 _1707_ (.A(\controller_i.ctrl_fsm_cs[0] ),
    .B(_0805_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand2_4 _1708_ (.A(_0848_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__o2111ai_4 _1709_ (.A1(_0465_),
    .A2(_0303_),
    .B1(_0466_),
    .C1(_0468_),
    .D1(_0790_),
    .Y(net467));
 sky130_fd_sc_hd__nand2_2 _1710_ (.A(_0466_),
    .B(_0468_),
    .Y(net469));
 sky130_fd_sc_hd__o21ai_4 _1711_ (.A1(net40),
    .A2(net358),
    .B1(_0467_),
    .Y(net471));
 sky130_fd_sc_hd__inv_1 _1712_ (.A(net358),
    .Y(_0469_));
 sky130_fd_sc_hd__a21oi_2 _1713_ (.A1(net40),
    .A2(_0469_),
    .B1(_0468_),
    .Y(net472));
 sky130_fd_sc_hd__and3_1 _1714_ (.A(net40),
    .B(_0469_),
    .C(_0467_),
    .X(net473));
 sky130_fd_sc_hd__nand2_4 _1715_ (.A(_0790_),
    .B(_0468_),
    .Y(net474));
 sky130_fd_sc_hd__nand2_2 _1716_ (.A(_0758_),
    .B(_0853_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor2_2 _1717_ (.A(_0622_),
    .B(_0470_),
    .Y(net476));
 sky130_fd_sc_hd__nor2_2 _1718_ (.A(_0760_),
    .B(_0779_),
    .Y(net478));
 sky130_fd_sc_hd__clkinv_2 _1719_ (.A(_0466_),
    .Y(net484));
 sky130_fd_sc_hd__or4_1 _1720_ (.A(net189),
    .B(net188),
    .C(net175),
    .D(net174),
    .X(_0471_));
 sky130_fd_sc_hd__nor3_1 _1721_ (.A(net177),
    .B(net176),
    .C(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__nor4_1 _1722_ (.A(net185),
    .B(net184),
    .C(net187),
    .D(net186),
    .Y(_0473_));
 sky130_fd_sc_hd__nor2_1 _1723_ (.A(net183),
    .B(net182),
    .Y(_0474_));
 sky130_fd_sc_hd__nor2_1 _1724_ (.A(net173),
    .B(net178),
    .Y(_0475_));
 sky130_fd_sc_hd__nand4_1 _1725_ (.A(_0472_),
    .B(_0473_),
    .C(_0474_),
    .D(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2b_1 _1726_ (.A_N(net671),
    .B(net171),
    .Y(_0477_));
 sky130_fd_sc_hd__o21ai_1 _1727_ (.A1(net181),
    .A2(_0476_),
    .B1(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_1 _1728_ (.A(net174),
    .Y(_0479_));
 sky130_fd_sc_hd__inv_1 _1729_ (.A(net186),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_1 _1730_ (.A(net182),
    .Y(_0481_));
 sky130_fd_sc_hd__a21oi_1 _1731_ (.A1(net181),
    .A2(_0481_),
    .B1(net183),
    .Y(_0482_));
 sky130_fd_sc_hd__o21bai_1 _1732_ (.A1(net184),
    .A2(_0482_),
    .B1_N(net185),
    .Y(_0483_));
 sky130_fd_sc_hd__a21oi_1 _1733_ (.A1(_0480_),
    .A2(_0483_),
    .B1(net187),
    .Y(_0484_));
 sky130_fd_sc_hd__o21bai_1 _1734_ (.A1(net188),
    .A2(_0484_),
    .B1_N(net189),
    .Y(_0485_));
 sky130_fd_sc_hd__a21oi_1 _1735_ (.A1(_0479_),
    .A2(_0485_),
    .B1(net175),
    .Y(_0486_));
 sky130_fd_sc_hd__o21bai_1 _1736_ (.A1(net176),
    .A2(_0486_),
    .B1_N(net177),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_1 _1737_ (.A(net178),
    .B(_0466_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _1738_ (.A(_0715_),
    .B(_0812_),
    .Y(_0489_));
 sky130_fd_sc_hd__and2_0 _1739_ (.A(_0693_),
    .B(_0699_),
    .X(_0490_));
 sky130_fd_sc_hd__nor4_1 _1740_ (.A(net155),
    .B(_0689_),
    .C(_0645_),
    .D(_0641_),
    .Y(_0491_));
 sky130_fd_sc_hd__nand4_4 _1741_ (.A(_0490_),
    .B(_0715_),
    .C(_0491_),
    .D(_0811_),
    .Y(_0492_));
 sky130_fd_sc_hd__nand2_1 _1742_ (.A(net258),
    .B(net259),
    .Y(_0493_));
 sky130_fd_sc_hd__o32ai_4 _1743_ (.A1(_0711_),
    .A2(_0787_),
    .A3(_0489_),
    .B1(_0492_),
    .B2(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__nor3_1 _1744_ (.A(_0315_),
    .B(_0307_),
    .C(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__nor2_1 _1745_ (.A(_0303_),
    .B(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__a221o_2 _1746_ (.A1(net484),
    .A2(_0478_),
    .B1(_0487_),
    .B2(_0488_),
    .C1(_0496_),
    .X(net479));
 sky130_fd_sc_hd__nand2_1 _1747_ (.A(_0720_),
    .B(_0715_),
    .Y(_0497_));
 sky130_fd_sc_hd__a211oi_2 _1748_ (.A1(\controller_i.store_err_q ),
    .A2(_0497_),
    .B1(_0494_),
    .C1(_0311_),
    .Y(_0498_));
 sky130_fd_sc_hd__nor3_1 _1749_ (.A(net185),
    .B(net184),
    .C(_0474_),
    .Y(_0499_));
 sky130_fd_sc_hd__nor3_1 _1750_ (.A(net187),
    .B(net186),
    .C(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__nor3_1 _1751_ (.A(net189),
    .B(net188),
    .C(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2_1 _1752_ (.A(net177),
    .B(net176),
    .Y(_0502_));
 sky130_fd_sc_hd__o31a_1 _1753_ (.A1(net175),
    .A2(net174),
    .A3(_0501_),
    .B1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__nor3_1 _1754_ (.A(net178),
    .B(_0478_),
    .C(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__o32ai_4 _1755_ (.A1(_0313_),
    .A2(_0303_),
    .A3(_0498_),
    .B1(_0504_),
    .B2(_0466_),
    .Y(net480));
 sky130_fd_sc_hd__nor2_1 _1756_ (.A(net181),
    .B(_0476_),
    .Y(_0505_));
 sky130_fd_sc_hd__nor2_1 _1757_ (.A(net180),
    .B(net179),
    .Y(_0506_));
 sky130_fd_sc_hd__nor2b_1 _1758_ (.A(net178),
    .B_N(_0477_),
    .Y(_0507_));
 sky130_fd_sc_hd__o211ai_1 _1759_ (.A1(_0471_),
    .A2(_0473_),
    .B1(_0507_),
    .C1(_0502_),
    .Y(_0508_));
 sky130_fd_sc_hd__a21oi_2 _1760_ (.A1(_0505_),
    .A2(_0506_),
    .B1(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nor2_2 _1761_ (.A(_0724_),
    .B(_0782_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand3_2 _1762_ (.A(_0304_),
    .B(_0510_),
    .C(_0308_),
    .Y(_0511_));
 sky130_fd_sc_hd__o21ai_4 _1763_ (.A1(_0466_),
    .A2(_0509_),
    .B1(_0511_),
    .Y(net481));
 sky130_fd_sc_hd__nand2_1 _1764_ (.A(net179),
    .B(_0505_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand3_1 _1765_ (.A(_0472_),
    .B(_0507_),
    .C(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _1766_ (.A(net484),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__o21ai_2 _1767_ (.A1(_0303_),
    .A2(_0492_),
    .B1(_0514_),
    .Y(net482));
 sky130_fd_sc_hd__a21oi_2 _1768_ (.A1(_0505_),
    .A2(_0477_),
    .B1(_0466_),
    .Y(net483));
 sky130_fd_sc_hd__a21boi_4 _1769_ (.A1(_0847_),
    .A2(_0510_),
    .B1_N(_0805_),
    .Y(net485));
 sky130_fd_sc_hd__o21ai_4 _1770_ (.A1(_0847_),
    .A2(_0303_),
    .B1(_0805_),
    .Y(net486));
 sky130_fd_sc_hd__o31a_2 _1771_ (.A1(_0624_),
    .A2(_0661_),
    .A3(_0700_),
    .B1(_0718_),
    .X(net560));
 sky130_fd_sc_hd__o21ai_1 _1772_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0788_),
    .Y(_0515_));
 sky130_fd_sc_hd__o21ai_4 _1773_ (.A1(_0704_),
    .A2(_0726_),
    .B1(_0515_),
    .Y(net561));
 sky130_fd_sc_hd__o21ai_1 _1774_ (.A1(_0703_),
    .A2(_0845_),
    .B1(\controller_i.ctrl_fsm_cs[2] ),
    .Y(_0516_));
 sky130_fd_sc_hd__a21oi_1 _1775_ (.A1(_0779_),
    .A2(_0849_),
    .B1(_0777_),
    .Y(_0517_));
 sky130_fd_sc_hd__a221o_4 _1776_ (.A1(_0792_),
    .A2(_0794_),
    .B1(_0516_),
    .B2(_0705_),
    .C1(_0517_),
    .X(net562));
 sky130_fd_sc_hd__nor3_4 _1777_ (.A(_0607_),
    .B(_0753_),
    .C(_0464_),
    .Y(net563));
 sky130_fd_sc_hd__nor3_2 _1778_ (.A(_0633_),
    .B(_0636_),
    .C(_0753_),
    .Y(net564));
 sky130_fd_sc_hd__nor2_1 _1779_ (.A(_0649_),
    .B(_0753_),
    .Y(net565));
 sky130_fd_sc_hd__nor3_2 _1780_ (.A(_0659_),
    .B(_0660_),
    .C(_0753_),
    .Y(net566));
 sky130_fd_sc_hd__nor2_8 _1781_ (.A(_0445_),
    .B(_0851_),
    .Y(net599));
 sky130_fd_sc_hd__nor2_2 _1782_ (.A(_0610_),
    .B(_0470_),
    .Y(net600));
 sky130_fd_sc_hd__nand2_1 _1783_ (.A(_0646_),
    .B(_0687_),
    .Y(_0518_));
 sky130_fd_sc_hd__or4_4 _1784_ (.A(_0683_),
    .B(_0648_),
    .C(_0642_),
    .D(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__a21oi_1 _1785_ (.A1(_0660_),
    .A2(_0644_),
    .B1(_0659_),
    .Y(_0520_));
 sky130_fd_sc_hd__nor2_2 _1786_ (.A(_0519_),
    .B(_0520_),
    .Y(net666));
 sky130_fd_sc_hd__nor2_2 _1787_ (.A(_0644_),
    .B(_0519_),
    .Y(net667));
 sky130_fd_sc_hd__o21ai_0 _1788_ (.A1(_0659_),
    .A2(_0633_),
    .B1(_0660_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _1789_ (.A(_0624_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nor2_2 _1790_ (.A(_0519_),
    .B(_0522_),
    .Y(net669));
 sky130_fd_sc_hd__mux2i_1 _1791_ (.A0(_0633_),
    .A1(_0634_),
    .S(_0660_),
    .Y(_0523_));
 sky130_fd_sc_hd__nor2_2 _1792_ (.A(_0519_),
    .B(_0523_),
    .Y(net670));
 sky130_fd_sc_hd__or2_1 _1793_ (.A(_0777_),
    .B(net466),
    .X(net672));
 sky130_fd_sc_hd__a21o_1 _1794_ (.A1(_0722_),
    .A2(_0808_),
    .B1(_0706_),
    .X(_0524_));
 sky130_fd_sc_hd__nand2_1 _1795_ (.A(_0805_),
    .B(_0524_),
    .Y(net673));
 sky130_fd_sc_hd__nor3_2 _1796_ (.A(_0697_),
    .B(_0737_),
    .C(_0783_),
    .Y(net674));
 sky130_fd_sc_hd__or2_1 _1797_ (.A(_0748_),
    .B(_0749_),
    .X(_0525_));
 sky130_fd_sc_hd__nand2_1 _1798_ (.A(_0722_),
    .B(_0704_),
    .Y(_0526_));
 sky130_fd_sc_hd__and3_2 _1799_ (.A(branch_set),
    .B(_0777_),
    .C(_0304_),
    .X(net682));
 sky130_fd_sc_hd__a211o_1 _1800_ (.A1(_0788_),
    .A2(_0526_),
    .B1(net682),
    .C1(net469),
    .X(_0527_));
 sky130_fd_sc_hd__a31oi_4 _1801_ (.A1(_0707_),
    .A2(_0829_),
    .A3(_0837_),
    .B1(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__o21ai_2 _1802_ (.A1(_0525_),
    .A2(_0302_),
    .B1(_0528_),
    .Y(net675));
 sky130_fd_sc_hd__nor2_4 _1803_ (.A(_0750_),
    .B(_0302_),
    .Y(net677));
 sky130_fd_sc_hd__a21oi_1 _1804_ (.A1(_0752_),
    .A2(_0753_),
    .B1(_0607_),
    .Y(_0529_));
 sky130_fd_sc_hd__a21o_2 _1805_ (.A1(net260),
    .A2(_0852_),
    .B1(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__nor3_4 _1806_ (.A(_0622_),
    .B(_0470_),
    .C(_0530_),
    .Y(net678));
 sky130_fd_sc_hd__nor3_4 _1807_ (.A(net224),
    .B(_0753_),
    .C(_0464_),
    .Y(net679));
 sky130_fd_sc_hd__nor2_4 _1808_ (.A(_0525_),
    .B(_0302_),
    .Y(net680));
 sky130_fd_sc_hd__nor3_4 _1809_ (.A(_0610_),
    .B(_0470_),
    .C(_0530_),
    .Y(net681));
 sky130_fd_sc_hd__or3_1 _1810_ (.A(_0633_),
    .B(_0445_),
    .C(_0677_),
    .X(_0531_));
 sky130_fd_sc_hd__a21oi_1 _1811_ (.A1(_0635_),
    .A2(_0531_),
    .B1(_0625_),
    .Y(_0532_));
 sky130_fd_sc_hd__a21oi_1 _1812_ (.A1(_0635_),
    .A2(_0671_),
    .B1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__nor3_4 _1813_ (.A(net165),
    .B(_0675_),
    .C(_0533_),
    .Y(net693));
 sky130_fd_sc_hd__a21oi_4 _1814_ (.A1(_0635_),
    .A2(_0628_),
    .B1(_0683_),
    .Y(net694));
 sky130_fd_sc_hd__clkbuf_4 _1815_ (.A(_0769_),
    .X(_0534_));
 sky130_fd_sc_hd__nand2_2 _1816_ (.A(net4),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__nand2_2 _1817_ (.A(net261),
    .B(_0632_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_8 _1818_ (.A(_0535_),
    .B(_0536_),
    .Y(net700));
 sky130_fd_sc_hd__nand2_1 _1819_ (.A(net5),
    .B(_0534_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_2 _1820_ (.A(net262),
    .B(_0632_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_8 _1821_ (.A(_0537_),
    .B(_0538_),
    .Y(net701));
 sky130_fd_sc_hd__nand2_1 _1822_ (.A(net6),
    .B(_0534_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _1823_ (.A(net263),
    .B(_0632_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_4 _1824_ (.A(_0539_),
    .B(_0540_),
    .Y(net702));
 sky130_fd_sc_hd__nand2_1 _1825_ (.A(net7),
    .B(_0534_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_2 _1826_ (.A(net264),
    .B(_0632_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_8 _1827_ (.A(_0541_),
    .B(_0542_),
    .Y(net703));
 sky130_fd_sc_hd__nand2_1 _1828_ (.A(net8),
    .B(_0534_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand2_1 _1829_ (.A(net265),
    .B(_0632_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_4 _1830_ (.A(_0543_),
    .B(_0544_),
    .Y(net704));
 sky130_fd_sc_hd__nand2_1 _1831_ (.A(net9),
    .B(_0534_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_2 _1832_ (.A(net266),
    .B(_0632_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_8 _1833_ (.A(_0545_),
    .B(_0546_),
    .Y(net705));
 sky130_fd_sc_hd__nand2_1 _1834_ (.A(net10),
    .B(_0534_),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _1835_ (.A(net267),
    .B(_0632_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_8 _1836_ (.A(_0547_),
    .B(_0548_),
    .Y(net706));
 sky130_fd_sc_hd__nand2_1 _1837_ (.A(net11),
    .B(_0534_),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_2 _1838_ (.A(net268),
    .B(_0632_),
    .Y(_0550_));
 sky130_fd_sc_hd__nand2_8 _1839_ (.A(_0549_),
    .B(_0550_),
    .Y(net707));
 sky130_fd_sc_hd__nand2_1 _1840_ (.A(net12),
    .B(_0534_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _1841_ (.A(net269),
    .B(_0632_),
    .Y(_0552_));
 sky130_fd_sc_hd__nand2_4 _1842_ (.A(_0551_),
    .B(_0552_),
    .Y(net708));
 sky130_fd_sc_hd__nand2_2 _1843_ (.A(net13),
    .B(_0534_),
    .Y(_0553_));
 sky130_fd_sc_hd__buf_4 _1844_ (.A(_0631_),
    .X(_0554_));
 sky130_fd_sc_hd__nand2_1 _1845_ (.A(net270),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand2_8 _1846_ (.A(_0553_),
    .B(_0555_),
    .Y(net709));
 sky130_fd_sc_hd__buf_4 _1847_ (.A(_0769_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_2 _1848_ (.A(net14),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__nand2_2 _1849_ (.A(net271),
    .B(_0554_),
    .Y(_0558_));
 sky130_fd_sc_hd__nand2_8 _1850_ (.A(_0557_),
    .B(_0558_),
    .Y(net710));
 sky130_fd_sc_hd__nand2_1 _1851_ (.A(net15),
    .B(_0556_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_2 _1852_ (.A(net272),
    .B(_0554_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_8 _1853_ (.A(_0559_),
    .B(_0560_),
    .Y(net711));
 sky130_fd_sc_hd__nand2_2 _1854_ (.A(net16),
    .B(_0556_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_2 _1855_ (.A(net273),
    .B(_0554_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_8 _1856_ (.A(_0561_),
    .B(_0562_),
    .Y(net712));
 sky130_fd_sc_hd__nand2_2 _1857_ (.A(net17),
    .B(_0556_),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2_2 _1858_ (.A(net274),
    .B(_0554_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_8 _1859_ (.A(_0563_),
    .B(_0564_),
    .Y(net713));
 sky130_fd_sc_hd__nand2_1 _1860_ (.A(net18),
    .B(_0556_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_2 _1861_ (.A(net275),
    .B(_0554_),
    .Y(_0566_));
 sky130_fd_sc_hd__nand2_8 _1862_ (.A(_0565_),
    .B(_0566_),
    .Y(net714));
 sky130_fd_sc_hd__nand2_1 _1863_ (.A(net19),
    .B(_0556_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_2 _1864_ (.A(net276),
    .B(_0554_),
    .Y(_0568_));
 sky130_fd_sc_hd__nand2_8 _1865_ (.A(_0567_),
    .B(_0568_),
    .Y(net715));
 sky130_fd_sc_hd__nand2_2 _1866_ (.A(net20),
    .B(_0556_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_2 _1867_ (.A(net277),
    .B(_0554_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_8 _1868_ (.A(_0569_),
    .B(_0570_),
    .Y(net716));
 sky130_fd_sc_hd__nand2_1 _1869_ (.A(net21),
    .B(_0556_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_2 _1870_ (.A(net278),
    .B(_0554_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2_8 _1871_ (.A(_0571_),
    .B(_0572_),
    .Y(net717));
 sky130_fd_sc_hd__nand2_1 _1872_ (.A(net22),
    .B(_0556_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_2 _1873_ (.A(net279),
    .B(_0554_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_8 _1874_ (.A(_0573_),
    .B(_0574_),
    .Y(net718));
 sky130_fd_sc_hd__nand2_2 _1875_ (.A(net23),
    .B(_0556_),
    .Y(_0575_));
 sky130_fd_sc_hd__buf_6 _1876_ (.A(_0631_),
    .X(_0576_));
 sky130_fd_sc_hd__nand2_2 _1877_ (.A(net280),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nand2_8 _1878_ (.A(_0575_),
    .B(_0577_),
    .Y(net719));
 sky130_fd_sc_hd__buf_4 _1879_ (.A(_0769_),
    .X(_0578_));
 sky130_fd_sc_hd__nand2_2 _1880_ (.A(net24),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_2 _1881_ (.A(net281),
    .B(_0576_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_8 _1882_ (.A(_0579_),
    .B(_0580_),
    .Y(net720));
 sky130_fd_sc_hd__nand2_2 _1883_ (.A(net25),
    .B(_0578_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_2 _1884_ (.A(net282),
    .B(_0576_),
    .Y(_0582_));
 sky130_fd_sc_hd__nand2_8 _1885_ (.A(_0581_),
    .B(_0582_),
    .Y(net721));
 sky130_fd_sc_hd__nand2_1 _1886_ (.A(net26),
    .B(_0578_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_2 _1887_ (.A(net283),
    .B(_0576_),
    .Y(_0584_));
 sky130_fd_sc_hd__nand2_8 _1888_ (.A(_0583_),
    .B(_0584_),
    .Y(net722));
 sky130_fd_sc_hd__nand2_1 _1889_ (.A(net27),
    .B(_0578_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_2 _1890_ (.A(net284),
    .B(_0576_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_8 _1891_ (.A(_0585_),
    .B(_0586_),
    .Y(net723));
 sky130_fd_sc_hd__nand2_1 _1892_ (.A(net28),
    .B(_0578_),
    .Y(_0587_));
 sky130_fd_sc_hd__nand2_2 _1893_ (.A(net285),
    .B(_0576_),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2_8 _1894_ (.A(_0587_),
    .B(_0588_),
    .Y(net724));
 sky130_fd_sc_hd__nand2_1 _1895_ (.A(net29),
    .B(_0578_),
    .Y(_0589_));
 sky130_fd_sc_hd__nand2_2 _1896_ (.A(net286),
    .B(_0576_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_8 _1897_ (.A(_0589_),
    .B(_0590_),
    .Y(net725));
 sky130_fd_sc_hd__nand2_2 _1898_ (.A(net30),
    .B(_0578_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_2 _1899_ (.A(net287),
    .B(_0576_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_8 _1900_ (.A(_0591_),
    .B(_0592_),
    .Y(net726));
 sky130_fd_sc_hd__nand2_1 _1901_ (.A(net31),
    .B(_0578_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(net288),
    .B(_0576_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_8 _1903_ (.A(_0593_),
    .B(_0594_),
    .Y(net727));
 sky130_fd_sc_hd__nand2_1 _1904_ (.A(net32),
    .B(_0578_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_2 _1905_ (.A(net289),
    .B(_0576_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_8 _1906_ (.A(_0595_),
    .B(_0596_),
    .Y(net728));
 sky130_fd_sc_hd__nand2_1 _1907_ (.A(net33),
    .B(_0578_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_2 _1908_ (.A(net290),
    .B(_0631_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2_8 _1909_ (.A(_0597_),
    .B(_0598_),
    .Y(net729));
 sky130_fd_sc_hd__nand2_1 _1910_ (.A(net34),
    .B(_0769_),
    .Y(_0599_));
 sky130_fd_sc_hd__nand2_2 _1911_ (.A(net291),
    .B(_0631_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_8 _1912_ (.A(_0599_),
    .B(_0600_),
    .Y(net730));
 sky130_fd_sc_hd__nand2_2 _1913_ (.A(net35),
    .B(_0769_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2_2 _1914_ (.A(net292),
    .B(_0631_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_8 _1915_ (.A(_0601_),
    .B(_0602_),
    .Y(net731));
 sky130_fd_sc_hd__o22ai_2 _1916_ (.A1(net165),
    .A2(_0648_),
    .B1(_0678_),
    .B2(net558),
    .Y(_0603_));
 sky130_fd_sc_hd__a31oi_2 _1917_ (.A1(net143),
    .A2(net153),
    .A3(_0603_),
    .B1(_0769_),
    .Y(_0604_));
 sky130_fd_sc_hd__o21ai_0 _1918_ (.A1(_0607_),
    .A2(_0753_),
    .B1(_0758_),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _1919_ (.A(net41),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor4_4 _1920_ (.A(net43),
    .B(_0464_),
    .C(_0604_),
    .D(_0606_),
    .Y(net732));
 sky130_fd_sc_hd__ha_1 _1921_ (.A(_0859_),
    .B(_0860_),
    .COUT(_0861_),
    .SUM(_0862_));
 sky130_fd_sc_hd__ha_1 _1922_ (.A(net237),
    .B(net248),
    .COUT(_0863_),
    .SUM(_0864_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__conb_1 _1992__802 (.HI(net802));
 sky130_fd_sc_hd__buf_4 _1925_ (.A(net733),
    .X(bt_a_operand_o[0]));
 sky130_fd_sc_hd__buf_4 _1926_ (.A(net734),
    .X(bt_a_operand_o[1]));
 sky130_fd_sc_hd__buf_4 _1927_ (.A(net735),
    .X(bt_a_operand_o[2]));
 sky130_fd_sc_hd__buf_4 _1928_ (.A(net736),
    .X(bt_a_operand_o[3]));
 sky130_fd_sc_hd__buf_4 _1929_ (.A(net737),
    .X(bt_a_operand_o[4]));
 sky130_fd_sc_hd__buf_4 _1930_ (.A(net738),
    .X(bt_a_operand_o[5]));
 sky130_fd_sc_hd__buf_4 _1931_ (.A(net739),
    .X(bt_a_operand_o[6]));
 sky130_fd_sc_hd__buf_4 _1932_ (.A(net740),
    .X(bt_a_operand_o[7]));
 sky130_fd_sc_hd__buf_4 _1933_ (.A(net741),
    .X(bt_a_operand_o[8]));
 sky130_fd_sc_hd__buf_4 _1934_ (.A(net742),
    .X(bt_a_operand_o[9]));
 sky130_fd_sc_hd__buf_4 _1935_ (.A(net743),
    .X(bt_a_operand_o[10]));
 sky130_fd_sc_hd__buf_4 _1936_ (.A(net744),
    .X(bt_a_operand_o[11]));
 sky130_fd_sc_hd__buf_4 _1937_ (.A(net745),
    .X(bt_a_operand_o[12]));
 sky130_fd_sc_hd__buf_4 _1938_ (.A(net746),
    .X(bt_a_operand_o[13]));
 sky130_fd_sc_hd__buf_4 _1939_ (.A(net747),
    .X(bt_a_operand_o[14]));
 sky130_fd_sc_hd__buf_4 _1940_ (.A(net748),
    .X(bt_a_operand_o[15]));
 sky130_fd_sc_hd__buf_4 _1941_ (.A(net749),
    .X(bt_a_operand_o[16]));
 sky130_fd_sc_hd__buf_4 _1942_ (.A(net750),
    .X(bt_a_operand_o[17]));
 sky130_fd_sc_hd__buf_4 _1943_ (.A(net751),
    .X(bt_a_operand_o[18]));
 sky130_fd_sc_hd__buf_4 _1944_ (.A(net752),
    .X(bt_a_operand_o[19]));
 sky130_fd_sc_hd__buf_4 _1945_ (.A(net753),
    .X(bt_a_operand_o[20]));
 sky130_fd_sc_hd__buf_4 _1946_ (.A(net754),
    .X(bt_a_operand_o[21]));
 sky130_fd_sc_hd__buf_4 _1947_ (.A(net755),
    .X(bt_a_operand_o[22]));
 sky130_fd_sc_hd__buf_4 _1948_ (.A(net756),
    .X(bt_a_operand_o[23]));
 sky130_fd_sc_hd__buf_4 _1949_ (.A(net757),
    .X(bt_a_operand_o[24]));
 sky130_fd_sc_hd__buf_4 _1950_ (.A(net758),
    .X(bt_a_operand_o[25]));
 sky130_fd_sc_hd__buf_4 _1951_ (.A(net759),
    .X(bt_a_operand_o[26]));
 sky130_fd_sc_hd__buf_4 _1952_ (.A(net760),
    .X(bt_a_operand_o[27]));
 sky130_fd_sc_hd__buf_4 _1953_ (.A(net761),
    .X(bt_a_operand_o[28]));
 sky130_fd_sc_hd__buf_4 _1954_ (.A(net762),
    .X(bt_a_operand_o[29]));
 sky130_fd_sc_hd__buf_4 _1955_ (.A(net763),
    .X(bt_a_operand_o[30]));
 sky130_fd_sc_hd__buf_4 _1956_ (.A(net764),
    .X(bt_a_operand_o[31]));
 sky130_fd_sc_hd__buf_4 _1957_ (.A(net765),
    .X(bt_b_operand_o[0]));
 sky130_fd_sc_hd__buf_4 _1958_ (.A(net766),
    .X(bt_b_operand_o[1]));
 sky130_fd_sc_hd__buf_4 _1959_ (.A(net767),
    .X(bt_b_operand_o[2]));
 sky130_fd_sc_hd__buf_4 _1960_ (.A(net768),
    .X(bt_b_operand_o[3]));
 sky130_fd_sc_hd__buf_4 _1961_ (.A(net769),
    .X(bt_b_operand_o[4]));
 sky130_fd_sc_hd__buf_4 _1962_ (.A(net770),
    .X(bt_b_operand_o[5]));
 sky130_fd_sc_hd__buf_4 _1963_ (.A(net771),
    .X(bt_b_operand_o[6]));
 sky130_fd_sc_hd__buf_4 _1964_ (.A(net772),
    .X(bt_b_operand_o[7]));
 sky130_fd_sc_hd__buf_4 _1965_ (.A(net773),
    .X(bt_b_operand_o[8]));
 sky130_fd_sc_hd__buf_4 _1966_ (.A(net774),
    .X(bt_b_operand_o[9]));
 sky130_fd_sc_hd__buf_4 _1967_ (.A(net775),
    .X(bt_b_operand_o[10]));
 sky130_fd_sc_hd__buf_4 _1968_ (.A(net776),
    .X(bt_b_operand_o[11]));
 sky130_fd_sc_hd__buf_4 _1969_ (.A(net777),
    .X(bt_b_operand_o[12]));
 sky130_fd_sc_hd__buf_4 _1970_ (.A(net778),
    .X(bt_b_operand_o[13]));
 sky130_fd_sc_hd__buf_4 _1971_ (.A(net779),
    .X(bt_b_operand_o[14]));
 sky130_fd_sc_hd__buf_4 _1972_ (.A(net780),
    .X(bt_b_operand_o[15]));
 sky130_fd_sc_hd__buf_4 _1973_ (.A(net781),
    .X(bt_b_operand_o[16]));
 sky130_fd_sc_hd__buf_4 _1974_ (.A(net782),
    .X(bt_b_operand_o[17]));
 sky130_fd_sc_hd__buf_4 _1975_ (.A(net783),
    .X(bt_b_operand_o[18]));
 sky130_fd_sc_hd__buf_4 _1976_ (.A(net784),
    .X(bt_b_operand_o[19]));
 sky130_fd_sc_hd__buf_4 _1977_ (.A(net785),
    .X(bt_b_operand_o[20]));
 sky130_fd_sc_hd__buf_4 _1978_ (.A(net786),
    .X(bt_b_operand_o[21]));
 sky130_fd_sc_hd__buf_4 _1979_ (.A(net787),
    .X(bt_b_operand_o[22]));
 sky130_fd_sc_hd__buf_4 _1980_ (.A(net788),
    .X(bt_b_operand_o[23]));
 sky130_fd_sc_hd__buf_4 _1981_ (.A(net789),
    .X(bt_b_operand_o[24]));
 sky130_fd_sc_hd__buf_4 _1982_ (.A(net790),
    .X(bt_b_operand_o[25]));
 sky130_fd_sc_hd__buf_4 _1983_ (.A(net791),
    .X(bt_b_operand_o[26]));
 sky130_fd_sc_hd__buf_4 _1984_ (.A(net792),
    .X(bt_b_operand_o[27]));
 sky130_fd_sc_hd__buf_4 _1985_ (.A(net793),
    .X(bt_b_operand_o[28]));
 sky130_fd_sc_hd__buf_4 _1986_ (.A(net794),
    .X(bt_b_operand_o[29]));
 sky130_fd_sc_hd__buf_4 _1987_ (.A(net795),
    .X(bt_b_operand_o[30]));
 sky130_fd_sc_hd__buf_4 _1988_ (.A(net796),
    .X(bt_b_operand_o[31]));
 sky130_fd_sc_hd__buf_4 _1989_ (.A(net797),
    .X(csr_save_wb_o));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1990_ (.A(net478),
    .X(net559));
 sky130_fd_sc_hd__buf_4 _1991_ (.A(net798),
    .X(instr_type_wb_o[0]));
 sky130_fd_sc_hd__buf_4 _1992_ (.A(net802),
    .X(instr_type_wb_o[1]));
 sky130_fd_sc_hd__buf_2 _1993_ (.A(net325),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 _1994_ (.A(net336),
    .X(net578));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1995_ (.A(net347),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_1 _1996_ (.A(net350),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_1 _1997_ (.A(net351),
    .X(net593));
 sky130_fd_sc_hd__buf_2 _1998_ (.A(net352),
    .X(net594));
 sky130_fd_sc_hd__buf_2 _1999_ (.A(net353),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_4 _2000_ (.A(net354),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_2 _2001_ (.A(net355),
    .X(net597));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2002_ (.A(net356),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_2 _2003_ (.A(net326),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_1 _2004_ (.A(net327),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_1 _2005_ (.A(net328),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_1 _2006_ (.A(net329),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 _2007_ (.A(net330),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_1 _2008_ (.A(net331),
    .X(net573));
 sky130_fd_sc_hd__buf_2 _2009_ (.A(net332),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 _2010_ (.A(net333),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_1 _2011_ (.A(net334),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_1 _2012_ (.A(net335),
    .X(net577));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2013_ (.A(net337),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_1 _2014_ (.A(net338),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 _2015_ (.A(net339),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 _2016_ (.A(net340),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 _2017_ (.A(net341),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_4 _2018_ (.A(net342),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_4 _2019_ (.A(net343),
    .X(net585));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2020_ (.A(net344),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_1 _2021_ (.A(net345),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 _2022_ (.A(net346),
    .X(net588));
 sky130_fd_sc_hd__buf_2 _2023_ (.A(net348),
    .X(net590));
 sky130_fd_sc_hd__buf_2 _2024_ (.A(net349),
    .X(net591));
 sky130_fd_sc_hd__buf_4 _2025_ (.A(net293),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_2 _2026_ (.A(net304),
    .X(net613));
 sky130_fd_sc_hd__buf_2 _2027_ (.A(net315),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_1 _2028_ (.A(net318),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_2 _2029_ (.A(net319),
    .X(net628));
 sky130_fd_sc_hd__buf_4 _2030_ (.A(net320),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 _2031_ (.A(net321),
    .X(net630));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2032_ (.A(net322),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_2 _2033_ (.A(net323),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_2 _2034_ (.A(net324),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_2 _2035_ (.A(net294),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_1 _2036_ (.A(net295),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_1 _2037_ (.A(net296),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_1 _2038_ (.A(net297),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_1 _2039_ (.A(net298),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_1 _2040_ (.A(net299),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 _2041_ (.A(net300),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 _2042_ (.A(net301),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_1 _2043_ (.A(net302),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_1 _2044_ (.A(net303),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_1 _2045_ (.A(net305),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_1 _2046_ (.A(net306),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_1 _2047_ (.A(net307),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 _2048_ (.A(net308),
    .X(net617));
 sky130_fd_sc_hd__buf_2 _2049_ (.A(net309),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_1 _2050_ (.A(net310),
    .X(net619));
 sky130_fd_sc_hd__buf_2 _2051_ (.A(net311),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_1 _2052_ (.A(net312),
    .X(net621));
 sky130_fd_sc_hd__buf_2 _2053_ (.A(net313),
    .X(net622));
 sky130_fd_sc_hd__buf_2 _2054_ (.A(net314),
    .X(net623));
 sky130_fd_sc_hd__buf_4 _2055_ (.A(net316),
    .X(net625));
 sky130_fd_sc_hd__buf_2 _2056_ (.A(net317),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_4 _2057_ (.A(net325),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_2 _2058_ (.A(net336),
    .X(net645));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2059_ (.A(net347),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_2 _2060_ (.A(net350),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_4 _2061_ (.A(net351),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_4 _2062_ (.A(net352),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_4 _2063_ (.A(net353),
    .X(net662));
 sky130_fd_sc_hd__buf_2 _2064_ (.A(net354),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_2 _2065_ (.A(net355),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_2 _2066_ (.A(net356),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_2 _2067_ (.A(net326),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_1 _2068_ (.A(net327),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 _2069_ (.A(net328),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_1 _2070_ (.A(net329),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_1 _2071_ (.A(net330),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_1 _2072_ (.A(net331),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_1 _2073_ (.A(net332),
    .X(net641));
 sky130_fd_sc_hd__buf_2 _2074_ (.A(net333),
    .X(net642));
 sky130_fd_sc_hd__buf_2 _2075_ (.A(net334),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_1 _2076_ (.A(net335),
    .X(net644));
 sky130_fd_sc_hd__buf_2 _2077_ (.A(net337),
    .X(net646));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2078_ (.A(net338),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_1 _2079_ (.A(net339),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_2 _2080_ (.A(net340),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_2 _2081_ (.A(net341),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 _2082_ (.A(net342),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_4 _2083_ (.A(net343),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_2 _2084_ (.A(net344),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_1 _2085_ (.A(net345),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_1 _2086_ (.A(net346),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_2 _2087_ (.A(net348),
    .X(net657));
 sky130_fd_sc_hd__buf_4 _2088_ (.A(net349),
    .X(net658));
 sky130_fd_sc_hd__buf_4 _2089_ (.A(net260),
    .X(net668));
 sky130_fd_sc_hd__buf_4 _2090_ (.A(net799),
    .X(nt_branch_mispredict_o));
 sky130_fd_sc_hd__clkbuf_1 _2091_ (.A(net675),
    .X(net676));
 sky130_fd_sc_hd__buf_4 _2092_ (.A(net148),
    .X(net683));
 sky130_fd_sc_hd__buf_6 _2093_ (.A(net149),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_8 _2094_ (.A(net150),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_8 _2095_ (.A(net151),
    .X(net686));
 sky130_fd_sc_hd__buf_6 _2096_ (.A(net152),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 _2097_ (.A(net154),
    .X(net688));
 sky130_fd_sc_hd__buf_4 _2098_ (.A(net155),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_4 _2099_ (.A(net156),
    .X(net690));
 sky130_fd_sc_hd__buf_6 _2100_ (.A(net157),
    .X(net691));
 sky130_fd_sc_hd__buf_6 _2101_ (.A(net158),
    .X(net692));
 sky130_fd_sc_hd__buf_4 _2102_ (.A(net800),
    .X(rf_rd_a_wb_match_o));
 sky130_fd_sc_hd__buf_4 _2103_ (.A(net801),
    .X(rf_rd_b_wb_match_o));
 sky130_fd_sc_hd__clkbuf_4 _2104_ (.A(net168),
    .X(net695));
 sky130_fd_sc_hd__buf_4 _2105_ (.A(net169),
    .X(net696));
 sky130_fd_sc_hd__buf_4 _2106_ (.A(net170),
    .X(net697));
 sky130_fd_sc_hd__buf_2 _2107_ (.A(net144),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_4 _2108_ (.A(net145),
    .X(net699));
 sky130_fd_sc_hd__dfrtp_4 \controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.D(_0000_),
    .Q(\controller_i.ctrl_fsm_cs[0] ),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.D(_0001_),
    .Q(\controller_i.ctrl_fsm_cs[1] ),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.D(_0002_),
    .Q(\controller_i.ctrl_fsm_cs[2] ),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.D(_0003_),
    .Q(\controller_i.ctrl_fsm_cs[3] ),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \controller_i.debug_mode_q$_DFFE_PN0P_  (.D(_0004_),
    .Q(net475),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \controller_i.exc_req_q$_DFF_PN0_  (.D(\controller_i.exc_req_d ),
    .Q(\controller_i.exc_req_q ),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \controller_i.illegal_insn_q$_DFF_PN0_  (.D(\controller_i.illegal_insn_d ),
    .Q(\controller_i.illegal_insn_q ),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \controller_i.load_err_q$_DFF_PN0_  (.D(net223),
    .Q(\controller_i.load_err_q ),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \controller_i.nmi_mode_q$_DFFE_PN0P_  (.D(_0005_),
    .Q(net671),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \controller_i.store_err_q$_DFF_PN0_  (.D(net225),
    .Q(\controller_i.store_err_q ),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \g_branch_set_flop.branch_set_q$_DFF_PN0_  (.D(branch_set_d),
    .Q(branch_set),
    .RESET_B(net357),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \id_fsm_q$_DFFE_PN0P_  (.D(_0006_),
    .Q(id_fsm_q),
    .RESET_B(net357),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[0]$_DFFE_PN0P_  (.D(_0007_),
    .Q(net490),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[10]$_DFFE_PN0P_  (.D(_0008_),
    .Q(net491),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[11]$_DFFE_PN0P_  (.D(_0009_),
    .Q(net492),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[12]$_DFFE_PN0P_  (.D(_0010_),
    .Q(net493),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[13]$_DFFE_PN0P_  (.D(_0011_),
    .Q(net494),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[14]$_DFFE_PN0P_  (.D(_0012_),
    .Q(net495),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[15]$_DFFE_PN0P_  (.D(_0013_),
    .Q(net496),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[16]$_DFFE_PN0P_  (.D(_0014_),
    .Q(net497),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[17]$_DFFE_PN0P_  (.D(_0015_),
    .Q(net498),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[18]$_DFFE_PN0P_  (.D(_0016_),
    .Q(net499),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[19]$_DFFE_PN0P_  (.D(_0017_),
    .Q(net500),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[1]$_DFFE_PN0P_  (.D(_0018_),
    .Q(net501),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[20]$_DFFE_PN0P_  (.D(_0019_),
    .Q(net502),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[21]$_DFFE_PN0P_  (.D(_0020_),
    .Q(net503),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[22]$_DFFE_PN0P_  (.D(_0021_),
    .Q(net504),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[23]$_DFFE_PN0P_  (.D(_0022_),
    .Q(net505),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[24]$_DFFE_PN0P_  (.D(_0023_),
    .Q(net506),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[25]$_DFFE_PN0P_  (.D(_0024_),
    .Q(net507),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[26]$_DFFE_PN0P_  (.D(_0025_),
    .Q(net508),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[27]$_DFFE_PN0P_  (.D(_0026_),
    .Q(net509),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[28]$_DFFE_PN0P_  (.D(_0027_),
    .Q(net510),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[29]$_DFFE_PN0P_  (.D(_0028_),
    .Q(net511),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[2]$_DFFE_PN0P_  (.D(_0029_),
    .Q(net512),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[30]$_DFFE_PN0P_  (.D(_0030_),
    .Q(net513),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[31]$_DFFE_PN0P_  (.D(_0031_),
    .Q(net514),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[32]$_DFFE_PN0P_  (.D(_0032_),
    .Q(net515),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[33]$_DFFE_PN0P_  (.D(_0033_),
    .Q(net516),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[34]$_DFFE_PN0P_  (.D(_0034_),
    .Q(net517),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[35]$_DFFE_PN0P_  (.D(_0035_),
    .Q(net518),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[36]$_DFFE_PN0P_  (.D(_0036_),
    .Q(net519),
    .RESET_B(net357),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[37]$_DFFE_PN0P_  (.D(_0037_),
    .Q(net520),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[38]$_DFFE_PN0P_  (.D(_0038_),
    .Q(net521),
    .RESET_B(net357),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[39]$_DFFE_PN0P_  (.D(_0039_),
    .Q(net522),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[3]$_DFFE_PN0P_  (.D(_0040_),
    .Q(net523),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[40]$_DFFE_PN0P_  (.D(_0041_),
    .Q(net524),
    .RESET_B(net357),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[41]$_DFFE_PN0P_  (.D(_0042_),
    .Q(net525),
    .RESET_B(net357),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[42]$_DFFE_PN0P_  (.D(_0043_),
    .Q(net526),
    .RESET_B(net357),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[43]$_DFFE_PN0P_  (.D(_0044_),
    .Q(net527),
    .RESET_B(net357),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[44]$_DFFE_PN0P_  (.D(_0045_),
    .Q(net528),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[45]$_DFFE_PN0P_  (.D(_0046_),
    .Q(net529),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[46]$_DFFE_PN0P_  (.D(_0047_),
    .Q(net530),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[47]$_DFFE_PN0P_  (.D(_0048_),
    .Q(net531),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[48]$_DFFE_PN0P_  (.D(_0049_),
    .Q(net532),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[49]$_DFFE_PN0P_  (.D(_0050_),
    .Q(net533),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[4]$_DFFE_PN0P_  (.D(_0051_),
    .Q(net534),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[50]$_DFFE_PN0P_  (.D(_0052_),
    .Q(net535),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[51]$_DFFE_PN0P_  (.D(_0053_),
    .Q(net536),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[52]$_DFFE_PN0P_  (.D(_0054_),
    .Q(net537),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[53]$_DFFE_PN0P_  (.D(_0055_),
    .Q(net538),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[54]$_DFFE_PN0P_  (.D(_0056_),
    .Q(net539),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[55]$_DFFE_PN0P_  (.D(_0057_),
    .Q(net540),
    .RESET_B(net357),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[56]$_DFFE_PN0P_  (.D(_0058_),
    .Q(net541),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[57]$_DFFE_PN0P_  (.D(_0059_),
    .Q(net542),
    .RESET_B(net357),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[58]$_DFFE_PN0P_  (.D(_0060_),
    .Q(net543),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \imd_val_q[59]$_DFFE_PN0P_  (.D(_0061_),
    .Q(net544),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[5]$_DFFE_PN0P_  (.D(_0062_),
    .Q(net545),
    .RESET_B(net357),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[60]$_DFFE_PN0P_  (.D(_0063_),
    .Q(net546),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[61]$_DFFE_PN0P_  (.D(_0064_),
    .Q(net547),
    .RESET_B(net357),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[62]$_DFFE_PN0P_  (.D(_0065_),
    .Q(net548),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[63]$_DFFE_PN0P_  (.D(_0066_),
    .Q(net549),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[64]$_DFFE_PN0P_  (.D(_0067_),
    .Q(net550),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[65]$_DFFE_PN0P_  (.D(_0068_),
    .Q(net551),
    .RESET_B(net357),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[66]$_DFFE_PN0P_  (.D(_0069_),
    .Q(net552),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[67]$_DFFE_PN0P_  (.D(_0070_),
    .Q(net553),
    .RESET_B(net357),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[6]$_DFFE_PN0P_  (.D(_0071_),
    .Q(net554),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[7]$_DFFE_PN0P_  (.D(_0072_),
    .Q(net555),
    .RESET_B(net357),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \imd_val_q[8]$_DFFE_PN0P_  (.D(_0073_),
    .Q(net556),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \imd_val_q[9]$_DFFE_PN0P_  (.D(_0074_),
    .Q(net557),
    .RESET_B(net357),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_1553 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(branch_decision_i),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(csr_mstatus_mie_i),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(csr_mstatus_tw_i),
    .X(net3));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input4 (.A(csr_rdata_i[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(csr_rdata_i[10]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(csr_rdata_i[11]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(csr_rdata_i[12]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(csr_rdata_i[13]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(csr_rdata_i[14]),
    .X(net9));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input10 (.A(csr_rdata_i[15]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(csr_rdata_i[16]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(csr_rdata_i[17]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(csr_rdata_i[18]),
    .X(net13));
 sky130_fd_sc_hd__buf_6 input14 (.A(csr_rdata_i[19]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(csr_rdata_i[1]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(csr_rdata_i[20]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(csr_rdata_i[21]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(csr_rdata_i[22]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(csr_rdata_i[23]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(csr_rdata_i[24]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(csr_rdata_i[25]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(csr_rdata_i[26]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(csr_rdata_i[27]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(csr_rdata_i[28]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(csr_rdata_i[29]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(csr_rdata_i[2]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(csr_rdata_i[30]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(csr_rdata_i[31]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(csr_rdata_i[3]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(csr_rdata_i[4]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(csr_rdata_i[5]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(csr_rdata_i[6]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(csr_rdata_i[7]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(csr_rdata_i[8]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(csr_rdata_i[9]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(data_ind_timing_i),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(debug_ebreakm_i),
    .X(net37));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input38 (.A(debug_ebreaku_i),
    .X(net38));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input39 (.A(debug_req_i),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input40 (.A(debug_single_step_i),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(ex_valid_i),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(illegal_c_insn_i),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(illegal_csr_insn_i),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(imd_val_d_ex_i[0]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(imd_val_d_ex_i[10]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(imd_val_d_ex_i[11]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(imd_val_d_ex_i[12]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(imd_val_d_ex_i[13]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(imd_val_d_ex_i[14]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(imd_val_d_ex_i[15]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(imd_val_d_ex_i[16]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(imd_val_d_ex_i[17]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(imd_val_d_ex_i[18]),
    .X(net53));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input54 (.A(imd_val_d_ex_i[19]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input55 (.A(imd_val_d_ex_i[1]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(imd_val_d_ex_i[20]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(imd_val_d_ex_i[21]),
    .X(net57));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input58 (.A(imd_val_d_ex_i[22]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(imd_val_d_ex_i[23]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(imd_val_d_ex_i[24]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(imd_val_d_ex_i[25]),
    .X(net61));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input62 (.A(imd_val_d_ex_i[26]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(imd_val_d_ex_i[27]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(imd_val_d_ex_i[28]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(imd_val_d_ex_i[29]),
    .X(net65));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input66 (.A(imd_val_d_ex_i[2]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(imd_val_d_ex_i[30]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(imd_val_d_ex_i[31]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(imd_val_d_ex_i[32]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(imd_val_d_ex_i[33]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(imd_val_d_ex_i[34]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(imd_val_d_ex_i[35]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(imd_val_d_ex_i[36]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(imd_val_d_ex_i[37]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(imd_val_d_ex_i[38]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(imd_val_d_ex_i[39]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(imd_val_d_ex_i[3]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(imd_val_d_ex_i[40]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(imd_val_d_ex_i[41]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(imd_val_d_ex_i[42]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(imd_val_d_ex_i[43]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(imd_val_d_ex_i[44]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(imd_val_d_ex_i[45]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(imd_val_d_ex_i[46]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(imd_val_d_ex_i[47]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(imd_val_d_ex_i[48]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(imd_val_d_ex_i[49]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(imd_val_d_ex_i[4]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(imd_val_d_ex_i[50]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(imd_val_d_ex_i[51]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(imd_val_d_ex_i[52]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(imd_val_d_ex_i[53]),
    .X(net92));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input93 (.A(imd_val_d_ex_i[54]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(imd_val_d_ex_i[55]),
    .X(net94));
 sky130_fd_sc_hd__buf_2 input95 (.A(imd_val_d_ex_i[56]),
    .X(net95));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input96 (.A(imd_val_d_ex_i[57]),
    .X(net96));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input97 (.A(imd_val_d_ex_i[58]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(imd_val_d_ex_i[59]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(imd_val_d_ex_i[5]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(imd_val_d_ex_i[60]),
    .X(net100));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input101 (.A(imd_val_d_ex_i[61]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(imd_val_d_ex_i[62]),
    .X(net102));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input103 (.A(imd_val_d_ex_i[63]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(imd_val_d_ex_i[64]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input105 (.A(imd_val_d_ex_i[65]),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input106 (.A(imd_val_d_ex_i[66]),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(imd_val_d_ex_i[67]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(imd_val_d_ex_i[6]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(imd_val_d_ex_i[7]),
    .X(net109));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input110 (.A(imd_val_d_ex_i[8]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input111 (.A(imd_val_d_ex_i[9]),
    .X(net111));
 sky130_fd_sc_hd__buf_6 input112 (.A(instr_fetch_err_plus2_i),
    .X(net112));
 sky130_fd_sc_hd__buf_6 input113 (.A(instr_is_compressed_i),
    .X(net113));
 sky130_fd_sc_hd__buf_2 input114 (.A(instr_rdata_alu_i[0]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(instr_rdata_alu_i[13]),
    .X(net115));
 sky130_fd_sc_hd__buf_4 input116 (.A(instr_rdata_alu_i[14]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(instr_rdata_alu_i[1]),
    .X(net117));
 sky130_fd_sc_hd__buf_4 input118 (.A(instr_rdata_alu_i[25]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(instr_rdata_alu_i[26]),
    .X(net119));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input120 (.A(instr_rdata_alu_i[27]),
    .X(net120));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input121 (.A(instr_rdata_alu_i[28]),
    .X(net121));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input122 (.A(instr_rdata_alu_i[29]),
    .X(net122));
 sky130_fd_sc_hd__buf_2 input123 (.A(instr_rdata_alu_i[30]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 input124 (.A(instr_rdata_alu_i[31]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(instr_rdata_alu_i[4]),
    .X(net125));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input126 (.A(instr_rdata_alu_i[6]),
    .X(net126));
 sky130_fd_sc_hd__buf_1 input127 (.A(instr_rdata_c_i[0]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(instr_rdata_c_i[10]),
    .X(net128));
 sky130_fd_sc_hd__buf_1 input129 (.A(instr_rdata_c_i[11]),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input130 (.A(instr_rdata_c_i[12]),
    .X(net130));
 sky130_fd_sc_hd__buf_2 input131 (.A(instr_rdata_c_i[13]),
    .X(net131));
 sky130_fd_sc_hd__buf_1 input132 (.A(instr_rdata_c_i[14]),
    .X(net132));
 sky130_fd_sc_hd__buf_1 input133 (.A(instr_rdata_c_i[15]),
    .X(net133));
 sky130_fd_sc_hd__buf_4 input134 (.A(instr_rdata_c_i[1]),
    .X(net134));
 sky130_fd_sc_hd__buf_4 input135 (.A(instr_rdata_c_i[2]),
    .X(net135));
 sky130_fd_sc_hd__buf_4 input136 (.A(instr_rdata_c_i[3]),
    .X(net136));
 sky130_fd_sc_hd__buf_4 input137 (.A(instr_rdata_c_i[4]),
    .X(net137));
 sky130_fd_sc_hd__buf_4 input138 (.A(instr_rdata_c_i[5]),
    .X(net138));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input139 (.A(instr_rdata_c_i[6]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input140 (.A(instr_rdata_c_i[7]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(instr_rdata_c_i[8]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(instr_rdata_c_i[9]),
    .X(net142));
 sky130_fd_sc_hd__buf_8 input143 (.A(instr_rdata_i[0]),
    .X(net143));
 sky130_fd_sc_hd__buf_4 input144 (.A(instr_rdata_i[10]),
    .X(net144));
 sky130_fd_sc_hd__buf_4 input145 (.A(instr_rdata_i[11]),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(instr_rdata_i[13]),
    .X(net146));
 sky130_fd_sc_hd__buf_4 input147 (.A(instr_rdata_i[14]),
    .X(net147));
 sky130_fd_sc_hd__buf_4 input148 (.A(instr_rdata_i[15]),
    .X(net148));
 sky130_fd_sc_hd__buf_4 input149 (.A(instr_rdata_i[16]),
    .X(net149));
 sky130_fd_sc_hd__buf_4 input150 (.A(instr_rdata_i[17]),
    .X(net150));
 sky130_fd_sc_hd__buf_4 input151 (.A(instr_rdata_i[18]),
    .X(net151));
 sky130_fd_sc_hd__buf_8 input152 (.A(instr_rdata_i[19]),
    .X(net152));
 sky130_fd_sc_hd__buf_6 input153 (.A(instr_rdata_i[1]),
    .X(net153));
 sky130_fd_sc_hd__buf_4 input154 (.A(instr_rdata_i[20]),
    .X(net154));
 sky130_fd_sc_hd__buf_8 input155 (.A(instr_rdata_i[21]),
    .X(net155));
 sky130_fd_sc_hd__buf_8 input156 (.A(instr_rdata_i[22]),
    .X(net156));
 sky130_fd_sc_hd__buf_8 input157 (.A(instr_rdata_i[23]),
    .X(net157));
 sky130_fd_sc_hd__buf_8 input158 (.A(instr_rdata_i[24]),
    .X(net158));
 sky130_fd_sc_hd__buf_8 input159 (.A(instr_rdata_i[26]),
    .X(net159));
 sky130_fd_sc_hd__buf_8 input160 (.A(instr_rdata_i[27]),
    .X(net160));
 sky130_fd_sc_hd__buf_8 input161 (.A(instr_rdata_i[28]),
    .X(net161));
 sky130_fd_sc_hd__buf_16 input162 (.A(instr_rdata_i[29]),
    .X(net162));
 sky130_fd_sc_hd__buf_2 input163 (.A(instr_rdata_i[30]),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(instr_rdata_i[31]),
    .X(net164));
 sky130_fd_sc_hd__buf_6 input165 (.A(instr_rdata_i[3]),
    .X(net165));
 sky130_fd_sc_hd__buf_4 input166 (.A(instr_rdata_i[4]),
    .X(net166));
 sky130_fd_sc_hd__buf_6 input167 (.A(instr_rdata_i[5]),
    .X(net167));
 sky130_fd_sc_hd__buf_4 input168 (.A(instr_rdata_i[7]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input169 (.A(instr_rdata_i[8]),
    .X(net169));
 sky130_fd_sc_hd__buf_4 input170 (.A(instr_rdata_i[9]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(irq_nm_i),
    .X(net171));
 sky130_fd_sc_hd__buf_2 input172 (.A(irq_pending_i),
    .X(net172));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input173 (.A(irqs_i[0]),
    .X(net173));
 sky130_fd_sc_hd__buf_2 input174 (.A(irqs_i[10]),
    .X(net174));
 sky130_fd_sc_hd__buf_2 input175 (.A(irqs_i[11]),
    .X(net175));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input176 (.A(irqs_i[12]),
    .X(net176));
 sky130_fd_sc_hd__buf_4 input177 (.A(irqs_i[13]),
    .X(net177));
 sky130_fd_sc_hd__buf_2 input178 (.A(irqs_i[14]),
    .X(net178));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input179 (.A(irqs_i[15]),
    .X(net179));
 sky130_fd_sc_hd__buf_1 input180 (.A(irqs_i[17]),
    .X(net180));
 sky130_fd_sc_hd__buf_2 input181 (.A(irqs_i[1]),
    .X(net181));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input182 (.A(irqs_i[2]),
    .X(net182));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input183 (.A(irqs_i[3]),
    .X(net183));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input184 (.A(irqs_i[4]),
    .X(net184));
 sky130_fd_sc_hd__buf_2 input185 (.A(irqs_i[5]),
    .X(net185));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input186 (.A(irqs_i[6]),
    .X(net186));
 sky130_fd_sc_hd__buf_2 input187 (.A(irqs_i[7]),
    .X(net187));
 sky130_fd_sc_hd__buf_2 input188 (.A(irqs_i[8]),
    .X(net188));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input189 (.A(irqs_i[9]),
    .X(net189));
 sky130_fd_sc_hd__buf_16 input190 (.A(lsu_addr_incr_req_i),
    .X(net190));
 sky130_fd_sc_hd__buf_1 input191 (.A(lsu_addr_last_i[0]),
    .X(net191));
 sky130_fd_sc_hd__buf_4 input192 (.A(lsu_addr_last_i[10]),
    .X(net192));
 sky130_fd_sc_hd__buf_1 input193 (.A(lsu_addr_last_i[11]),
    .X(net193));
 sky130_fd_sc_hd__buf_1 input194 (.A(lsu_addr_last_i[12]),
    .X(net194));
 sky130_fd_sc_hd__buf_1 input195 (.A(lsu_addr_last_i[13]),
    .X(net195));
 sky130_fd_sc_hd__buf_2 input196 (.A(lsu_addr_last_i[14]),
    .X(net196));
 sky130_fd_sc_hd__buf_1 input197 (.A(lsu_addr_last_i[15]),
    .X(net197));
 sky130_fd_sc_hd__buf_1 input198 (.A(lsu_addr_last_i[16]),
    .X(net198));
 sky130_fd_sc_hd__buf_1 input199 (.A(lsu_addr_last_i[17]),
    .X(net199));
 sky130_fd_sc_hd__buf_1 input200 (.A(lsu_addr_last_i[18]),
    .X(net200));
 sky130_fd_sc_hd__buf_1 input201 (.A(lsu_addr_last_i[19]),
    .X(net201));
 sky130_fd_sc_hd__buf_2 input202 (.A(lsu_addr_last_i[1]),
    .X(net202));
 sky130_fd_sc_hd__buf_1 input203 (.A(lsu_addr_last_i[20]),
    .X(net203));
 sky130_fd_sc_hd__buf_1 input204 (.A(lsu_addr_last_i[21]),
    .X(net204));
 sky130_fd_sc_hd__buf_1 input205 (.A(lsu_addr_last_i[22]),
    .X(net205));
 sky130_fd_sc_hd__buf_1 input206 (.A(lsu_addr_last_i[23]),
    .X(net206));
 sky130_fd_sc_hd__buf_1 input207 (.A(lsu_addr_last_i[24]),
    .X(net207));
 sky130_fd_sc_hd__buf_1 input208 (.A(lsu_addr_last_i[25]),
    .X(net208));
 sky130_fd_sc_hd__buf_1 input209 (.A(lsu_addr_last_i[26]),
    .X(net209));
 sky130_fd_sc_hd__buf_1 input210 (.A(lsu_addr_last_i[27]),
    .X(net210));
 sky130_fd_sc_hd__buf_1 input211 (.A(lsu_addr_last_i[28]),
    .X(net211));
 sky130_fd_sc_hd__buf_4 input212 (.A(lsu_addr_last_i[29]),
    .X(net212));
 sky130_fd_sc_hd__buf_4 input213 (.A(lsu_addr_last_i[2]),
    .X(net213));
 sky130_fd_sc_hd__buf_4 input214 (.A(lsu_addr_last_i[30]),
    .X(net214));
 sky130_fd_sc_hd__buf_6 input215 (.A(lsu_addr_last_i[31]),
    .X(net215));
 sky130_fd_sc_hd__buf_4 input216 (.A(lsu_addr_last_i[3]),
    .X(net216));
 sky130_fd_sc_hd__buf_2 input217 (.A(lsu_addr_last_i[4]),
    .X(net217));
 sky130_fd_sc_hd__buf_6 input218 (.A(lsu_addr_last_i[5]),
    .X(net218));
 sky130_fd_sc_hd__buf_2 input219 (.A(lsu_addr_last_i[6]),
    .X(net219));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input220 (.A(lsu_addr_last_i[7]),
    .X(net220));
 sky130_fd_sc_hd__buf_6 input221 (.A(lsu_addr_last_i[8]),
    .X(net221));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input222 (.A(lsu_addr_last_i[9]),
    .X(net222));
 sky130_fd_sc_hd__buf_4 input223 (.A(lsu_load_err_i),
    .X(net223));
 sky130_fd_sc_hd__buf_6 input224 (.A(lsu_resp_valid_i),
    .X(net224));
 sky130_fd_sc_hd__buf_2 input225 (.A(lsu_store_err_i),
    .X(net225));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input226 (.A(pc_id_i[0]),
    .X(net226));
 sky130_fd_sc_hd__buf_4 input227 (.A(pc_id_i[10]),
    .X(net227));
 sky130_fd_sc_hd__buf_4 input228 (.A(pc_id_i[11]),
    .X(net228));
 sky130_fd_sc_hd__buf_6 input229 (.A(pc_id_i[12]),
    .X(net229));
 sky130_fd_sc_hd__buf_2 input230 (.A(pc_id_i[13]),
    .X(net230));
 sky130_fd_sc_hd__buf_2 input231 (.A(pc_id_i[14]),
    .X(net231));
 sky130_fd_sc_hd__buf_2 input232 (.A(pc_id_i[15]),
    .X(net232));
 sky130_fd_sc_hd__buf_2 input233 (.A(pc_id_i[16]),
    .X(net233));
 sky130_fd_sc_hd__buf_2 input234 (.A(pc_id_i[17]),
    .X(net234));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input235 (.A(pc_id_i[18]),
    .X(net235));
 sky130_fd_sc_hd__buf_2 input236 (.A(pc_id_i[19]),
    .X(net236));
 sky130_fd_sc_hd__buf_4 input237 (.A(pc_id_i[1]),
    .X(net237));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input238 (.A(pc_id_i[20]),
    .X(net238));
 sky130_fd_sc_hd__buf_1 input239 (.A(pc_id_i[21]),
    .X(net239));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input240 (.A(pc_id_i[22]),
    .X(net240));
 sky130_fd_sc_hd__buf_4 input241 (.A(pc_id_i[23]),
    .X(net241));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input242 (.A(pc_id_i[24]),
    .X(net242));
 sky130_fd_sc_hd__buf_4 input243 (.A(pc_id_i[25]),
    .X(net243));
 sky130_fd_sc_hd__buf_4 input244 (.A(pc_id_i[26]),
    .X(net244));
 sky130_fd_sc_hd__buf_2 input245 (.A(pc_id_i[27]),
    .X(net245));
 sky130_fd_sc_hd__buf_4 input246 (.A(pc_id_i[28]),
    .X(net246));
 sky130_fd_sc_hd__buf_4 input247 (.A(pc_id_i[29]),
    .X(net247));
 sky130_fd_sc_hd__buf_4 input248 (.A(pc_id_i[2]),
    .X(net248));
 sky130_fd_sc_hd__buf_4 input249 (.A(pc_id_i[30]),
    .X(net249));
 sky130_fd_sc_hd__buf_4 input250 (.A(pc_id_i[31]),
    .X(net250));
 sky130_fd_sc_hd__buf_6 input251 (.A(pc_id_i[3]),
    .X(net251));
 sky130_fd_sc_hd__buf_6 input252 (.A(pc_id_i[4]),
    .X(net252));
 sky130_fd_sc_hd__buf_6 input253 (.A(pc_id_i[5]),
    .X(net253));
 sky130_fd_sc_hd__buf_4 input254 (.A(pc_id_i[6]),
    .X(net254));
 sky130_fd_sc_hd__buf_4 input255 (.A(pc_id_i[7]),
    .X(net255));
 sky130_fd_sc_hd__buf_4 input256 (.A(pc_id_i[8]),
    .X(net256));
 sky130_fd_sc_hd__buf_4 input257 (.A(pc_id_i[9]),
    .X(net257));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input258 (.A(priv_mode_i[0]),
    .X(net258));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input259 (.A(priv_mode_i[1]),
    .X(net259));
 sky130_fd_sc_hd__buf_8 input260 (.A(ready_wb_i),
    .X(net260));
 sky130_fd_sc_hd__buf_1 input261 (.A(result_ex_i[0]),
    .X(net261));
 sky130_fd_sc_hd__buf_1 input262 (.A(result_ex_i[10]),
    .X(net262));
 sky130_fd_sc_hd__buf_1 input263 (.A(result_ex_i[11]),
    .X(net263));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input264 (.A(result_ex_i[12]),
    .X(net264));
 sky130_fd_sc_hd__buf_1 input265 (.A(result_ex_i[13]),
    .X(net265));
 sky130_fd_sc_hd__buf_2 input266 (.A(result_ex_i[14]),
    .X(net266));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input267 (.A(result_ex_i[15]),
    .X(net267));
 sky130_fd_sc_hd__buf_4 input268 (.A(result_ex_i[16]),
    .X(net268));
 sky130_fd_sc_hd__buf_1 input269 (.A(result_ex_i[17]),
    .X(net269));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input270 (.A(result_ex_i[18]),
    .X(net270));
 sky130_fd_sc_hd__buf_2 input271 (.A(result_ex_i[19]),
    .X(net271));
 sky130_fd_sc_hd__buf_4 input272 (.A(result_ex_i[1]),
    .X(net272));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input273 (.A(result_ex_i[20]),
    .X(net273));
 sky130_fd_sc_hd__buf_1 input274 (.A(result_ex_i[21]),
    .X(net274));
 sky130_fd_sc_hd__buf_2 input275 (.A(result_ex_i[22]),
    .X(net275));
 sky130_fd_sc_hd__buf_1 input276 (.A(result_ex_i[23]),
    .X(net276));
 sky130_fd_sc_hd__buf_2 input277 (.A(result_ex_i[24]),
    .X(net277));
 sky130_fd_sc_hd__buf_4 input278 (.A(result_ex_i[25]),
    .X(net278));
 sky130_fd_sc_hd__buf_1 input279 (.A(result_ex_i[26]),
    .X(net279));
 sky130_fd_sc_hd__buf_4 input280 (.A(result_ex_i[27]),
    .X(net280));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input281 (.A(result_ex_i[28]),
    .X(net281));
 sky130_fd_sc_hd__buf_4 input282 (.A(result_ex_i[29]),
    .X(net282));
 sky130_fd_sc_hd__buf_4 input283 (.A(result_ex_i[2]),
    .X(net283));
 sky130_fd_sc_hd__buf_4 input284 (.A(result_ex_i[30]),
    .X(net284));
 sky130_fd_sc_hd__buf_4 input285 (.A(result_ex_i[31]),
    .X(net285));
 sky130_fd_sc_hd__buf_4 input286 (.A(result_ex_i[3]),
    .X(net286));
 sky130_fd_sc_hd__buf_4 input287 (.A(result_ex_i[4]),
    .X(net287));
 sky130_fd_sc_hd__buf_4 input288 (.A(result_ex_i[5]),
    .X(net288));
 sky130_fd_sc_hd__buf_4 input289 (.A(result_ex_i[6]),
    .X(net289));
 sky130_fd_sc_hd__buf_4 input290 (.A(result_ex_i[7]),
    .X(net290));
 sky130_fd_sc_hd__buf_4 input291 (.A(result_ex_i[8]),
    .X(net291));
 sky130_fd_sc_hd__buf_4 input292 (.A(result_ex_i[9]),
    .X(net292));
 sky130_fd_sc_hd__buf_4 input293 (.A(rf_rdata_a_i[0]),
    .X(net293));
 sky130_fd_sc_hd__buf_4 input294 (.A(rf_rdata_a_i[10]),
    .X(net294));
 sky130_fd_sc_hd__buf_4 input295 (.A(rf_rdata_a_i[11]),
    .X(net295));
 sky130_fd_sc_hd__buf_4 input296 (.A(rf_rdata_a_i[12]),
    .X(net296));
 sky130_fd_sc_hd__buf_4 input297 (.A(rf_rdata_a_i[13]),
    .X(net297));
 sky130_fd_sc_hd__buf_4 input298 (.A(rf_rdata_a_i[14]),
    .X(net298));
 sky130_fd_sc_hd__buf_4 input299 (.A(rf_rdata_a_i[15]),
    .X(net299));
 sky130_fd_sc_hd__buf_4 input300 (.A(rf_rdata_a_i[16]),
    .X(net300));
 sky130_fd_sc_hd__buf_4 input301 (.A(rf_rdata_a_i[17]),
    .X(net301));
 sky130_fd_sc_hd__buf_4 input302 (.A(rf_rdata_a_i[18]),
    .X(net302));
 sky130_fd_sc_hd__buf_4 input303 (.A(rf_rdata_a_i[19]),
    .X(net303));
 sky130_fd_sc_hd__buf_4 input304 (.A(rf_rdata_a_i[1]),
    .X(net304));
 sky130_fd_sc_hd__buf_4 input305 (.A(rf_rdata_a_i[20]),
    .X(net305));
 sky130_fd_sc_hd__buf_4 input306 (.A(rf_rdata_a_i[21]),
    .X(net306));
 sky130_fd_sc_hd__buf_4 input307 (.A(rf_rdata_a_i[22]),
    .X(net307));
 sky130_fd_sc_hd__buf_4 input308 (.A(rf_rdata_a_i[23]),
    .X(net308));
 sky130_fd_sc_hd__buf_2 input309 (.A(rf_rdata_a_i[24]),
    .X(net309));
 sky130_fd_sc_hd__buf_4 input310 (.A(rf_rdata_a_i[25]),
    .X(net310));
 sky130_fd_sc_hd__buf_4 input311 (.A(rf_rdata_a_i[26]),
    .X(net311));
 sky130_fd_sc_hd__buf_2 input312 (.A(rf_rdata_a_i[27]),
    .X(net312));
 sky130_fd_sc_hd__buf_2 input313 (.A(rf_rdata_a_i[28]),
    .X(net313));
 sky130_fd_sc_hd__buf_2 input314 (.A(rf_rdata_a_i[29]),
    .X(net314));
 sky130_fd_sc_hd__buf_4 input315 (.A(rf_rdata_a_i[2]),
    .X(net315));
 sky130_fd_sc_hd__buf_4 input316 (.A(rf_rdata_a_i[30]),
    .X(net316));
 sky130_fd_sc_hd__buf_4 input317 (.A(rf_rdata_a_i[31]),
    .X(net317));
 sky130_fd_sc_hd__buf_2 input318 (.A(rf_rdata_a_i[3]),
    .X(net318));
 sky130_fd_sc_hd__buf_2 input319 (.A(rf_rdata_a_i[4]),
    .X(net319));
 sky130_fd_sc_hd__buf_4 input320 (.A(rf_rdata_a_i[5]),
    .X(net320));
 sky130_fd_sc_hd__buf_4 input321 (.A(rf_rdata_a_i[6]),
    .X(net321));
 sky130_fd_sc_hd__buf_4 input322 (.A(rf_rdata_a_i[7]),
    .X(net322));
 sky130_fd_sc_hd__buf_4 input323 (.A(rf_rdata_a_i[8]),
    .X(net323));
 sky130_fd_sc_hd__buf_6 input324 (.A(rf_rdata_a_i[9]),
    .X(net324));
 sky130_fd_sc_hd__buf_4 input325 (.A(rf_rdata_b_i[0]),
    .X(net325));
 sky130_fd_sc_hd__buf_2 input326 (.A(rf_rdata_b_i[10]),
    .X(net326));
 sky130_fd_sc_hd__buf_4 input327 (.A(rf_rdata_b_i[11]),
    .X(net327));
 sky130_fd_sc_hd__buf_4 input328 (.A(rf_rdata_b_i[12]),
    .X(net328));
 sky130_fd_sc_hd__buf_4 input329 (.A(rf_rdata_b_i[13]),
    .X(net329));
 sky130_fd_sc_hd__buf_4 input330 (.A(rf_rdata_b_i[14]),
    .X(net330));
 sky130_fd_sc_hd__buf_4 input331 (.A(rf_rdata_b_i[15]),
    .X(net331));
 sky130_fd_sc_hd__buf_4 input332 (.A(rf_rdata_b_i[16]),
    .X(net332));
 sky130_fd_sc_hd__buf_4 input333 (.A(rf_rdata_b_i[17]),
    .X(net333));
 sky130_fd_sc_hd__buf_4 input334 (.A(rf_rdata_b_i[18]),
    .X(net334));
 sky130_fd_sc_hd__buf_2 input335 (.A(rf_rdata_b_i[19]),
    .X(net335));
 sky130_fd_sc_hd__buf_2 input336 (.A(rf_rdata_b_i[1]),
    .X(net336));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input337 (.A(rf_rdata_b_i[20]),
    .X(net337));
 sky130_fd_sc_hd__buf_2 input338 (.A(rf_rdata_b_i[21]),
    .X(net338));
 sky130_fd_sc_hd__buf_2 input339 (.A(rf_rdata_b_i[22]),
    .X(net339));
 sky130_fd_sc_hd__buf_2 input340 (.A(rf_rdata_b_i[23]),
    .X(net340));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input341 (.A(rf_rdata_b_i[24]),
    .X(net341));
 sky130_fd_sc_hd__buf_2 input342 (.A(rf_rdata_b_i[25]),
    .X(net342));
 sky130_fd_sc_hd__buf_4 input343 (.A(rf_rdata_b_i[26]),
    .X(net343));
 sky130_fd_sc_hd__buf_2 input344 (.A(rf_rdata_b_i[27]),
    .X(net344));
 sky130_fd_sc_hd__buf_2 input345 (.A(rf_rdata_b_i[28]),
    .X(net345));
 sky130_fd_sc_hd__buf_4 input346 (.A(rf_rdata_b_i[29]),
    .X(net346));
 sky130_fd_sc_hd__buf_4 input347 (.A(rf_rdata_b_i[2]),
    .X(net347));
 sky130_fd_sc_hd__buf_2 input348 (.A(rf_rdata_b_i[30]),
    .X(net348));
 sky130_fd_sc_hd__buf_2 input349 (.A(rf_rdata_b_i[31]),
    .X(net349));
 sky130_fd_sc_hd__buf_2 input350 (.A(rf_rdata_b_i[3]),
    .X(net350));
 sky130_fd_sc_hd__buf_2 input351 (.A(rf_rdata_b_i[4]),
    .X(net351));
 sky130_fd_sc_hd__buf_2 input352 (.A(rf_rdata_b_i[5]),
    .X(net352));
 sky130_fd_sc_hd__buf_4 input353 (.A(rf_rdata_b_i[6]),
    .X(net353));
 sky130_fd_sc_hd__buf_2 input354 (.A(rf_rdata_b_i[7]),
    .X(net354));
 sky130_fd_sc_hd__buf_2 input355 (.A(rf_rdata_b_i[8]),
    .X(net355));
 sky130_fd_sc_hd__buf_4 input356 (.A(rf_rdata_b_i[9]),
    .X(net356));
 sky130_fd_sc_hd__buf_16 input357 (.A(rst_ni),
    .X(net357));
 sky130_fd_sc_hd__buf_4 input358 (.A(trigger_match_i),
    .X(net358));
 sky130_fd_sc_hd__buf_1 output359 (.A(net359),
    .X(alu_operand_a_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output360 (.A(net360),
    .X(alu_operand_a_ex_o[10]));
 sky130_fd_sc_hd__buf_1 output361 (.A(net361),
    .X(alu_operand_a_ex_o[11]));
 sky130_fd_sc_hd__buf_1 output362 (.A(net362),
    .X(alu_operand_a_ex_o[12]));
 sky130_fd_sc_hd__buf_1 output363 (.A(net363),
    .X(alu_operand_a_ex_o[13]));
 sky130_fd_sc_hd__buf_1 output364 (.A(net364),
    .X(alu_operand_a_ex_o[14]));
 sky130_fd_sc_hd__buf_1 output365 (.A(net365),
    .X(alu_operand_a_ex_o[15]));
 sky130_fd_sc_hd__buf_1 output366 (.A(net366),
    .X(alu_operand_a_ex_o[16]));
 sky130_fd_sc_hd__buf_1 output367 (.A(net367),
    .X(alu_operand_a_ex_o[17]));
 sky130_fd_sc_hd__buf_1 output368 (.A(net368),
    .X(alu_operand_a_ex_o[18]));
 sky130_fd_sc_hd__buf_1 output369 (.A(net369),
    .X(alu_operand_a_ex_o[19]));
 sky130_fd_sc_hd__buf_1 output370 (.A(net370),
    .X(alu_operand_a_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output371 (.A(net371),
    .X(alu_operand_a_ex_o[20]));
 sky130_fd_sc_hd__buf_1 output372 (.A(net372),
    .X(alu_operand_a_ex_o[21]));
 sky130_fd_sc_hd__buf_1 output373 (.A(net373),
    .X(alu_operand_a_ex_o[22]));
 sky130_fd_sc_hd__buf_1 output374 (.A(net374),
    .X(alu_operand_a_ex_o[23]));
 sky130_fd_sc_hd__buf_1 output375 (.A(net375),
    .X(alu_operand_a_ex_o[24]));
 sky130_fd_sc_hd__buf_1 output376 (.A(net376),
    .X(alu_operand_a_ex_o[25]));
 sky130_fd_sc_hd__buf_1 output377 (.A(net377),
    .X(alu_operand_a_ex_o[26]));
 sky130_fd_sc_hd__buf_1 output378 (.A(net378),
    .X(alu_operand_a_ex_o[27]));
 sky130_fd_sc_hd__buf_1 output379 (.A(net379),
    .X(alu_operand_a_ex_o[28]));
 sky130_fd_sc_hd__buf_1 output380 (.A(net380),
    .X(alu_operand_a_ex_o[29]));
 sky130_fd_sc_hd__buf_1 output381 (.A(net381),
    .X(alu_operand_a_ex_o[2]));
 sky130_fd_sc_hd__buf_1 output382 (.A(net382),
    .X(alu_operand_a_ex_o[30]));
 sky130_fd_sc_hd__buf_1 output383 (.A(net383),
    .X(alu_operand_a_ex_o[31]));
 sky130_fd_sc_hd__buf_1 output384 (.A(net384),
    .X(alu_operand_a_ex_o[3]));
 sky130_fd_sc_hd__buf_1 output385 (.A(net385),
    .X(alu_operand_a_ex_o[4]));
 sky130_fd_sc_hd__buf_1 output386 (.A(net386),
    .X(alu_operand_a_ex_o[5]));
 sky130_fd_sc_hd__buf_1 output387 (.A(net387),
    .X(alu_operand_a_ex_o[6]));
 sky130_fd_sc_hd__buf_1 output388 (.A(net388),
    .X(alu_operand_a_ex_o[7]));
 sky130_fd_sc_hd__buf_1 output389 (.A(net389),
    .X(alu_operand_a_ex_o[8]));
 sky130_fd_sc_hd__buf_1 output390 (.A(net390),
    .X(alu_operand_a_ex_o[9]));
 sky130_fd_sc_hd__buf_1 output391 (.A(net391),
    .X(alu_operand_b_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output392 (.A(net392),
    .X(alu_operand_b_ex_o[10]));
 sky130_fd_sc_hd__buf_1 output393 (.A(net393),
    .X(alu_operand_b_ex_o[11]));
 sky130_fd_sc_hd__buf_1 output394 (.A(net394),
    .X(alu_operand_b_ex_o[12]));
 sky130_fd_sc_hd__buf_1 output395 (.A(net395),
    .X(alu_operand_b_ex_o[13]));
 sky130_fd_sc_hd__buf_1 output396 (.A(net396),
    .X(alu_operand_b_ex_o[14]));
 sky130_fd_sc_hd__buf_1 output397 (.A(net397),
    .X(alu_operand_b_ex_o[15]));
 sky130_fd_sc_hd__buf_1 output398 (.A(net398),
    .X(alu_operand_b_ex_o[16]));
 sky130_fd_sc_hd__buf_1 output399 (.A(net399),
    .X(alu_operand_b_ex_o[17]));
 sky130_fd_sc_hd__buf_1 output400 (.A(net400),
    .X(alu_operand_b_ex_o[18]));
 sky130_fd_sc_hd__buf_1 output401 (.A(net401),
    .X(alu_operand_b_ex_o[19]));
 sky130_fd_sc_hd__buf_1 output402 (.A(net402),
    .X(alu_operand_b_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output403 (.A(net403),
    .X(alu_operand_b_ex_o[20]));
 sky130_fd_sc_hd__buf_1 output404 (.A(net404),
    .X(alu_operand_b_ex_o[21]));
 sky130_fd_sc_hd__buf_1 output405 (.A(net405),
    .X(alu_operand_b_ex_o[22]));
 sky130_fd_sc_hd__buf_1 output406 (.A(net406),
    .X(alu_operand_b_ex_o[23]));
 sky130_fd_sc_hd__buf_1 output407 (.A(net407),
    .X(alu_operand_b_ex_o[24]));
 sky130_fd_sc_hd__buf_1 output408 (.A(net408),
    .X(alu_operand_b_ex_o[25]));
 sky130_fd_sc_hd__buf_1 output409 (.A(net409),
    .X(alu_operand_b_ex_o[26]));
 sky130_fd_sc_hd__buf_1 output410 (.A(net410),
    .X(alu_operand_b_ex_o[27]));
 sky130_fd_sc_hd__buf_1 output411 (.A(net411),
    .X(alu_operand_b_ex_o[28]));
 sky130_fd_sc_hd__buf_1 output412 (.A(net412),
    .X(alu_operand_b_ex_o[29]));
 sky130_fd_sc_hd__buf_1 output413 (.A(net413),
    .X(alu_operand_b_ex_o[2]));
 sky130_fd_sc_hd__buf_1 output414 (.A(net414),
    .X(alu_operand_b_ex_o[30]));
 sky130_fd_sc_hd__buf_1 output415 (.A(net415),
    .X(alu_operand_b_ex_o[31]));
 sky130_fd_sc_hd__buf_1 output416 (.A(net416),
    .X(alu_operand_b_ex_o[3]));
 sky130_fd_sc_hd__buf_1 output417 (.A(net417),
    .X(alu_operand_b_ex_o[4]));
 sky130_fd_sc_hd__buf_1 output418 (.A(net418),
    .X(alu_operand_b_ex_o[5]));
 sky130_fd_sc_hd__buf_1 output419 (.A(net419),
    .X(alu_operand_b_ex_o[6]));
 sky130_fd_sc_hd__buf_1 output420 (.A(net420),
    .X(alu_operand_b_ex_o[7]));
 sky130_fd_sc_hd__buf_1 output421 (.A(net421),
    .X(alu_operand_b_ex_o[8]));
 sky130_fd_sc_hd__buf_1 output422 (.A(net422),
    .X(alu_operand_b_ex_o[9]));
 sky130_fd_sc_hd__buf_1 output423 (.A(net423),
    .X(alu_operator_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output424 (.A(net424),
    .X(alu_operator_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output425 (.A(net425),
    .X(alu_operator_ex_o[2]));
 sky130_fd_sc_hd__buf_1 output426 (.A(net426),
    .X(alu_operator_ex_o[3]));
 sky130_fd_sc_hd__buf_1 output427 (.A(net427),
    .X(alu_operator_ex_o[4]));
 sky130_fd_sc_hd__buf_1 output428 (.A(net428),
    .X(alu_operator_ex_o[5]));
 sky130_fd_sc_hd__buf_1 output429 (.A(net429),
    .X(csr_access_o));
 sky130_fd_sc_hd__buf_1 output430 (.A(net430),
    .X(csr_mtval_o[0]));
 sky130_fd_sc_hd__buf_1 output431 (.A(net431),
    .X(csr_mtval_o[10]));
 sky130_fd_sc_hd__buf_1 output432 (.A(net432),
    .X(csr_mtval_o[11]));
 sky130_fd_sc_hd__buf_1 output433 (.A(net433),
    .X(csr_mtval_o[12]));
 sky130_fd_sc_hd__buf_1 output434 (.A(net434),
    .X(csr_mtval_o[13]));
 sky130_fd_sc_hd__buf_1 output435 (.A(net435),
    .X(csr_mtval_o[14]));
 sky130_fd_sc_hd__buf_1 output436 (.A(net436),
    .X(csr_mtval_o[15]));
 sky130_fd_sc_hd__buf_1 output437 (.A(net437),
    .X(csr_mtval_o[16]));
 sky130_fd_sc_hd__buf_1 output438 (.A(net438),
    .X(csr_mtval_o[17]));
 sky130_fd_sc_hd__buf_1 output439 (.A(net439),
    .X(csr_mtval_o[18]));
 sky130_fd_sc_hd__buf_1 output440 (.A(net440),
    .X(csr_mtval_o[19]));
 sky130_fd_sc_hd__buf_1 output441 (.A(net441),
    .X(csr_mtval_o[1]));
 sky130_fd_sc_hd__buf_1 output442 (.A(net442),
    .X(csr_mtval_o[20]));
 sky130_fd_sc_hd__buf_1 output443 (.A(net443),
    .X(csr_mtval_o[21]));
 sky130_fd_sc_hd__buf_1 output444 (.A(net444),
    .X(csr_mtval_o[22]));
 sky130_fd_sc_hd__buf_1 output445 (.A(net445),
    .X(csr_mtval_o[23]));
 sky130_fd_sc_hd__buf_1 output446 (.A(net446),
    .X(csr_mtval_o[24]));
 sky130_fd_sc_hd__buf_1 output447 (.A(net447),
    .X(csr_mtval_o[25]));
 sky130_fd_sc_hd__buf_1 output448 (.A(net448),
    .X(csr_mtval_o[26]));
 sky130_fd_sc_hd__buf_1 output449 (.A(net449),
    .X(csr_mtval_o[27]));
 sky130_fd_sc_hd__buf_1 output450 (.A(net450),
    .X(csr_mtval_o[28]));
 sky130_fd_sc_hd__buf_1 output451 (.A(net451),
    .X(csr_mtval_o[29]));
 sky130_fd_sc_hd__buf_1 output452 (.A(net452),
    .X(csr_mtval_o[2]));
 sky130_fd_sc_hd__buf_1 output453 (.A(net453),
    .X(csr_mtval_o[30]));
 sky130_fd_sc_hd__buf_1 output454 (.A(net454),
    .X(csr_mtval_o[31]));
 sky130_fd_sc_hd__buf_1 output455 (.A(net455),
    .X(csr_mtval_o[3]));
 sky130_fd_sc_hd__buf_1 output456 (.A(net456),
    .X(csr_mtval_o[4]));
 sky130_fd_sc_hd__buf_1 output457 (.A(net457),
    .X(csr_mtval_o[5]));
 sky130_fd_sc_hd__buf_1 output458 (.A(net458),
    .X(csr_mtval_o[6]));
 sky130_fd_sc_hd__buf_1 output459 (.A(net459),
    .X(csr_mtval_o[7]));
 sky130_fd_sc_hd__buf_1 output460 (.A(net460),
    .X(csr_mtval_o[8]));
 sky130_fd_sc_hd__buf_1 output461 (.A(net461),
    .X(csr_mtval_o[9]));
 sky130_fd_sc_hd__buf_1 output462 (.A(net462),
    .X(csr_op_en_o));
 sky130_fd_sc_hd__buf_1 output463 (.A(net463),
    .X(csr_op_o[0]));
 sky130_fd_sc_hd__buf_1 output464 (.A(net464),
    .X(csr_op_o[1]));
 sky130_fd_sc_hd__buf_1 output465 (.A(net465),
    .X(csr_restore_dret_id_o));
 sky130_fd_sc_hd__buf_1 output466 (.A(net466),
    .X(csr_restore_mret_id_o));
 sky130_fd_sc_hd__buf_1 output467 (.A(net467),
    .X(csr_save_cause_o));
 sky130_fd_sc_hd__buf_1 output468 (.A(net468),
    .X(csr_save_id_o));
 sky130_fd_sc_hd__buf_1 output469 (.A(net469),
    .X(csr_save_if_o));
 sky130_fd_sc_hd__buf_1 output470 (.A(net470),
    .X(ctrl_busy_o));
 sky130_fd_sc_hd__buf_1 output471 (.A(net471),
    .X(debug_cause_o[0]));
 sky130_fd_sc_hd__buf_1 output472 (.A(net472),
    .X(debug_cause_o[1]));
 sky130_fd_sc_hd__buf_1 output473 (.A(net473),
    .X(debug_cause_o[2]));
 sky130_fd_sc_hd__buf_1 output474 (.A(net474),
    .X(debug_csr_save_o));
 sky130_fd_sc_hd__buf_1 output475 (.A(net475),
    .X(debug_mode_o));
 sky130_fd_sc_hd__buf_1 output476 (.A(net476),
    .X(div_en_ex_o));
 sky130_fd_sc_hd__buf_1 output477 (.A(net477),
    .X(div_sel_ex_o));
 sky130_fd_sc_hd__buf_1 output478 (.A(net478),
    .X(en_wb_o));
 sky130_fd_sc_hd__buf_1 output479 (.A(net479),
    .X(exc_cause_o[0]));
 sky130_fd_sc_hd__buf_1 output480 (.A(net480),
    .X(exc_cause_o[1]));
 sky130_fd_sc_hd__buf_1 output481 (.A(net481),
    .X(exc_cause_o[2]));
 sky130_fd_sc_hd__buf_1 output482 (.A(net482),
    .X(exc_cause_o[3]));
 sky130_fd_sc_hd__buf_1 output483 (.A(net483),
    .X(exc_cause_o[4]));
 sky130_fd_sc_hd__buf_1 output484 (.A(net484),
    .X(exc_cause_o[5]));
 sky130_fd_sc_hd__buf_1 output485 (.A(net485),
    .X(exc_pc_mux_o[0]));
 sky130_fd_sc_hd__buf_1 output486 (.A(net486),
    .X(exc_pc_mux_o[1]));
 sky130_fd_sc_hd__buf_1 output487 (.A(net487),
    .X(icache_inval_o));
 sky130_fd_sc_hd__buf_1 output488 (.A(net488),
    .X(id_in_ready_o));
 sky130_fd_sc_hd__buf_1 output489 (.A(net489),
    .X(illegal_insn_o));
 sky130_fd_sc_hd__buf_1 output490 (.A(net490),
    .X(imd_val_q_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output491 (.A(net491),
    .X(imd_val_q_ex_o[10]));
 sky130_fd_sc_hd__buf_1 output492 (.A(net492),
    .X(imd_val_q_ex_o[11]));
 sky130_fd_sc_hd__buf_1 output493 (.A(net493),
    .X(imd_val_q_ex_o[12]));
 sky130_fd_sc_hd__buf_1 output494 (.A(net494),
    .X(imd_val_q_ex_o[13]));
 sky130_fd_sc_hd__buf_1 output495 (.A(net495),
    .X(imd_val_q_ex_o[14]));
 sky130_fd_sc_hd__buf_1 output496 (.A(net496),
    .X(imd_val_q_ex_o[15]));
 sky130_fd_sc_hd__buf_1 output497 (.A(net497),
    .X(imd_val_q_ex_o[16]));
 sky130_fd_sc_hd__buf_1 output498 (.A(net498),
    .X(imd_val_q_ex_o[17]));
 sky130_fd_sc_hd__buf_1 output499 (.A(net499),
    .X(imd_val_q_ex_o[18]));
 sky130_fd_sc_hd__buf_1 output500 (.A(net500),
    .X(imd_val_q_ex_o[19]));
 sky130_fd_sc_hd__buf_1 output501 (.A(net501),
    .X(imd_val_q_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output502 (.A(net502),
    .X(imd_val_q_ex_o[20]));
 sky130_fd_sc_hd__buf_1 output503 (.A(net503),
    .X(imd_val_q_ex_o[21]));
 sky130_fd_sc_hd__buf_1 output504 (.A(net504),
    .X(imd_val_q_ex_o[22]));
 sky130_fd_sc_hd__buf_1 output505 (.A(net505),
    .X(imd_val_q_ex_o[23]));
 sky130_fd_sc_hd__buf_1 output506 (.A(net506),
    .X(imd_val_q_ex_o[24]));
 sky130_fd_sc_hd__buf_1 output507 (.A(net507),
    .X(imd_val_q_ex_o[25]));
 sky130_fd_sc_hd__buf_1 output508 (.A(net508),
    .X(imd_val_q_ex_o[26]));
 sky130_fd_sc_hd__buf_1 output509 (.A(net509),
    .X(imd_val_q_ex_o[27]));
 sky130_fd_sc_hd__buf_1 output510 (.A(net510),
    .X(imd_val_q_ex_o[28]));
 sky130_fd_sc_hd__buf_1 output511 (.A(net511),
    .X(imd_val_q_ex_o[29]));
 sky130_fd_sc_hd__buf_1 output512 (.A(net512),
    .X(imd_val_q_ex_o[2]));
 sky130_fd_sc_hd__buf_1 output513 (.A(net513),
    .X(imd_val_q_ex_o[30]));
 sky130_fd_sc_hd__buf_1 output514 (.A(net514),
    .X(imd_val_q_ex_o[31]));
 sky130_fd_sc_hd__buf_1 output515 (.A(net515),
    .X(imd_val_q_ex_o[32]));
 sky130_fd_sc_hd__buf_1 output516 (.A(net516),
    .X(imd_val_q_ex_o[33]));
 sky130_fd_sc_hd__buf_1 output517 (.A(net517),
    .X(imd_val_q_ex_o[34]));
 sky130_fd_sc_hd__buf_1 output518 (.A(net518),
    .X(imd_val_q_ex_o[35]));
 sky130_fd_sc_hd__buf_1 output519 (.A(net519),
    .X(imd_val_q_ex_o[36]));
 sky130_fd_sc_hd__buf_1 output520 (.A(net520),
    .X(imd_val_q_ex_o[37]));
 sky130_fd_sc_hd__buf_1 output521 (.A(net521),
    .X(imd_val_q_ex_o[38]));
 sky130_fd_sc_hd__buf_1 output522 (.A(net522),
    .X(imd_val_q_ex_o[39]));
 sky130_fd_sc_hd__buf_1 output523 (.A(net523),
    .X(imd_val_q_ex_o[3]));
 sky130_fd_sc_hd__buf_1 output524 (.A(net524),
    .X(imd_val_q_ex_o[40]));
 sky130_fd_sc_hd__buf_1 output525 (.A(net525),
    .X(imd_val_q_ex_o[41]));
 sky130_fd_sc_hd__buf_1 output526 (.A(net526),
    .X(imd_val_q_ex_o[42]));
 sky130_fd_sc_hd__buf_1 output527 (.A(net527),
    .X(imd_val_q_ex_o[43]));
 sky130_fd_sc_hd__buf_1 output528 (.A(net528),
    .X(imd_val_q_ex_o[44]));
 sky130_fd_sc_hd__buf_1 output529 (.A(net529),
    .X(imd_val_q_ex_o[45]));
 sky130_fd_sc_hd__buf_1 output530 (.A(net530),
    .X(imd_val_q_ex_o[46]));
 sky130_fd_sc_hd__buf_1 output531 (.A(net531),
    .X(imd_val_q_ex_o[47]));
 sky130_fd_sc_hd__buf_1 output532 (.A(net532),
    .X(imd_val_q_ex_o[48]));
 sky130_fd_sc_hd__buf_1 output533 (.A(net533),
    .X(imd_val_q_ex_o[49]));
 sky130_fd_sc_hd__buf_1 output534 (.A(net534),
    .X(imd_val_q_ex_o[4]));
 sky130_fd_sc_hd__buf_1 output535 (.A(net535),
    .X(imd_val_q_ex_o[50]));
 sky130_fd_sc_hd__buf_1 output536 (.A(net536),
    .X(imd_val_q_ex_o[51]));
 sky130_fd_sc_hd__buf_1 output537 (.A(net537),
    .X(imd_val_q_ex_o[52]));
 sky130_fd_sc_hd__buf_1 output538 (.A(net538),
    .X(imd_val_q_ex_o[53]));
 sky130_fd_sc_hd__buf_1 output539 (.A(net539),
    .X(imd_val_q_ex_o[54]));
 sky130_fd_sc_hd__buf_1 output540 (.A(net540),
    .X(imd_val_q_ex_o[55]));
 sky130_fd_sc_hd__buf_1 output541 (.A(net541),
    .X(imd_val_q_ex_o[56]));
 sky130_fd_sc_hd__buf_1 output542 (.A(net542),
    .X(imd_val_q_ex_o[57]));
 sky130_fd_sc_hd__buf_1 output543 (.A(net543),
    .X(imd_val_q_ex_o[58]));
 sky130_fd_sc_hd__buf_1 output544 (.A(net544),
    .X(imd_val_q_ex_o[59]));
 sky130_fd_sc_hd__buf_1 output545 (.A(net545),
    .X(imd_val_q_ex_o[5]));
 sky130_fd_sc_hd__buf_1 output546 (.A(net546),
    .X(imd_val_q_ex_o[60]));
 sky130_fd_sc_hd__buf_1 output547 (.A(net547),
    .X(imd_val_q_ex_o[61]));
 sky130_fd_sc_hd__buf_1 output548 (.A(net548),
    .X(imd_val_q_ex_o[62]));
 sky130_fd_sc_hd__buf_1 output549 (.A(net549),
    .X(imd_val_q_ex_o[63]));
 sky130_fd_sc_hd__buf_1 output550 (.A(net550),
    .X(imd_val_q_ex_o[64]));
 sky130_fd_sc_hd__buf_1 output551 (.A(net551),
    .X(imd_val_q_ex_o[65]));
 sky130_fd_sc_hd__buf_1 output552 (.A(net552),
    .X(imd_val_q_ex_o[66]));
 sky130_fd_sc_hd__buf_1 output553 (.A(net553),
    .X(imd_val_q_ex_o[67]));
 sky130_fd_sc_hd__buf_1 output554 (.A(net554),
    .X(imd_val_q_ex_o[6]));
 sky130_fd_sc_hd__buf_1 output555 (.A(net555),
    .X(imd_val_q_ex_o[7]));
 sky130_fd_sc_hd__buf_1 output556 (.A(net556),
    .X(imd_val_q_ex_o[8]));
 sky130_fd_sc_hd__buf_1 output557 (.A(net557),
    .X(imd_val_q_ex_o[9]));
 sky130_fd_sc_hd__buf_1 output558 (.A(net558),
    .X(instr_first_cycle_id_o));
 sky130_fd_sc_hd__buf_1 output559 (.A(net559),
    .X(instr_id_done_o));
 sky130_fd_sc_hd__buf_1 output560 (.A(net560),
    .X(instr_perf_count_id_o));
 sky130_fd_sc_hd__buf_1 output561 (.A(net561),
    .X(instr_req_o));
 sky130_fd_sc_hd__buf_1 output562 (.A(net562),
    .X(instr_valid_clear_o));
 sky130_fd_sc_hd__buf_1 output563 (.A(net563),
    .X(lsu_req_o));
 sky130_fd_sc_hd__buf_1 output564 (.A(net564),
    .X(lsu_sign_ext_o));
 sky130_fd_sc_hd__buf_1 output565 (.A(net565),
    .X(lsu_type_o[0]));
 sky130_fd_sc_hd__buf_1 output566 (.A(net566),
    .X(lsu_type_o[1]));
 sky130_fd_sc_hd__buf_1 output567 (.A(net567),
    .X(lsu_wdata_o[0]));
 sky130_fd_sc_hd__buf_1 output568 (.A(net568),
    .X(lsu_wdata_o[10]));
 sky130_fd_sc_hd__buf_1 output569 (.A(net569),
    .X(lsu_wdata_o[11]));
 sky130_fd_sc_hd__buf_1 output570 (.A(net570),
    .X(lsu_wdata_o[12]));
 sky130_fd_sc_hd__buf_1 output571 (.A(net571),
    .X(lsu_wdata_o[13]));
 sky130_fd_sc_hd__buf_1 output572 (.A(net572),
    .X(lsu_wdata_o[14]));
 sky130_fd_sc_hd__buf_1 output573 (.A(net573),
    .X(lsu_wdata_o[15]));
 sky130_fd_sc_hd__buf_1 output574 (.A(net574),
    .X(lsu_wdata_o[16]));
 sky130_fd_sc_hd__buf_1 output575 (.A(net575),
    .X(lsu_wdata_o[17]));
 sky130_fd_sc_hd__buf_1 output576 (.A(net576),
    .X(lsu_wdata_o[18]));
 sky130_fd_sc_hd__buf_1 output577 (.A(net577),
    .X(lsu_wdata_o[19]));
 sky130_fd_sc_hd__buf_1 output578 (.A(net578),
    .X(lsu_wdata_o[1]));
 sky130_fd_sc_hd__buf_1 output579 (.A(net579),
    .X(lsu_wdata_o[20]));
 sky130_fd_sc_hd__buf_1 output580 (.A(net580),
    .X(lsu_wdata_o[21]));
 sky130_fd_sc_hd__buf_1 output581 (.A(net581),
    .X(lsu_wdata_o[22]));
 sky130_fd_sc_hd__buf_1 output582 (.A(net582),
    .X(lsu_wdata_o[23]));
 sky130_fd_sc_hd__buf_1 output583 (.A(net583),
    .X(lsu_wdata_o[24]));
 sky130_fd_sc_hd__buf_1 output584 (.A(net584),
    .X(lsu_wdata_o[25]));
 sky130_fd_sc_hd__buf_1 output585 (.A(net585),
    .X(lsu_wdata_o[26]));
 sky130_fd_sc_hd__buf_1 output586 (.A(net586),
    .X(lsu_wdata_o[27]));
 sky130_fd_sc_hd__buf_1 output587 (.A(net587),
    .X(lsu_wdata_o[28]));
 sky130_fd_sc_hd__buf_1 output588 (.A(net588),
    .X(lsu_wdata_o[29]));
 sky130_fd_sc_hd__buf_1 output589 (.A(net589),
    .X(lsu_wdata_o[2]));
 sky130_fd_sc_hd__buf_1 output590 (.A(net590),
    .X(lsu_wdata_o[30]));
 sky130_fd_sc_hd__buf_1 output591 (.A(net591),
    .X(lsu_wdata_o[31]));
 sky130_fd_sc_hd__buf_1 output592 (.A(net592),
    .X(lsu_wdata_o[3]));
 sky130_fd_sc_hd__buf_1 output593 (.A(net593),
    .X(lsu_wdata_o[4]));
 sky130_fd_sc_hd__buf_1 output594 (.A(net594),
    .X(lsu_wdata_o[5]));
 sky130_fd_sc_hd__buf_1 output595 (.A(net595),
    .X(lsu_wdata_o[6]));
 sky130_fd_sc_hd__buf_1 output596 (.A(net596),
    .X(lsu_wdata_o[7]));
 sky130_fd_sc_hd__buf_1 output597 (.A(net597),
    .X(lsu_wdata_o[8]));
 sky130_fd_sc_hd__buf_1 output598 (.A(net598),
    .X(lsu_wdata_o[9]));
 sky130_fd_sc_hd__buf_1 output599 (.A(net599),
    .X(lsu_we_o));
 sky130_fd_sc_hd__buf_1 output600 (.A(net600),
    .X(mult_en_ex_o));
 sky130_fd_sc_hd__buf_1 output601 (.A(net601),
    .X(mult_sel_ex_o));
 sky130_fd_sc_hd__buf_1 output602 (.A(net602),
    .X(multdiv_operand_a_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output603 (.A(net603),
    .X(multdiv_operand_a_ex_o[10]));
 sky130_fd_sc_hd__buf_1 output604 (.A(net604),
    .X(multdiv_operand_a_ex_o[11]));
 sky130_fd_sc_hd__buf_1 output605 (.A(net605),
    .X(multdiv_operand_a_ex_o[12]));
 sky130_fd_sc_hd__buf_1 output606 (.A(net606),
    .X(multdiv_operand_a_ex_o[13]));
 sky130_fd_sc_hd__buf_1 output607 (.A(net607),
    .X(multdiv_operand_a_ex_o[14]));
 sky130_fd_sc_hd__buf_1 output608 (.A(net608),
    .X(multdiv_operand_a_ex_o[15]));
 sky130_fd_sc_hd__buf_1 output609 (.A(net609),
    .X(multdiv_operand_a_ex_o[16]));
 sky130_fd_sc_hd__buf_1 output610 (.A(net610),
    .X(multdiv_operand_a_ex_o[17]));
 sky130_fd_sc_hd__buf_1 output611 (.A(net611),
    .X(multdiv_operand_a_ex_o[18]));
 sky130_fd_sc_hd__buf_1 output612 (.A(net612),
    .X(multdiv_operand_a_ex_o[19]));
 sky130_fd_sc_hd__buf_1 output613 (.A(net613),
    .X(multdiv_operand_a_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output614 (.A(net614),
    .X(multdiv_operand_a_ex_o[20]));
 sky130_fd_sc_hd__buf_1 output615 (.A(net615),
    .X(multdiv_operand_a_ex_o[21]));
 sky130_fd_sc_hd__buf_1 output616 (.A(net616),
    .X(multdiv_operand_a_ex_o[22]));
 sky130_fd_sc_hd__buf_1 output617 (.A(net617),
    .X(multdiv_operand_a_ex_o[23]));
 sky130_fd_sc_hd__buf_1 output618 (.A(net618),
    .X(multdiv_operand_a_ex_o[24]));
 sky130_fd_sc_hd__buf_1 output619 (.A(net619),
    .X(multdiv_operand_a_ex_o[25]));
 sky130_fd_sc_hd__buf_1 output620 (.A(net620),
    .X(multdiv_operand_a_ex_o[26]));
 sky130_fd_sc_hd__buf_1 output621 (.A(net621),
    .X(multdiv_operand_a_ex_o[27]));
 sky130_fd_sc_hd__buf_1 output622 (.A(net622),
    .X(multdiv_operand_a_ex_o[28]));
 sky130_fd_sc_hd__buf_1 output623 (.A(net623),
    .X(multdiv_operand_a_ex_o[29]));
 sky130_fd_sc_hd__buf_1 output624 (.A(net624),
    .X(multdiv_operand_a_ex_o[2]));
 sky130_fd_sc_hd__buf_1 output625 (.A(net625),
    .X(multdiv_operand_a_ex_o[30]));
 sky130_fd_sc_hd__buf_1 output626 (.A(net626),
    .X(multdiv_operand_a_ex_o[31]));
 sky130_fd_sc_hd__buf_1 output627 (.A(net627),
    .X(multdiv_operand_a_ex_o[3]));
 sky130_fd_sc_hd__buf_1 output628 (.A(net628),
    .X(multdiv_operand_a_ex_o[4]));
 sky130_fd_sc_hd__buf_1 output629 (.A(net629),
    .X(multdiv_operand_a_ex_o[5]));
 sky130_fd_sc_hd__buf_1 output630 (.A(net630),
    .X(multdiv_operand_a_ex_o[6]));
 sky130_fd_sc_hd__buf_1 output631 (.A(net631),
    .X(multdiv_operand_a_ex_o[7]));
 sky130_fd_sc_hd__buf_1 output632 (.A(net632),
    .X(multdiv_operand_a_ex_o[8]));
 sky130_fd_sc_hd__buf_1 output633 (.A(net633),
    .X(multdiv_operand_a_ex_o[9]));
 sky130_fd_sc_hd__buf_1 output634 (.A(net634),
    .X(multdiv_operand_b_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output635 (.A(net635),
    .X(multdiv_operand_b_ex_o[10]));
 sky130_fd_sc_hd__buf_1 output636 (.A(net636),
    .X(multdiv_operand_b_ex_o[11]));
 sky130_fd_sc_hd__buf_1 output637 (.A(net637),
    .X(multdiv_operand_b_ex_o[12]));
 sky130_fd_sc_hd__buf_1 output638 (.A(net638),
    .X(multdiv_operand_b_ex_o[13]));
 sky130_fd_sc_hd__buf_1 output639 (.A(net639),
    .X(multdiv_operand_b_ex_o[14]));
 sky130_fd_sc_hd__buf_1 output640 (.A(net640),
    .X(multdiv_operand_b_ex_o[15]));
 sky130_fd_sc_hd__buf_1 output641 (.A(net641),
    .X(multdiv_operand_b_ex_o[16]));
 sky130_fd_sc_hd__buf_1 output642 (.A(net642),
    .X(multdiv_operand_b_ex_o[17]));
 sky130_fd_sc_hd__buf_1 output643 (.A(net643),
    .X(multdiv_operand_b_ex_o[18]));
 sky130_fd_sc_hd__buf_1 output644 (.A(net644),
    .X(multdiv_operand_b_ex_o[19]));
 sky130_fd_sc_hd__buf_1 output645 (.A(net645),
    .X(multdiv_operand_b_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output646 (.A(net646),
    .X(multdiv_operand_b_ex_o[20]));
 sky130_fd_sc_hd__buf_1 output647 (.A(net647),
    .X(multdiv_operand_b_ex_o[21]));
 sky130_fd_sc_hd__buf_1 output648 (.A(net648),
    .X(multdiv_operand_b_ex_o[22]));
 sky130_fd_sc_hd__buf_1 output649 (.A(net649),
    .X(multdiv_operand_b_ex_o[23]));
 sky130_fd_sc_hd__buf_1 output650 (.A(net650),
    .X(multdiv_operand_b_ex_o[24]));
 sky130_fd_sc_hd__buf_1 output651 (.A(net651),
    .X(multdiv_operand_b_ex_o[25]));
 sky130_fd_sc_hd__buf_1 output652 (.A(net652),
    .X(multdiv_operand_b_ex_o[26]));
 sky130_fd_sc_hd__buf_1 output653 (.A(net653),
    .X(multdiv_operand_b_ex_o[27]));
 sky130_fd_sc_hd__buf_1 output654 (.A(net654),
    .X(multdiv_operand_b_ex_o[28]));
 sky130_fd_sc_hd__buf_1 output655 (.A(net655),
    .X(multdiv_operand_b_ex_o[29]));
 sky130_fd_sc_hd__buf_1 output656 (.A(net656),
    .X(multdiv_operand_b_ex_o[2]));
 sky130_fd_sc_hd__buf_1 output657 (.A(net657),
    .X(multdiv_operand_b_ex_o[30]));
 sky130_fd_sc_hd__buf_1 output658 (.A(net658),
    .X(multdiv_operand_b_ex_o[31]));
 sky130_fd_sc_hd__buf_1 output659 (.A(net659),
    .X(multdiv_operand_b_ex_o[3]));
 sky130_fd_sc_hd__buf_1 output660 (.A(net660),
    .X(multdiv_operand_b_ex_o[4]));
 sky130_fd_sc_hd__buf_1 output661 (.A(net661),
    .X(multdiv_operand_b_ex_o[5]));
 sky130_fd_sc_hd__buf_1 output662 (.A(net662),
    .X(multdiv_operand_b_ex_o[6]));
 sky130_fd_sc_hd__buf_1 output663 (.A(net663),
    .X(multdiv_operand_b_ex_o[7]));
 sky130_fd_sc_hd__buf_1 output664 (.A(net664),
    .X(multdiv_operand_b_ex_o[8]));
 sky130_fd_sc_hd__buf_1 output665 (.A(net665),
    .X(multdiv_operand_b_ex_o[9]));
 sky130_fd_sc_hd__buf_1 output666 (.A(net666),
    .X(multdiv_operator_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output667 (.A(net667),
    .X(multdiv_operator_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output668 (.A(net668),
    .X(multdiv_ready_id_o));
 sky130_fd_sc_hd__buf_1 output669 (.A(net669),
    .X(multdiv_signed_mode_ex_o[0]));
 sky130_fd_sc_hd__buf_1 output670 (.A(net670),
    .X(multdiv_signed_mode_ex_o[1]));
 sky130_fd_sc_hd__buf_1 output671 (.A(net671),
    .X(nmi_mode_o));
 sky130_fd_sc_hd__buf_1 output672 (.A(net672),
    .X(pc_mux_o[0]));
 sky130_fd_sc_hd__buf_1 output673 (.A(net673),
    .X(pc_mux_o[1]));
 sky130_fd_sc_hd__buf_1 output674 (.A(net674),
    .X(pc_mux_o[2]));
 sky130_fd_sc_hd__buf_1 output675 (.A(net675),
    .X(pc_set_o));
 sky130_fd_sc_hd__buf_1 output676 (.A(net676),
    .X(pc_set_spec_o));
 sky130_fd_sc_hd__buf_1 output677 (.A(net677),
    .X(perf_branch_o));
 sky130_fd_sc_hd__buf_1 output678 (.A(net678),
    .X(perf_div_wait_o));
 sky130_fd_sc_hd__buf_1 output679 (.A(net679),
    .X(perf_dside_wait_o));
 sky130_fd_sc_hd__buf_1 output680 (.A(net680),
    .X(perf_jump_o));
 sky130_fd_sc_hd__buf_1 output681 (.A(net681),
    .X(perf_mul_wait_o));
 sky130_fd_sc_hd__buf_1 output682 (.A(net682),
    .X(perf_tbranch_o));
 sky130_fd_sc_hd__buf_1 output683 (.A(net683),
    .X(rf_raddr_a_o[0]));
 sky130_fd_sc_hd__buf_1 output684 (.A(net684),
    .X(rf_raddr_a_o[1]));
 sky130_fd_sc_hd__buf_1 output685 (.A(net685),
    .X(rf_raddr_a_o[2]));
 sky130_fd_sc_hd__buf_1 output686 (.A(net686),
    .X(rf_raddr_a_o[3]));
 sky130_fd_sc_hd__buf_1 output687 (.A(net687),
    .X(rf_raddr_a_o[4]));
 sky130_fd_sc_hd__buf_1 output688 (.A(net688),
    .X(rf_raddr_b_o[0]));
 sky130_fd_sc_hd__buf_1 output689 (.A(net689),
    .X(rf_raddr_b_o[1]));
 sky130_fd_sc_hd__buf_1 output690 (.A(net690),
    .X(rf_raddr_b_o[2]));
 sky130_fd_sc_hd__buf_1 output691 (.A(net691),
    .X(rf_raddr_b_o[3]));
 sky130_fd_sc_hd__buf_1 output692 (.A(net692),
    .X(rf_raddr_b_o[4]));
 sky130_fd_sc_hd__buf_1 output693 (.A(net693),
    .X(rf_ren_a_o));
 sky130_fd_sc_hd__buf_1 output694 (.A(net694),
    .X(rf_ren_b_o));
 sky130_fd_sc_hd__buf_1 output695 (.A(net695),
    .X(rf_waddr_id_o[0]));
 sky130_fd_sc_hd__buf_1 output696 (.A(net696),
    .X(rf_waddr_id_o[1]));
 sky130_fd_sc_hd__buf_1 output697 (.A(net697),
    .X(rf_waddr_id_o[2]));
 sky130_fd_sc_hd__buf_1 output698 (.A(net698),
    .X(rf_waddr_id_o[3]));
 sky130_fd_sc_hd__buf_1 output699 (.A(net699),
    .X(rf_waddr_id_o[4]));
 sky130_fd_sc_hd__buf_1 output700 (.A(net700),
    .X(rf_wdata_id_o[0]));
 sky130_fd_sc_hd__buf_1 output701 (.A(net701),
    .X(rf_wdata_id_o[10]));
 sky130_fd_sc_hd__buf_1 output702 (.A(net702),
    .X(rf_wdata_id_o[11]));
 sky130_fd_sc_hd__buf_1 output703 (.A(net703),
    .X(rf_wdata_id_o[12]));
 sky130_fd_sc_hd__buf_1 output704 (.A(net704),
    .X(rf_wdata_id_o[13]));
 sky130_fd_sc_hd__buf_1 output705 (.A(net705),
    .X(rf_wdata_id_o[14]));
 sky130_fd_sc_hd__buf_1 output706 (.A(net706),
    .X(rf_wdata_id_o[15]));
 sky130_fd_sc_hd__buf_1 output707 (.A(net707),
    .X(rf_wdata_id_o[16]));
 sky130_fd_sc_hd__buf_1 output708 (.A(net708),
    .X(rf_wdata_id_o[17]));
 sky130_fd_sc_hd__buf_1 output709 (.A(net709),
    .X(rf_wdata_id_o[18]));
 sky130_fd_sc_hd__buf_1 output710 (.A(net710),
    .X(rf_wdata_id_o[19]));
 sky130_fd_sc_hd__buf_1 output711 (.A(net711),
    .X(rf_wdata_id_o[1]));
 sky130_fd_sc_hd__buf_1 output712 (.A(net712),
    .X(rf_wdata_id_o[20]));
 sky130_fd_sc_hd__buf_1 output713 (.A(net713),
    .X(rf_wdata_id_o[21]));
 sky130_fd_sc_hd__buf_1 output714 (.A(net714),
    .X(rf_wdata_id_o[22]));
 sky130_fd_sc_hd__buf_1 output715 (.A(net715),
    .X(rf_wdata_id_o[23]));
 sky130_fd_sc_hd__buf_1 output716 (.A(net716),
    .X(rf_wdata_id_o[24]));
 sky130_fd_sc_hd__buf_1 output717 (.A(net717),
    .X(rf_wdata_id_o[25]));
 sky130_fd_sc_hd__buf_1 output718 (.A(net718),
    .X(rf_wdata_id_o[26]));
 sky130_fd_sc_hd__buf_1 output719 (.A(net719),
    .X(rf_wdata_id_o[27]));
 sky130_fd_sc_hd__buf_1 output720 (.A(net720),
    .X(rf_wdata_id_o[28]));
 sky130_fd_sc_hd__buf_1 output721 (.A(net721),
    .X(rf_wdata_id_o[29]));
 sky130_fd_sc_hd__buf_1 output722 (.A(net722),
    .X(rf_wdata_id_o[2]));
 sky130_fd_sc_hd__buf_1 output723 (.A(net723),
    .X(rf_wdata_id_o[30]));
 sky130_fd_sc_hd__buf_1 output724 (.A(net724),
    .X(rf_wdata_id_o[31]));
 sky130_fd_sc_hd__buf_1 output725 (.A(net725),
    .X(rf_wdata_id_o[3]));
 sky130_fd_sc_hd__buf_1 output726 (.A(net726),
    .X(rf_wdata_id_o[4]));
 sky130_fd_sc_hd__buf_1 output727 (.A(net727),
    .X(rf_wdata_id_o[5]));
 sky130_fd_sc_hd__buf_1 output728 (.A(net728),
    .X(rf_wdata_id_o[6]));
 sky130_fd_sc_hd__buf_1 output729 (.A(net729),
    .X(rf_wdata_id_o[7]));
 sky130_fd_sc_hd__buf_1 output730 (.A(net730),
    .X(rf_wdata_id_o[8]));
 sky130_fd_sc_hd__buf_1 output731 (.A(net731),
    .X(rf_wdata_id_o[9]));
 sky130_fd_sc_hd__buf_1 output732 (.A(net732),
    .X(rf_we_id_o));
 sky130_fd_sc_hd__conb_1 _1925__733 (.LO(net733));
 sky130_fd_sc_hd__conb_1 _1926__734 (.LO(net734));
 sky130_fd_sc_hd__conb_1 _1927__735 (.LO(net735));
 sky130_fd_sc_hd__conb_1 _1928__736 (.LO(net736));
 sky130_fd_sc_hd__conb_1 _1929__737 (.LO(net737));
 sky130_fd_sc_hd__conb_1 _1930__738 (.LO(net738));
 sky130_fd_sc_hd__conb_1 _1931__739 (.LO(net739));
 sky130_fd_sc_hd__conb_1 _1932__740 (.LO(net740));
 sky130_fd_sc_hd__conb_1 _1933__741 (.LO(net741));
 sky130_fd_sc_hd__conb_1 _1934__742 (.LO(net742));
 sky130_fd_sc_hd__conb_1 _1935__743 (.LO(net743));
 sky130_fd_sc_hd__conb_1 _1936__744 (.LO(net744));
 sky130_fd_sc_hd__conb_1 _1937__745 (.LO(net745));
 sky130_fd_sc_hd__conb_1 _1938__746 (.LO(net746));
 sky130_fd_sc_hd__conb_1 _1939__747 (.LO(net747));
 sky130_fd_sc_hd__conb_1 _1940__748 (.LO(net748));
 sky130_fd_sc_hd__conb_1 _1941__749 (.LO(net749));
 sky130_fd_sc_hd__conb_1 _1942__750 (.LO(net750));
 sky130_fd_sc_hd__conb_1 _1943__751 (.LO(net751));
 sky130_fd_sc_hd__conb_1 _1944__752 (.LO(net752));
 sky130_fd_sc_hd__conb_1 _1945__753 (.LO(net753));
 sky130_fd_sc_hd__conb_1 _1946__754 (.LO(net754));
 sky130_fd_sc_hd__conb_1 _1947__755 (.LO(net755));
 sky130_fd_sc_hd__conb_1 _1948__756 (.LO(net756));
 sky130_fd_sc_hd__conb_1 _1949__757 (.LO(net757));
 sky130_fd_sc_hd__conb_1 _1950__758 (.LO(net758));
 sky130_fd_sc_hd__conb_1 _1951__759 (.LO(net759));
 sky130_fd_sc_hd__conb_1 _1952__760 (.LO(net760));
 sky130_fd_sc_hd__conb_1 _1953__761 (.LO(net761));
 sky130_fd_sc_hd__conb_1 _1954__762 (.LO(net762));
 sky130_fd_sc_hd__conb_1 _1955__763 (.LO(net763));
 sky130_fd_sc_hd__conb_1 _1956__764 (.LO(net764));
 sky130_fd_sc_hd__conb_1 _1957__765 (.LO(net765));
 sky130_fd_sc_hd__conb_1 _1958__766 (.LO(net766));
 sky130_fd_sc_hd__conb_1 _1959__767 (.LO(net767));
 sky130_fd_sc_hd__conb_1 _1960__768 (.LO(net768));
 sky130_fd_sc_hd__conb_1 _1961__769 (.LO(net769));
 sky130_fd_sc_hd__conb_1 _1962__770 (.LO(net770));
 sky130_fd_sc_hd__conb_1 _1963__771 (.LO(net771));
 sky130_fd_sc_hd__conb_1 _1964__772 (.LO(net772));
 sky130_fd_sc_hd__conb_1 _1965__773 (.LO(net773));
 sky130_fd_sc_hd__conb_1 _1966__774 (.LO(net774));
 sky130_fd_sc_hd__conb_1 _1967__775 (.LO(net775));
 sky130_fd_sc_hd__conb_1 _1968__776 (.LO(net776));
 sky130_fd_sc_hd__conb_1 _1969__777 (.LO(net777));
 sky130_fd_sc_hd__conb_1 _1970__778 (.LO(net778));
 sky130_fd_sc_hd__conb_1 _1971__779 (.LO(net779));
 sky130_fd_sc_hd__conb_1 _1972__780 (.LO(net780));
 sky130_fd_sc_hd__conb_1 _1973__781 (.LO(net781));
 sky130_fd_sc_hd__conb_1 _1974__782 (.LO(net782));
 sky130_fd_sc_hd__conb_1 _1975__783 (.LO(net783));
 sky130_fd_sc_hd__conb_1 _1976__784 (.LO(net784));
 sky130_fd_sc_hd__conb_1 _1977__785 (.LO(net785));
 sky130_fd_sc_hd__conb_1 _1978__786 (.LO(net786));
 sky130_fd_sc_hd__conb_1 _1979__787 (.LO(net787));
 sky130_fd_sc_hd__conb_1 _1980__788 (.LO(net788));
 sky130_fd_sc_hd__conb_1 _1981__789 (.LO(net789));
 sky130_fd_sc_hd__conb_1 _1982__790 (.LO(net790));
 sky130_fd_sc_hd__conb_1 _1983__791 (.LO(net791));
 sky130_fd_sc_hd__conb_1 _1984__792 (.LO(net792));
 sky130_fd_sc_hd__conb_1 _1985__793 (.LO(net793));
 sky130_fd_sc_hd__conb_1 _1986__794 (.LO(net794));
 sky130_fd_sc_hd__conb_1 _1987__795 (.LO(net795));
 sky130_fd_sc_hd__conb_1 _1988__796 (.LO(net796));
 sky130_fd_sc_hd__conb_1 _1989__797 (.LO(net797));
 sky130_fd_sc_hd__conb_1 _1991__798 (.LO(net798));
 sky130_fd_sc_hd__conb_1 _2090__799 (.LO(net799));
 sky130_fd_sc_hd__conb_1 _2102__800 (.LO(net800));
 sky130_fd_sc_hd__conb_1 _2103__801 (.LO(net801));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_6_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_3_0_0_clk_i));
 sky130_fd_sc_hd__inv_8 clkload1 (.A(clknet_3_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_3_2_0_clk_i));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload4 (.A(clknet_3_4_0_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload5 (.A(clknet_3_5_0_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_3_7_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net189));
 sky130_fd_sc_hd__fill_4 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_247_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_249_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_249_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_253_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_254_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_254_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_255_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_255_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_256_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_256_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_256_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_256_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_256_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_256_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_379 ();
endmodule
