module riscv_top (clk,
    memwrite,
    ready,
    reset,
    suspend,
    valid,
    valid_reg,
    dataadr,
    instr,
    pc,
    writedata);
 input clk;
 output memwrite;
 output ready;
 input reset;
 output suspend;
 input valid;
 input valid_reg;
 output [31:0] dataadr;
 input [31:0] instr;
 output [31:0] pc;
 output [31:0] writedata;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire clknet_leaf_0_clk;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire \readdata[0] ;
 wire \readdata[10] ;
 wire \readdata[11] ;
 wire \readdata[12] ;
 wire \readdata[13] ;
 wire \readdata[14] ;
 wire \readdata[15] ;
 wire \readdata[16] ;
 wire \readdata[17] ;
 wire \readdata[18] ;
 wire \readdata[19] ;
 wire \readdata[1] ;
 wire \readdata[20] ;
 wire \readdata[21] ;
 wire \readdata[22] ;
 wire \readdata[23] ;
 wire \readdata[24] ;
 wire \readdata[25] ;
 wire \readdata[26] ;
 wire \readdata[27] ;
 wire \readdata[28] ;
 wire \readdata[29] ;
 wire \readdata[2] ;
 wire \readdata[30] ;
 wire \readdata[31] ;
 wire \readdata[3] ;
 wire \readdata[4] ;
 wire \readdata[5] ;
 wire \readdata[6] ;
 wire \readdata[7] ;
 wire \readdata[8] ;
 wire \readdata[9] ;
 wire net97;
 wire \riscv.dp.ISRmux.d0[10] ;
 wire \riscv.dp.ISRmux.d0[11] ;
 wire \riscv.dp.ISRmux.d0[12] ;
 wire \riscv.dp.ISRmux.d0[13] ;
 wire \riscv.dp.ISRmux.d0[14] ;
 wire \riscv.dp.ISRmux.d0[15] ;
 wire \riscv.dp.ISRmux.d0[16] ;
 wire \riscv.dp.ISRmux.d0[17] ;
 wire \riscv.dp.ISRmux.d0[18] ;
 wire \riscv.dp.ISRmux.d0[19] ;
 wire \riscv.dp.ISRmux.d0[20] ;
 wire \riscv.dp.ISRmux.d0[21] ;
 wire \riscv.dp.ISRmux.d0[22] ;
 wire \riscv.dp.ISRmux.d0[23] ;
 wire \riscv.dp.ISRmux.d0[24] ;
 wire \riscv.dp.ISRmux.d0[25] ;
 wire \riscv.dp.ISRmux.d0[26] ;
 wire \riscv.dp.ISRmux.d0[27] ;
 wire \riscv.dp.ISRmux.d0[28] ;
 wire \riscv.dp.ISRmux.d0[29] ;
 wire \riscv.dp.ISRmux.d0[2] ;
 wire \riscv.dp.ISRmux.d0[30] ;
 wire \riscv.dp.ISRmux.d0[31] ;
 wire \riscv.dp.ISRmux.d0[3] ;
 wire \riscv.dp.ISRmux.d0[4] ;
 wire \riscv.dp.ISRmux.d0[5] ;
 wire \riscv.dp.ISRmux.d0[6] ;
 wire \riscv.dp.ISRmux.d0[7] ;
 wire \riscv.dp.ISRmux.d0[8] ;
 wire \riscv.dp.ISRmux.d0[9] ;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire \dmem/_000_ ;
 wire \dmem/_001_ ;
 wire \dmem/_002_ ;
 wire \dmem/_003_ ;
 wire \dmem/_004_ ;
 wire \dmem/_005_ ;
 wire \dmem/_006_ ;
 wire \dmem/_007_ ;
 wire \dmem/_008_ ;
 wire \dmem/_009_ ;
 wire \dmem/_010_ ;
 wire \dmem/_011_ ;
 wire \dmem/_012_ ;
 wire \dmem/_013_ ;
 wire \dmem/_014_ ;
 wire \dmem/_015_ ;
 wire \dmem/_016_ ;
 wire \dmem/_017_ ;
 wire \dmem/_018_ ;
 wire \dmem/_019_ ;
 wire \dmem/_020_ ;
 wire \dmem/_021_ ;
 wire \dmem/_022_ ;
 wire \dmem/_023_ ;
 wire \dmem/_024_ ;
 wire \dmem/_025_ ;
 wire \dmem/_026_ ;
 wire \dmem/_027_ ;
 wire \dmem/_028_ ;
 wire \dmem/_029_ ;
 wire \dmem/_030_ ;
 wire \dmem/_031_ ;
 wire \dmem/_032_ ;
 wire \dmem/_033_ ;
 wire \dmem/_034_ ;
 wire \dmem/_035_ ;
 wire \dmem/_036_ ;
 wire \dmem/_037_ ;
 wire \dmem/_038_ ;
 wire \dmem/_039_ ;
 wire \dmem/_040_ ;
 wire \dmem/_041_ ;
 wire \dmem/_042_ ;
 wire \dmem/_043_ ;
 wire \dmem/_044_ ;
 wire \dmem/_045_ ;
 wire \dmem/_046_ ;
 wire \dmem/_047_ ;
 wire \dmem/_048_ ;
 wire \dmem/_049_ ;
 wire \dmem/_050_ ;
 wire \dmem/_051_ ;
 wire \dmem/_052_ ;
 wire \dmem/_053_ ;
 wire \dmem/_054_ ;
 wire \dmem/_055_ ;
 wire \dmem/_056_ ;
 wire \dmem/_057_ ;
 wire \dmem/_058_ ;
 wire \dmem/_059_ ;
 wire \dmem/_060_ ;
 wire \dmem/_061_ ;
 wire \dmem/_062_ ;
 wire \dmem/_063_ ;
 wire \dmem/_064_ ;
 wire \dmem/_065_ ;
 wire \dmem/_066_ ;
 wire \dmem/_067_ ;
 wire \dmem/_068_ ;
 wire \dmem/_069_ ;
 wire \dmem/_070_ ;
 wire \dmem/_071_ ;
 wire \dmem/_072_ ;
 wire \dmem/_073_ ;
 wire \dmem/_074_ ;
 wire \dmem/_075_ ;
 wire \dmem/_076_ ;
 wire \dmem/_077_ ;
 wire \dmem/_078_ ;
 wire \dmem/_079_ ;
 wire \dmem/_080_ ;
 wire \dmem/_081_ ;
 wire \dmem/_082_ ;
 wire \dmem/_083_ ;
 wire \dmem/_084_ ;
 wire \dmem/_085_ ;
 wire \dmem/_086_ ;
 wire \dmem/_087_ ;
 wire \dmem/_088_ ;
 wire \dmem/_089_ ;
 wire \dmem/_090_ ;
 wire \dmem/_091_ ;
 wire \dmem/_092_ ;
 wire \dmem/_093_ ;
 wire \dmem/_094_ ;
 wire \dmem/_095_ ;
 wire \dmem/_096_ ;
 wire \dmem/_097_ ;
 wire \dmem/_098_ ;
 wire \dmem/_099_ ;
 wire \dmem/_100_ ;
 wire \dmem/_101_ ;
 wire \dmem/_102_ ;
 wire \dmem/_103_ ;
 wire \dmem/_104_ ;
 wire \dmem/_105_ ;
 wire \dmem/_106_ ;
 wire \dmem/_107_ ;
 wire \dmem/_108_ ;
 wire \dmem/_109_ ;
 wire \dmem/_110_ ;
 wire \dmem/_111_ ;
 wire \dmem/_112_ ;
 wire \dmem/_113_ ;
 wire \dmem/_114_ ;
 wire \dmem/_115_ ;
 wire \dmem/_116_ ;
 wire \dmem/_117_ ;
 wire \dmem/_118_ ;
 wire \dmem/_119_ ;
 wire \dmem/_120_ ;
 wire \dmem/_121_ ;
 wire \dmem/_122_ ;
 wire \dmem/_123_ ;
 wire \dmem/_124_ ;
 wire \dmem/_125_ ;
 wire \dmem/_126_ ;
 wire \dmem/_127_ ;
 wire \dmem/_128_ ;
 wire \dmem/_129_ ;
 wire \dmem/_130_ ;
 wire \dmem/_131_ ;
 wire \dmem/_132_ ;
 wire \dmem/_133_ ;
 wire \dmem/_134_ ;
 wire \dmem/_135_ ;
 wire \dmem/_136_ ;
 wire \dmem/_137_ ;
 wire \dmem/_138_ ;
 wire \dmem/_139_ ;
 wire \dmem/_140_ ;
 wire \dmem/_141_ ;
 wire \dmem/_142_ ;
 wire \dmem/_143_ ;
 wire \dmem/_144_ ;
 wire \dmem/_145_ ;
 wire \dmem/_146_ ;
 wire \dmem/_147_ ;
 wire \dmem/_148_ ;
 wire \dmem/_149_ ;
 wire \dmem/_150_ ;
 wire \dmem/_151_ ;
 wire \dmem/_152_ ;
 wire \dmem/ce_mem[0] ;
 wire \dmem/ce_mem[1] ;
 wire \dmem/ce_mem[2] ;
 wire \dmem/inter_dmem0[0] ;
 wire \dmem/inter_dmem0[10] ;
 wire \dmem/inter_dmem0[11] ;
 wire \dmem/inter_dmem0[12] ;
 wire \dmem/inter_dmem0[13] ;
 wire \dmem/inter_dmem0[14] ;
 wire \dmem/inter_dmem0[15] ;
 wire \dmem/inter_dmem0[16] ;
 wire \dmem/inter_dmem0[17] ;
 wire \dmem/inter_dmem0[18] ;
 wire \dmem/inter_dmem0[19] ;
 wire \dmem/inter_dmem0[1] ;
 wire \dmem/inter_dmem0[20] ;
 wire \dmem/inter_dmem0[21] ;
 wire \dmem/inter_dmem0[22] ;
 wire \dmem/inter_dmem0[23] ;
 wire \dmem/inter_dmem0[24] ;
 wire \dmem/inter_dmem0[25] ;
 wire \dmem/inter_dmem0[26] ;
 wire \dmem/inter_dmem0[27] ;
 wire \dmem/inter_dmem0[28] ;
 wire \dmem/inter_dmem0[29] ;
 wire \dmem/inter_dmem0[2] ;
 wire \dmem/inter_dmem0[30] ;
 wire \dmem/inter_dmem0[31] ;
 wire \dmem/inter_dmem0[3] ;
 wire \dmem/inter_dmem0[4] ;
 wire \dmem/inter_dmem0[5] ;
 wire \dmem/inter_dmem0[6] ;
 wire \dmem/inter_dmem0[7] ;
 wire \dmem/inter_dmem0[8] ;
 wire \dmem/inter_dmem0[9] ;
 wire \dmem/inter_dmem1[0] ;
 wire \dmem/inter_dmem1[10] ;
 wire \dmem/inter_dmem1[11] ;
 wire \dmem/inter_dmem1[12] ;
 wire \dmem/inter_dmem1[13] ;
 wire \dmem/inter_dmem1[14] ;
 wire \dmem/inter_dmem1[15] ;
 wire \dmem/inter_dmem1[16] ;
 wire \dmem/inter_dmem1[17] ;
 wire \dmem/inter_dmem1[18] ;
 wire \dmem/inter_dmem1[19] ;
 wire \dmem/inter_dmem1[1] ;
 wire \dmem/inter_dmem1[20] ;
 wire \dmem/inter_dmem1[21] ;
 wire \dmem/inter_dmem1[22] ;
 wire \dmem/inter_dmem1[23] ;
 wire \dmem/inter_dmem1[24] ;
 wire \dmem/inter_dmem1[25] ;
 wire \dmem/inter_dmem1[26] ;
 wire \dmem/inter_dmem1[27] ;
 wire \dmem/inter_dmem1[28] ;
 wire \dmem/inter_dmem1[29] ;
 wire \dmem/inter_dmem1[2] ;
 wire \dmem/inter_dmem1[30] ;
 wire \dmem/inter_dmem1[31] ;
 wire \dmem/inter_dmem1[3] ;
 wire \dmem/inter_dmem1[4] ;
 wire \dmem/inter_dmem1[5] ;
 wire \dmem/inter_dmem1[6] ;
 wire \dmem/inter_dmem1[7] ;
 wire \dmem/inter_dmem1[8] ;
 wire \dmem/inter_dmem1[9] ;
 wire \dmem/inter_dmem2[0] ;
 wire \dmem/inter_dmem2[10] ;
 wire \dmem/inter_dmem2[11] ;
 wire \dmem/inter_dmem2[12] ;
 wire \dmem/inter_dmem2[13] ;
 wire \dmem/inter_dmem2[14] ;
 wire \dmem/inter_dmem2[15] ;
 wire \dmem/inter_dmem2[16] ;
 wire \dmem/inter_dmem2[17] ;
 wire \dmem/inter_dmem2[18] ;
 wire \dmem/inter_dmem2[19] ;
 wire \dmem/inter_dmem2[1] ;
 wire \dmem/inter_dmem2[20] ;
 wire \dmem/inter_dmem2[21] ;
 wire \dmem/inter_dmem2[22] ;
 wire \dmem/inter_dmem2[23] ;
 wire \dmem/inter_dmem2[24] ;
 wire \dmem/inter_dmem2[25] ;
 wire \dmem/inter_dmem2[26] ;
 wire \dmem/inter_dmem2[27] ;
 wire \dmem/inter_dmem2[28] ;
 wire \dmem/inter_dmem2[29] ;
 wire \dmem/inter_dmem2[2] ;
 wire \dmem/inter_dmem2[30] ;
 wire \dmem/inter_dmem2[31] ;
 wire \dmem/inter_dmem2[3] ;
 wire \dmem/inter_dmem2[4] ;
 wire \dmem/inter_dmem2[5] ;
 wire \dmem/inter_dmem2[6] ;
 wire \dmem/inter_dmem2[7] ;
 wire \dmem/inter_dmem2[8] ;
 wire \dmem/inter_dmem2[9] ;
 wire \dmem/inter_dmem3[0] ;
 wire \dmem/inter_dmem3[10] ;
 wire \dmem/inter_dmem3[11] ;
 wire \dmem/inter_dmem3[12] ;
 wire \dmem/inter_dmem3[13] ;
 wire \dmem/inter_dmem3[14] ;
 wire \dmem/inter_dmem3[15] ;
 wire \dmem/inter_dmem3[16] ;
 wire \dmem/inter_dmem3[17] ;
 wire \dmem/inter_dmem3[18] ;
 wire \dmem/inter_dmem3[19] ;
 wire \dmem/inter_dmem3[1] ;
 wire \dmem/inter_dmem3[20] ;
 wire \dmem/inter_dmem3[21] ;
 wire \dmem/inter_dmem3[22] ;
 wire \dmem/inter_dmem3[23] ;
 wire \dmem/inter_dmem3[24] ;
 wire \dmem/inter_dmem3[25] ;
 wire \dmem/inter_dmem3[26] ;
 wire \dmem/inter_dmem3[27] ;
 wire \dmem/inter_dmem3[28] ;
 wire \dmem/inter_dmem3[29] ;
 wire \dmem/inter_dmem3[2] ;
 wire \dmem/inter_dmem3[30] ;
 wire \dmem/inter_dmem3[31] ;
 wire \dmem/inter_dmem3[3] ;
 wire \dmem/inter_dmem3[4] ;
 wire \dmem/inter_dmem3[5] ;
 wire \dmem/inter_dmem3[6] ;
 wire \dmem/inter_dmem3[7] ;
 wire \dmem/inter_dmem3[8] ;
 wire \dmem/inter_dmem3[9] ;
 wire \dmem/we_mem[0] ;
 wire \dmem/we_mem[1] ;
 wire \dmem/we_mem[2] ;
 wire \dmem/we_mem[3] ;
 wire net3;
 wire net4;
 wire net1;
 wire net2;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;

 CKINVDCx10_ASAP7_75t_R _09778_ (.A(net168),
    .Y(_03016_));
 BUFx12f_ASAP7_75t_R _09779_ (.A(_03016_),
    .Y(_03017_));
 BUFx16f_ASAP7_75t_R _09780_ (.A(_03017_),
    .Y(_03018_));
 BUFx12_ASAP7_75t_R _09781_ (.A(_03018_),
    .Y(_03019_));
 BUFx6f_ASAP7_75t_R _09782_ (.A(_03019_),
    .Y(_03020_));
 BUFx12f_ASAP7_75t_R _09783_ (.A(_03020_),
    .Y(_03021_));
 BUFx10_ASAP7_75t_R _09784_ (.A(_03021_),
    .Y(_03022_));
 BUFx6f_ASAP7_75t_R _09785_ (.A(_03022_),
    .Y(_03023_));
 BUFx6f_ASAP7_75t_R _09786_ (.A(_03023_),
    .Y(_03024_));
 BUFx10_ASAP7_75t_R _09787_ (.A(_03024_),
    .Y(_03025_));
 BUFx4f_ASAP7_75t_R _09788_ (.A(_03025_),
    .Y(net89));
 INVx5_ASAP7_75t_R _09789_ (.A(net12),
    .Y(_03026_));
 BUFx12f_ASAP7_75t_R _09790_ (.A(_03026_),
    .Y(_03027_));
 BUFx6f_ASAP7_75t_R _09791_ (.A(_03027_),
    .Y(_03028_));
 BUFx10_ASAP7_75t_R _09792_ (.A(_03028_),
    .Y(_03029_));
 INVx1_ASAP7_75t_R _09793_ (.A(_00023_),
    .Y(_03030_));
 BUFx10_ASAP7_75t_R _09794_ (.A(_03018_),
    .Y(_03031_));
 NAND2x2_ASAP7_75t_R _09795_ (.A(net15),
    .B(_03031_),
    .Y(_03032_));
 BUFx6f_ASAP7_75t_R _09796_ (.A(net15),
    .Y(_03033_));
 BUFx6f_ASAP7_75t_R _09797_ (.A(_03019_),
    .Y(_03034_));
 INVx2_ASAP7_75t_R _09798_ (.A(_00007_),
    .Y(_03035_));
 AO21x1_ASAP7_75t_R _09799_ (.A1(_03033_),
    .A2(_03034_),
    .B(_03035_),
    .Y(_03036_));
 BUFx6f_ASAP7_75t_R _09800_ (.A(instr[20]),
    .Y(_03037_));
 BUFx6f_ASAP7_75t_R _09801_ (.A(_03037_),
    .Y(_03038_));
 BUFx6f_ASAP7_75t_R _09802_ (.A(_03038_),
    .Y(_03039_));
 BUFx10_ASAP7_75t_R _09803_ (.A(_03039_),
    .Y(_03040_));
 BUFx10_ASAP7_75t_R _09804_ (.A(_03040_),
    .Y(_03041_));
 OA211x2_ASAP7_75t_R _09805_ (.A1(_03030_),
    .A2(_03032_),
    .B(_03036_),
    .C(_03041_),
    .Y(_03042_));
 BUFx10_ASAP7_75t_R _09806_ (.A(_03018_),
    .Y(_03043_));
 BUFx12f_ASAP7_75t_R _09807_ (.A(_03043_),
    .Y(_03044_));
 BUFx12f_ASAP7_75t_R _09808_ (.A(_03044_),
    .Y(_03045_));
 AND3x1_ASAP7_75t_R _09809_ (.A(_03033_),
    .B(_00022_),
    .C(_03045_),
    .Y(_03046_));
 BUFx10_ASAP7_75t_R _09810_ (.A(_03038_),
    .Y(_03047_));
 BUFx10_ASAP7_75t_R _09811_ (.A(_03047_),
    .Y(_03048_));
 BUFx6f_ASAP7_75t_R _09812_ (.A(_03048_),
    .Y(_03049_));
 AOI211x1_ASAP7_75t_R _09813_ (.A1(_00006_),
    .A2(_03032_),
    .B(_03046_),
    .C(_03049_),
    .Y(_03050_));
 OR3x1_ASAP7_75t_R _09814_ (.A(_03029_),
    .B(_03042_),
    .C(_03050_),
    .Y(_03051_));
 INVx5_ASAP7_75t_R _09815_ (.A(net13),
    .Y(_03052_));
 INVx4_ASAP7_75t_R _09816_ (.A(_03037_),
    .Y(_03053_));
 BUFx6f_ASAP7_75t_R _09817_ (.A(_03053_),
    .Y(_03054_));
 BUFx10_ASAP7_75t_R _09818_ (.A(_03054_),
    .Y(_03055_));
 BUFx10_ASAP7_75t_R _09819_ (.A(_03055_),
    .Y(_03056_));
 BUFx6f_ASAP7_75t_R _09820_ (.A(_03038_),
    .Y(_03057_));
 BUFx6f_ASAP7_75t_R _09821_ (.A(_03057_),
    .Y(_03058_));
 AND2x2_ASAP7_75t_R _09822_ (.A(_03058_),
    .B(_00021_),
    .Y(_03059_));
 AO21x1_ASAP7_75t_R _09823_ (.A1(_03056_),
    .A2(_00020_),
    .B(_03059_),
    .Y(_03060_));
 BUFx12_ASAP7_75t_R _09824_ (.A(_03053_),
    .Y(_03061_));
 BUFx12_ASAP7_75t_R _09825_ (.A(_03061_),
    .Y(_03062_));
 BUFx12f_ASAP7_75t_R _09826_ (.A(_03043_),
    .Y(_03063_));
 BUFx12f_ASAP7_75t_R _09827_ (.A(_03063_),
    .Y(_03064_));
 BUFx6f_ASAP7_75t_R _09828_ (.A(_03057_),
    .Y(_03065_));
 AO21x1_ASAP7_75t_R _09829_ (.A1(_03065_),
    .A2(_00005_),
    .B(net15),
    .Y(_03066_));
 AO22x1_ASAP7_75t_R _09830_ (.A1(_03062_),
    .A2(_00004_),
    .B1(_03064_),
    .B2(_03066_),
    .Y(_03067_));
 BUFx10_ASAP7_75t_R _09831_ (.A(_03027_),
    .Y(_03068_));
 OA211x2_ASAP7_75t_R _09832_ (.A1(_03032_),
    .A2(_03060_),
    .B(_03067_),
    .C(_03068_),
    .Y(_03069_));
 NOR2x1_ASAP7_75t_R _09833_ (.A(_03052_),
    .B(_03069_),
    .Y(_03070_));
 BUFx6f_ASAP7_75t_R _09834_ (.A(_03048_),
    .Y(_03071_));
 BUFx10_ASAP7_75t_R _09835_ (.A(net12),
    .Y(_03072_));
 BUFx6f_ASAP7_75t_R _09836_ (.A(_03072_),
    .Y(_03073_));
 BUFx12_ASAP7_75t_R _09837_ (.A(_03073_),
    .Y(_03074_));
 OR2x2_ASAP7_75t_R _09838_ (.A(_03071_),
    .B(_03074_),
    .Y(_03075_));
 INVx1_ASAP7_75t_R _09839_ (.A(_00000_),
    .Y(_01222_));
 AO21x1_ASAP7_75t_R _09840_ (.A1(_03022_),
    .A2(_03075_),
    .B(_01222_),
    .Y(_03076_));
 BUFx10_ASAP7_75t_R _09841_ (.A(net13),
    .Y(_03077_));
 BUFx6f_ASAP7_75t_R _09842_ (.A(_03077_),
    .Y(_03078_));
 NOR2x1_ASAP7_75t_R _09843_ (.A(_03078_),
    .B(_03033_),
    .Y(_03079_));
 BUFx12_ASAP7_75t_R _09844_ (.A(_03053_),
    .Y(_03080_));
 BUFx10_ASAP7_75t_R _09845_ (.A(_03080_),
    .Y(_03081_));
 BUFx10_ASAP7_75t_R _09846_ (.A(_03081_),
    .Y(_03082_));
 NAND2x1_ASAP7_75t_R _09847_ (.A(_03074_),
    .B(_00002_),
    .Y(_03083_));
 INVx1_ASAP7_75t_R _09848_ (.A(_00001_),
    .Y(_03084_));
 BUFx6f_ASAP7_75t_R _09849_ (.A(net12),
    .Y(_03085_));
 BUFx10_ASAP7_75t_R _09850_ (.A(_03085_),
    .Y(_03086_));
 BUFx12f_ASAP7_75t_R _09851_ (.A(_03086_),
    .Y(_03087_));
 BUFx6f_ASAP7_75t_R _09852_ (.A(_03085_),
    .Y(_03088_));
 NAND2x1_ASAP7_75t_R _09853_ (.A(_03088_),
    .B(_00003_),
    .Y(_03089_));
 BUFx12_ASAP7_75t_R _09854_ (.A(_03037_),
    .Y(_03090_));
 BUFx12_ASAP7_75t_R _09855_ (.A(_03090_),
    .Y(_03091_));
 BUFx10_ASAP7_75t_R _09856_ (.A(_03091_),
    .Y(_03092_));
 OA211x2_ASAP7_75t_R _09857_ (.A1(_03084_),
    .A2(_03087_),
    .B(_03089_),
    .C(_03092_),
    .Y(_03093_));
 AO21x1_ASAP7_75t_R _09858_ (.A1(_03082_),
    .A2(_03083_),
    .B(_03093_),
    .Y(_03094_));
 BUFx16f_ASAP7_75t_R _09859_ (.A(net168),
    .Y(_03095_));
 BUFx16f_ASAP7_75t_R _09860_ (.A(_03095_),
    .Y(_03096_));
 BUFx12f_ASAP7_75t_R _09861_ (.A(_03096_),
    .Y(_03097_));
 BUFx10_ASAP7_75t_R _09862_ (.A(_03097_),
    .Y(_03098_));
 BUFx10_ASAP7_75t_R _09863_ (.A(_03098_),
    .Y(_03099_));
 AO21x1_ASAP7_75t_R _09864_ (.A1(_03079_),
    .A2(_03094_),
    .B(_03099_),
    .Y(_03100_));
 INVx1_ASAP7_75t_R _09865_ (.A(_00019_),
    .Y(_03101_));
 INVx1_ASAP7_75t_R _09866_ (.A(_00017_),
    .Y(_03102_));
 BUFx12f_ASAP7_75t_R _09867_ (.A(_03095_),
    .Y(_03103_));
 BUFx12f_ASAP7_75t_R _09868_ (.A(_03103_),
    .Y(_03104_));
 OR3x1_ASAP7_75t_R _09869_ (.A(_03073_),
    .B(_03102_),
    .C(_03104_),
    .Y(_03105_));
 OA211x2_ASAP7_75t_R _09870_ (.A1(_03028_),
    .A2(_03101_),
    .B(_03105_),
    .C(_03041_),
    .Y(_03106_));
 BUFx12_ASAP7_75t_R _09871_ (.A(_03073_),
    .Y(_03107_));
 INVx1_ASAP7_75t_R _09872_ (.A(_00016_),
    .Y(_03108_));
 BUFx10_ASAP7_75t_R _09873_ (.A(_03086_),
    .Y(_03109_));
 NAND2x1_ASAP7_75t_R _09874_ (.A(_03109_),
    .B(_00018_),
    .Y(_03110_));
 BUFx10_ASAP7_75t_R _09875_ (.A(_03054_),
    .Y(_03111_));
 BUFx10_ASAP7_75t_R _09876_ (.A(_03111_),
    .Y(_03112_));
 OA211x2_ASAP7_75t_R _09877_ (.A1(_03107_),
    .A2(_03108_),
    .B(_03110_),
    .C(_03112_),
    .Y(_03113_));
 OA211x2_ASAP7_75t_R _09878_ (.A1(_03106_),
    .A2(_03113_),
    .B(_03052_),
    .C(_03033_),
    .Y(_03114_));
 AO221x1_ASAP7_75t_R _09879_ (.A1(_03051_),
    .A2(_03070_),
    .B1(_03076_),
    .B2(_03100_),
    .C(_03114_),
    .Y(_03115_));
 BUFx10_ASAP7_75t_R _09880_ (.A(_03017_),
    .Y(_03116_));
 BUFx6f_ASAP7_75t_R _09881_ (.A(_03116_),
    .Y(_03117_));
 AND2x6_ASAP7_75t_R _09882_ (.A(net14),
    .B(_03117_),
    .Y(_03118_));
 BUFx12_ASAP7_75t_R _09883_ (.A(_03118_),
    .Y(_03119_));
 NAND2x2_ASAP7_75t_R _09884_ (.A(net14),
    .B(_03019_),
    .Y(_03120_));
 NAND2x2_ASAP7_75t_R _09885_ (.A(net12),
    .B(_03116_),
    .Y(_03121_));
 NAND2x2_ASAP7_75t_R _09886_ (.A(_03037_),
    .B(_03018_),
    .Y(_03122_));
 BUFx10_ASAP7_75t_R _09887_ (.A(_03122_),
    .Y(_03123_));
 NAND2x2_ASAP7_75t_R _09888_ (.A(net13),
    .B(_03018_),
    .Y(_03124_));
 BUFx6f_ASAP7_75t_R _09889_ (.A(_03124_),
    .Y(_03125_));
 AND5x2_ASAP7_75t_R _09890_ (.A(_03032_),
    .B(_03120_),
    .C(_03121_),
    .D(_03123_),
    .E(_03125_),
    .Y(_03126_));
 BUFx10_ASAP7_75t_R _09891_ (.A(_03126_),
    .Y(_03127_));
 NOR2x2_ASAP7_75t_R _09892_ (.A(_03119_),
    .B(_03127_),
    .Y(_03128_));
 INVx2_ASAP7_75t_R _09893_ (.A(_00008_),
    .Y(_03129_));
 BUFx10_ASAP7_75t_R _09894_ (.A(_03096_),
    .Y(_03130_));
 BUFx6f_ASAP7_75t_R _09895_ (.A(_03130_),
    .Y(_03131_));
 BUFx12f_ASAP7_75t_R _09896_ (.A(_03027_),
    .Y(_03132_));
 AND2x2_ASAP7_75t_R _09897_ (.A(_03058_),
    .B(_00011_),
    .Y(_03133_));
 AOI21x1_ASAP7_75t_R _09898_ (.A1(_03056_),
    .A2(_00010_),
    .B(_03133_),
    .Y(_03134_));
 OA211x2_ASAP7_75t_R _09899_ (.A1(_03132_),
    .A2(_03134_),
    .B(_03021_),
    .C(_03052_),
    .Y(_03135_));
 AO21x1_ASAP7_75t_R _09900_ (.A1(_03129_),
    .A2(_03131_),
    .B(_03135_),
    .Y(_03136_));
 BUFx6f_ASAP7_75t_R _09901_ (.A(_03132_),
    .Y(_03137_));
 BUFx6f_ASAP7_75t_R _09902_ (.A(_03055_),
    .Y(_03138_));
 BUFx10_ASAP7_75t_R _09903_ (.A(_03138_),
    .Y(_03139_));
 AND3x1_ASAP7_75t_R _09904_ (.A(_03041_),
    .B(_00009_),
    .C(_03021_),
    .Y(_03140_));
 AO21x1_ASAP7_75t_R _09905_ (.A1(_03139_),
    .A2(_00008_),
    .B(_03140_),
    .Y(_03141_));
 AND2x6_ASAP7_75t_R _09906_ (.A(_03033_),
    .B(_03064_),
    .Y(_03142_));
 BUFx12f_ASAP7_75t_R _09907_ (.A(_03142_),
    .Y(_03143_));
 AOI21x1_ASAP7_75t_R _09908_ (.A1(_03137_),
    .A2(_03141_),
    .B(_03143_),
    .Y(_03144_));
 BUFx6f_ASAP7_75t_R _09909_ (.A(_03044_),
    .Y(_03145_));
 AND3x1_ASAP7_75t_R _09910_ (.A(_03033_),
    .B(_00030_),
    .C(_03145_),
    .Y(_03146_));
 AOI211x1_ASAP7_75t_R _09911_ (.A1(_00014_),
    .A2(_03032_),
    .B(_03146_),
    .C(_03049_),
    .Y(_03147_));
 INVx3_ASAP7_75t_R _09912_ (.A(_00031_),
    .Y(_03148_));
 BUFx12_ASAP7_75t_R _09913_ (.A(_03117_),
    .Y(_03149_));
 INVx2_ASAP7_75t_R _09914_ (.A(_00015_),
    .Y(_03150_));
 AO21x1_ASAP7_75t_R _09915_ (.A1(_03033_),
    .A2(_03149_),
    .B(_03150_),
    .Y(_03151_));
 OA211x2_ASAP7_75t_R _09916_ (.A1(_03148_),
    .A2(_03032_),
    .B(_03151_),
    .C(_03041_),
    .Y(_03152_));
 OR3x1_ASAP7_75t_R _09917_ (.A(_03029_),
    .B(_03147_),
    .C(_03152_),
    .Y(_03153_));
 BUFx12f_ASAP7_75t_R _09918_ (.A(_03032_),
    .Y(_03154_));
 BUFx10_ASAP7_75t_R _09919_ (.A(_03057_),
    .Y(_03155_));
 AND2x2_ASAP7_75t_R _09920_ (.A(_03155_),
    .B(_00029_),
    .Y(_03156_));
 AO21x1_ASAP7_75t_R _09921_ (.A1(_03056_),
    .A2(_00028_),
    .B(_03156_),
    .Y(_03157_));
 AO21x1_ASAP7_75t_R _09922_ (.A1(_03058_),
    .A2(_00013_),
    .B(_03033_),
    .Y(_03158_));
 AO22x1_ASAP7_75t_R _09923_ (.A1(_03081_),
    .A2(_00012_),
    .B1(_03045_),
    .B2(_03158_),
    .Y(_03159_));
 BUFx12_ASAP7_75t_R _09924_ (.A(_03026_),
    .Y(_03160_));
 BUFx12f_ASAP7_75t_R _09925_ (.A(_03160_),
    .Y(_03161_));
 OA211x2_ASAP7_75t_R _09926_ (.A1(_03154_),
    .A2(_03157_),
    .B(_03159_),
    .C(_03161_),
    .Y(_03162_));
 NOR2x1_ASAP7_75t_R _09927_ (.A(_03052_),
    .B(_03162_),
    .Y(_03163_));
 INVx3_ASAP7_75t_R _09928_ (.A(_00027_),
    .Y(_03164_));
 INVx3_ASAP7_75t_R _09929_ (.A(_00025_),
    .Y(_03165_));
 OR3x1_ASAP7_75t_R _09930_ (.A(_03073_),
    .B(_03165_),
    .C(_03104_),
    .Y(_03166_));
 OA211x2_ASAP7_75t_R _09931_ (.A1(_03028_),
    .A2(_03164_),
    .B(_03166_),
    .C(_03041_),
    .Y(_03167_));
 INVx3_ASAP7_75t_R _09932_ (.A(_00024_),
    .Y(_03168_));
 NAND2x1_ASAP7_75t_R _09933_ (.A(_03109_),
    .B(_00026_),
    .Y(_03169_));
 OA211x2_ASAP7_75t_R _09934_ (.A1(_03107_),
    .A2(_03168_),
    .B(_03169_),
    .C(_03112_),
    .Y(_03170_));
 OA211x2_ASAP7_75t_R _09935_ (.A1(_03167_),
    .A2(_03170_),
    .B(_03052_),
    .C(_03033_),
    .Y(_03171_));
 AO221x1_ASAP7_75t_R _09936_ (.A1(_03136_),
    .A2(_03144_),
    .B1(_03153_),
    .B2(_03163_),
    .C(_03171_),
    .Y(_03172_));
 BUFx6f_ASAP7_75t_R _09937_ (.A(_03118_),
    .Y(_03173_));
 BUFx6f_ASAP7_75t_R _09938_ (.A(_03173_),
    .Y(_03174_));
 BUFx6f_ASAP7_75t_R _09939_ (.A(_03174_),
    .Y(_03175_));
 AOI22x1_ASAP7_75t_R _09940_ (.A1(_03115_),
    .A2(_03128_),
    .B1(_03172_),
    .B2(_03175_),
    .Y(_03176_));
 CKINVDCx20_ASAP7_75t_R _09941_ (.A(_03176_),
    .Y(net99));
 INVx3_ASAP7_75t_R _09942_ (.A(_01114_),
    .Y(net73));
 INVx2_ASAP7_75t_R _09943_ (.A(_01111_),
    .Y(net72));
 INVx2_ASAP7_75t_R _09944_ (.A(_01120_),
    .Y(net75));
 INVx3_ASAP7_75t_R _09945_ (.A(_01117_),
    .Y(net74));
 INVx3_ASAP7_75t_R _09946_ (.A(_01126_),
    .Y(net78));
 INVx3_ASAP7_75t_R _09947_ (.A(_01123_),
    .Y(net77));
 INVx2_ASAP7_75t_R _09948_ (.A(_01132_),
    .Y(net80));
 INVx3_ASAP7_75t_R _09949_ (.A(_01129_),
    .Y(net79));
 INVx3_ASAP7_75t_R _09950_ (.A(_01138_),
    .Y(net82));
 INVx2_ASAP7_75t_R _09951_ (.A(_01135_),
    .Y(net81));
 INVx2_ASAP7_75t_R _09952_ (.A(_01144_),
    .Y(net84));
 INVx3_ASAP7_75t_R _09953_ (.A(_01141_),
    .Y(net83));
 INVx3_ASAP7_75t_R _09954_ (.A(_01150_),
    .Y(net86));
 INVx2_ASAP7_75t_R _09955_ (.A(_01147_),
    .Y(net85));
 INVx2_ASAP7_75t_R _09956_ (.A(_01153_),
    .Y(net88));
 INVx3_ASAP7_75t_R _09957_ (.A(_01090_),
    .Y(net96));
 INVx3_ASAP7_75t_R _09958_ (.A(_01087_),
    .Y(net95));
 INVx3_ASAP7_75t_R _09959_ (.A(_01096_),
    .Y(net67));
 INVx3_ASAP7_75t_R _09960_ (.A(_01093_),
    .Y(net66));
 INVx3_ASAP7_75t_R _09961_ (.A(_01102_),
    .Y(net69));
 INVx3_ASAP7_75t_R _09962_ (.A(_01099_),
    .Y(net68));
 INVx3_ASAP7_75t_R _09963_ (.A(_01108_),
    .Y(net71));
 INVx3_ASAP7_75t_R _09964_ (.A(_01105_),
    .Y(net70));
 INVx3_ASAP7_75t_R _09965_ (.A(_01078_),
    .Y(net92));
 INVx2_ASAP7_75t_R _09966_ (.A(_01075_),
    .Y(net91));
 INVx2_ASAP7_75t_R _09967_ (.A(_01084_),
    .Y(net94));
 INVx2_ASAP7_75t_R _09968_ (.A(_01081_),
    .Y(net93));
 INVx3_ASAP7_75t_R _09969_ (.A(_01068_),
    .Y(net76));
 INVx2_ASAP7_75t_R _09970_ (.A(_01066_),
    .Y(net65));
 NAND2x2_ASAP7_75t_R _09971_ (.A(net1),
    .B(net11),
    .Y(_03177_));
 AND2x2_ASAP7_75t_R _09972_ (.A(_00032_),
    .B(_00033_),
    .Y(_03178_));
 AND4x2_ASAP7_75t_R _09973_ (.A(_01132_),
    .B(_01135_),
    .C(_01138_),
    .D(_01153_),
    .Y(_03179_));
 AND4x2_ASAP7_75t_R _09974_ (.A(_01141_),
    .B(_01144_),
    .C(_01147_),
    .D(_01150_),
    .Y(_03180_));
 NAND2x1_ASAP7_75t_R _09975_ (.A(_03179_),
    .B(_03180_),
    .Y(_03181_));
 AND4x2_ASAP7_75t_R _09976_ (.A(_01157_),
    .B(_01111_),
    .C(_01114_),
    .D(_01129_),
    .Y(_03182_));
 AND4x2_ASAP7_75t_R _09977_ (.A(_01117_),
    .B(_01120_),
    .C(_01123_),
    .D(_01126_),
    .Y(_03183_));
 NAND2x1_ASAP7_75t_R _09978_ (.A(_03182_),
    .B(_03183_),
    .Y(_03184_));
 AND4x1_ASAP7_75t_R _09979_ (.A(_01084_),
    .B(_01090_),
    .C(_01093_),
    .D(_01108_),
    .Y(_03185_));
 AND4x1_ASAP7_75t_R _09980_ (.A(_01096_),
    .B(_01099_),
    .C(_01102_),
    .D(_01105_),
    .Y(_03186_));
 NAND2x1_ASAP7_75t_R _09981_ (.A(_03185_),
    .B(_03186_),
    .Y(_03187_));
 AND4x2_ASAP7_75t_R _09982_ (.A(_01068_),
    .B(_01075_),
    .C(_01078_),
    .D(_01081_),
    .Y(_03188_));
 AND2x2_ASAP7_75t_R _09983_ (.A(_01066_),
    .B(_01087_),
    .Y(_03189_));
 NAND2x1_ASAP7_75t_R _09984_ (.A(_03188_),
    .B(_03189_),
    .Y(_03190_));
 OR5x1_ASAP7_75t_R _09985_ (.A(_03178_),
    .B(_03181_),
    .C(_03184_),
    .D(_03187_),
    .E(_03190_),
    .Y(_03191_));
 BUFx3_ASAP7_75t_R _09986_ (.A(_03191_),
    .Y(_03192_));
 OR5x2_ASAP7_75t_R _09987_ (.A(_00032_),
    .B(_03181_),
    .C(_03184_),
    .D(_03187_),
    .E(_03190_),
    .Y(_03193_));
 INVx2_ASAP7_75t_R _09988_ (.A(net25),
    .Y(_03194_));
 INVx1_ASAP7_75t_R _09989_ (.A(net26),
    .Y(_03195_));
 OR3x1_ASAP7_75t_R _09990_ (.A(_03131_),
    .B(_03194_),
    .C(_03195_),
    .Y(_03196_));
 BUFx12_ASAP7_75t_R _09991_ (.A(net24),
    .Y(_03197_));
 OR3x2_ASAP7_75t_R _09992_ (.A(_03095_),
    .B(net21),
    .C(_03197_),
    .Y(_03198_));
 AOI221x1_ASAP7_75t_R _09993_ (.A1(_03177_),
    .A2(_03192_),
    .B1(_03193_),
    .B2(_03196_),
    .C(_03198_),
    .Y(_03199_));
 BUFx12_ASAP7_75t_R _09994_ (.A(_03044_),
    .Y(_03200_));
 BUFx12f_ASAP7_75t_R _09995_ (.A(_03200_),
    .Y(_03201_));
 NAND2x2_ASAP7_75t_R _09996_ (.A(_03201_),
    .B(net27),
    .Y(_03202_));
 INVx1_ASAP7_75t_R _09997_ (.A(_00033_),
    .Y(_03203_));
 NAND2x1_ASAP7_75t_R _09998_ (.A(_00032_),
    .B(_03203_),
    .Y(_03204_));
 OR5x2_ASAP7_75t_R _09999_ (.A(_03181_),
    .B(_03184_),
    .C(_03187_),
    .D(_03190_),
    .E(_03204_),
    .Y(_03205_));
 BUFx6f_ASAP7_75t_R _10000_ (.A(_03205_),
    .Y(_03206_));
 BUFx6f_ASAP7_75t_R _10001_ (.A(_03206_),
    .Y(_03207_));
 BUFx6f_ASAP7_75t_R _10002_ (.A(_03207_),
    .Y(_03208_));
 BUFx16f_ASAP7_75t_R _10003_ (.A(_03208_),
    .Y(_03209_));
 BUFx10_ASAP7_75t_R _10004_ (.A(_03209_),
    .Y(_03210_));
 AND3x1_ASAP7_75t_R _10005_ (.A(net22),
    .B(_03202_),
    .C(_03210_),
    .Y(_03211_));
 BUFx4f_ASAP7_75t_R _10006_ (.A(instr[13]),
    .Y(_03212_));
 INVx1_ASAP7_75t_R _10007_ (.A(_03212_),
    .Y(_03213_));
 AOI21x1_ASAP7_75t_R _10008_ (.A1(_03199_),
    .A2(_03211_),
    .B(_03213_),
    .Y(_03214_));
 BUFx10_ASAP7_75t_R _10009_ (.A(_03149_),
    .Y(_03215_));
 BUFx6f_ASAP7_75t_R _10010_ (.A(_03215_),
    .Y(_03216_));
 BUFx4f_ASAP7_75t_R _10011_ (.A(instr[12]),
    .Y(_03217_));
 NAND2x2_ASAP7_75t_R _10012_ (.A(_03216_),
    .B(_03217_),
    .Y(_03218_));
 AND4x1_ASAP7_75t_R _10013_ (.A(_03213_),
    .B(_03199_),
    .C(_03211_),
    .D(_03218_),
    .Y(_03219_));
 NOR2x1_ASAP7_75t_R _10014_ (.A(_03214_),
    .B(_03219_),
    .Y(_03220_));
 OR3x1_ASAP7_75t_R _10015_ (.A(_03103_),
    .B(net27),
    .C(net26),
    .Y(_03221_));
 AOI211x1_ASAP7_75t_R _10016_ (.A1(_03177_),
    .A2(_03192_),
    .B(_03198_),
    .C(_03221_),
    .Y(_03222_));
 OA21x2_ASAP7_75t_R _10017_ (.A1(_03099_),
    .A2(_03194_),
    .B(_03193_),
    .Y(_03223_));
 BUFx4f_ASAP7_75t_R _10018_ (.A(_03223_),
    .Y(_03224_));
 BUFx6f_ASAP7_75t_R _10019_ (.A(_03197_),
    .Y(_03225_));
 BUFx12_ASAP7_75t_R _10020_ (.A(_03225_),
    .Y(_03226_));
 OR3x2_ASAP7_75t_R _10021_ (.A(_03103_),
    .B(net25),
    .C(_03195_),
    .Y(_03227_));
 OR5x1_ASAP7_75t_R _10022_ (.A(_03130_),
    .B(net21),
    .C(_03226_),
    .D(net27),
    .E(_03227_),
    .Y(_03228_));
 AO21x2_ASAP7_75t_R _10023_ (.A1(_03177_),
    .A2(_03192_),
    .B(_03228_),
    .Y(_03229_));
 INVx13_ASAP7_75t_R _10024_ (.A(_03229_),
    .Y(net64));
 AO21x1_ASAP7_75t_R _10025_ (.A1(_03222_),
    .A2(_03224_),
    .B(net64),
    .Y(_03230_));
 OR3x4_ASAP7_75t_R _10026_ (.A(_03095_),
    .B(net27),
    .C(_03194_),
    .Y(_03231_));
 NAND2x2_ASAP7_75t_R _10027_ (.A(_03193_),
    .B(_03231_),
    .Y(_03232_));
 BUFx6f_ASAP7_75t_R _10028_ (.A(_03232_),
    .Y(_03233_));
 NAND2x1_ASAP7_75t_R _10029_ (.A(_00032_),
    .B(_00033_),
    .Y(_03234_));
 AND2x2_ASAP7_75t_R _10030_ (.A(_03179_),
    .B(_03180_),
    .Y(_03235_));
 AND2x2_ASAP7_75t_R _10031_ (.A(_03182_),
    .B(_03183_),
    .Y(_03236_));
 AND4x1_ASAP7_75t_R _10032_ (.A(_03185_),
    .B(_03186_),
    .C(_03188_),
    .D(_03189_),
    .Y(_03237_));
 AND4x2_ASAP7_75t_R _10033_ (.A(_03234_),
    .B(_03235_),
    .C(_03236_),
    .D(_03237_),
    .Y(_03238_));
 AND2x2_ASAP7_75t_R _10034_ (.A(net1),
    .B(net11),
    .Y(_03239_));
 AND3x2_ASAP7_75t_R _10035_ (.A(_03016_),
    .B(net21),
    .C(_03239_),
    .Y(_03240_));
 NAND2x2_ASAP7_75t_R _10036_ (.A(_03017_),
    .B(net24),
    .Y(_03241_));
 OA21x2_ASAP7_75t_R _10037_ (.A1(_03238_),
    .A2(_03240_),
    .B(_03241_),
    .Y(_03242_));
 BUFx6f_ASAP7_75t_R _10038_ (.A(_03242_),
    .Y(_03243_));
 NAND2x2_ASAP7_75t_R _10039_ (.A(_03233_),
    .B(_03243_),
    .Y(_03244_));
 BUFx10_ASAP7_75t_R _10040_ (.A(_03244_),
    .Y(_03245_));
 BUFx6f_ASAP7_75t_R _10041_ (.A(_03245_),
    .Y(_03246_));
 BUFx6f_ASAP7_75t_R _10042_ (.A(_03246_),
    .Y(_03247_));
 AO21x1_ASAP7_75t_R _10043_ (.A1(_03177_),
    .A2(_03192_),
    .B(_03198_),
    .Y(_03248_));
 BUFx4f_ASAP7_75t_R _10044_ (.A(_03248_),
    .Y(_03249_));
 BUFx10_ASAP7_75t_R _10045_ (.A(_03207_),
    .Y(_03250_));
 BUFx16f_ASAP7_75t_R _10046_ (.A(_03250_),
    .Y(_03251_));
 INVx1_ASAP7_75t_R _10047_ (.A(net27),
    .Y(_03252_));
 OR4x2_ASAP7_75t_R _10048_ (.A(_03095_),
    .B(_03252_),
    .C(net25),
    .D(_03195_),
    .Y(_03253_));
 AND2x4_ASAP7_75t_R _10049_ (.A(_03251_),
    .B(_03253_),
    .Y(_03254_));
 OR2x2_ASAP7_75t_R _10050_ (.A(_03249_),
    .B(_03254_),
    .Y(_03255_));
 BUFx4f_ASAP7_75t_R _10051_ (.A(_03255_),
    .Y(_03256_));
 NAND2x2_ASAP7_75t_R _10052_ (.A(_03247_),
    .B(_03256_),
    .Y(_03257_));
 OR5x2_ASAP7_75t_R _10053_ (.A(_03099_),
    .B(net6),
    .C(_03220_),
    .D(_03230_),
    .E(_03257_),
    .Y(_03258_));
 BUFx12f_ASAP7_75t_R _10054_ (.A(_03258_),
    .Y(_03259_));
 BUFx10_ASAP7_75t_R _10055_ (.A(_03206_),
    .Y(_03260_));
 BUFx12f_ASAP7_75t_R _10056_ (.A(_03260_),
    .Y(_03261_));
 AND3x1_ASAP7_75t_R _10057_ (.A(_03261_),
    .B(_03221_),
    .C(_03227_),
    .Y(_03262_));
 INVx1_ASAP7_75t_R _10058_ (.A(net21),
    .Y(_03263_));
 OR3x2_ASAP7_75t_R _10059_ (.A(net170),
    .B(_03263_),
    .C(_03177_),
    .Y(_03264_));
 OR3x2_ASAP7_75t_R _10060_ (.A(_03264_),
    .B(_03241_),
    .C(_03253_),
    .Y(_03265_));
 AO21x1_ASAP7_75t_R _10061_ (.A1(_03231_),
    .A2(_03253_),
    .B(_03264_),
    .Y(_03266_));
 AND2x2_ASAP7_75t_R _10062_ (.A(_03016_),
    .B(net24),
    .Y(_03267_));
 AO21x1_ASAP7_75t_R _10063_ (.A1(_03192_),
    .A2(_03266_),
    .B(_03267_),
    .Y(_03268_));
 AND2x2_ASAP7_75t_R _10064_ (.A(_03265_),
    .B(_03268_),
    .Y(_03269_));
 OAI21x1_ASAP7_75t_R _10065_ (.A1(_03249_),
    .A2(_03262_),
    .B(_03269_),
    .Y(_03270_));
 AND2x6_ASAP7_75t_R _10066_ (.A(_03193_),
    .B(_03231_),
    .Y(_03271_));
 BUFx6f_ASAP7_75t_R _10067_ (.A(_03271_),
    .Y(_03272_));
 BUFx6f_ASAP7_75t_R _10068_ (.A(_03272_),
    .Y(_03273_));
 AND2x2_ASAP7_75t_R _10069_ (.A(_03267_),
    .B(_03253_),
    .Y(_03274_));
 AO221x2_ASAP7_75t_R _10070_ (.A1(_03192_),
    .A2(_03264_),
    .B1(_03273_),
    .B2(_03241_),
    .C(_03274_),
    .Y(_03275_));
 AND5x2_ASAP7_75t_R _10071_ (.A(_00032_),
    .B(_03203_),
    .C(_03235_),
    .D(_03236_),
    .E(_03237_),
    .Y(_03276_));
 BUFx12f_ASAP7_75t_R _10072_ (.A(_03276_),
    .Y(_03277_));
 BUFx12_ASAP7_75t_R _10073_ (.A(_03277_),
    .Y(_03278_));
 AO21x2_ASAP7_75t_R _10074_ (.A1(_03216_),
    .A2(net28),
    .B(_03278_),
    .Y(_03279_));
 OA22x2_ASAP7_75t_R _10075_ (.A1(_03249_),
    .A2(_03254_),
    .B1(_03279_),
    .B2(_03229_),
    .Y(_03280_));
 NAND2x2_ASAP7_75t_R _10076_ (.A(_03275_),
    .B(_03280_),
    .Y(_03281_));
 OA211x2_ASAP7_75t_R _10077_ (.A1(_03249_),
    .A2(_03262_),
    .B(_03268_),
    .C(_03265_),
    .Y(_03282_));
 BUFx4f_ASAP7_75t_R _10078_ (.A(_03282_),
    .Y(_03283_));
 BUFx4f_ASAP7_75t_R _10079_ (.A(_03273_),
    .Y(_03284_));
 AO21x2_ASAP7_75t_R _10080_ (.A1(_03192_),
    .A2(_03264_),
    .B(_03267_),
    .Y(_03285_));
 BUFx6f_ASAP7_75t_R _10081_ (.A(_03285_),
    .Y(_03286_));
 BUFx6f_ASAP7_75t_R _10082_ (.A(_03286_),
    .Y(_03287_));
 BUFx4f_ASAP7_75t_R _10083_ (.A(_03287_),
    .Y(_03288_));
 BUFx10_ASAP7_75t_R _10084_ (.A(_03122_),
    .Y(_03289_));
 BUFx10_ASAP7_75t_R _10085_ (.A(_03289_),
    .Y(_03290_));
 BUFx6f_ASAP7_75t_R _10086_ (.A(_03290_),
    .Y(_03291_));
 OA211x2_ASAP7_75t_R _10087_ (.A1(_03284_),
    .A2(_03288_),
    .B(_03291_),
    .C(_03229_),
    .Y(_03292_));
 OR2x2_ASAP7_75t_R _10088_ (.A(_03283_),
    .B(_03292_),
    .Y(_03293_));
 OAI22x1_ASAP7_75t_R _10089_ (.A1(_03176_),
    .A2(_03270_),
    .B1(_03281_),
    .B2(_03293_),
    .Y(_03294_));
 BUFx4f_ASAP7_75t_R _10090_ (.A(_03294_),
    .Y(_03295_));
 BUFx4f_ASAP7_75t_R _10091_ (.A(_03295_),
    .Y(_03296_));
 BUFx6f_ASAP7_75t_R _10092_ (.A(_03296_),
    .Y(_03297_));
 XNOR2x1_ASAP7_75t_R _10093_ (.B(_03297_),
    .Y(_09556_),
    .A(_03259_));
 INVx1_ASAP7_75t_R _10094_ (.A(_09556_),
    .Y(_09558_));
 NAND2x2_ASAP7_75t_R _10095_ (.A(_03018_),
    .B(net9),
    .Y(_03298_));
 BUFx10_ASAP7_75t_R _10096_ (.A(_03298_),
    .Y(_03299_));
 BUFx10_ASAP7_75t_R _10097_ (.A(_03299_),
    .Y(_03300_));
 BUFx12f_ASAP7_75t_R _10098_ (.A(instr[15]),
    .Y(_03301_));
 AND2x4_ASAP7_75t_R _10099_ (.A(_03016_),
    .B(_03301_),
    .Y(_03302_));
 BUFx10_ASAP7_75t_R _10100_ (.A(_03302_),
    .Y(_03303_));
 BUFx6f_ASAP7_75t_R _10101_ (.A(_03303_),
    .Y(_03304_));
 BUFx12_ASAP7_75t_R _10102_ (.A(_03304_),
    .Y(_03305_));
 BUFx16f_ASAP7_75t_R _10103_ (.A(_03305_),
    .Y(_03306_));
 NOR2x1_ASAP7_75t_R _10104_ (.A(_00002_),
    .B(_03306_),
    .Y(_03307_));
 OR5x2_ASAP7_75t_R _10105_ (.A(net169),
    .B(_03263_),
    .C(net27),
    .D(_03194_),
    .E(_03177_),
    .Y(_03308_));
 BUFx6f_ASAP7_75t_R _10106_ (.A(_03308_),
    .Y(_03309_));
 BUFx6f_ASAP7_75t_R _10107_ (.A(_03309_),
    .Y(_03310_));
 BUFx12_ASAP7_75t_R _10108_ (.A(_03310_),
    .Y(_03311_));
 BUFx10_ASAP7_75t_R _10109_ (.A(_03303_),
    .Y(_03312_));
 BUFx12f_ASAP7_75t_R _10110_ (.A(_03312_),
    .Y(_03313_));
 INVx1_ASAP7_75t_R _10111_ (.A(_00003_),
    .Y(_03314_));
 OA211x2_ASAP7_75t_R _10112_ (.A1(_03226_),
    .A2(_03311_),
    .B(_03313_),
    .C(_03314_),
    .Y(_03315_));
 BUFx10_ASAP7_75t_R _10113_ (.A(_03207_),
    .Y(_03316_));
 BUFx6f_ASAP7_75t_R _10114_ (.A(_03316_),
    .Y(_03317_));
 NAND2x2_ASAP7_75t_R _10115_ (.A(_03016_),
    .B(net8),
    .Y(_03318_));
 BUFx6f_ASAP7_75t_R _10116_ (.A(_03318_),
    .Y(_03319_));
 BUFx6f_ASAP7_75t_R _10117_ (.A(_03319_),
    .Y(_03320_));
 BUFx10_ASAP7_75t_R _10118_ (.A(_03320_),
    .Y(_03321_));
 BUFx6f_ASAP7_75t_R _10119_ (.A(_03321_),
    .Y(_03322_));
 OA211x2_ASAP7_75t_R _10120_ (.A1(_03307_),
    .A2(_03315_),
    .B(_03317_),
    .C(_03322_),
    .Y(_03323_));
 BUFx6f_ASAP7_75t_R _10121_ (.A(_03206_),
    .Y(_03324_));
 BUFx10_ASAP7_75t_R _10122_ (.A(_03324_),
    .Y(_03325_));
 BUFx10_ASAP7_75t_R _10123_ (.A(_03325_),
    .Y(_03326_));
 BUFx10_ASAP7_75t_R _10124_ (.A(_03303_),
    .Y(_03327_));
 BUFx12_ASAP7_75t_R _10125_ (.A(_03327_),
    .Y(_03328_));
 BUFx10_ASAP7_75t_R _10126_ (.A(_03328_),
    .Y(_03329_));
 BUFx12f_ASAP7_75t_R _10127_ (.A(_03329_),
    .Y(_03330_));
 NAND2x1_ASAP7_75t_R _10128_ (.A(_03016_),
    .B(_03301_),
    .Y(_03331_));
 BUFx6f_ASAP7_75t_R _10129_ (.A(_03331_),
    .Y(_03332_));
 BUFx12_ASAP7_75t_R _10130_ (.A(_03332_),
    .Y(_03333_));
 BUFx16f_ASAP7_75t_R _10131_ (.A(_03333_),
    .Y(_03334_));
 BUFx16f_ASAP7_75t_R _10132_ (.A(_03334_),
    .Y(_03335_));
 AND2x2_ASAP7_75t_R _10133_ (.A(_00006_),
    .B(_03335_),
    .Y(_03336_));
 AOI221x1_ASAP7_75t_R _10134_ (.A1(_03326_),
    .A2(_03322_),
    .B1(_03330_),
    .B2(_00007_),
    .C(_03336_),
    .Y(_03337_));
 NAND2x2_ASAP7_75t_R _10135_ (.A(_03016_),
    .B(net7),
    .Y(_03338_));
 NAND2x2_ASAP7_75t_R _10136_ (.A(_03206_),
    .B(_03338_),
    .Y(_03339_));
 BUFx12_ASAP7_75t_R _10137_ (.A(_03339_),
    .Y(_03340_));
 BUFx10_ASAP7_75t_R _10138_ (.A(_03340_),
    .Y(_03341_));
 OAI21x1_ASAP7_75t_R _10139_ (.A1(_03323_),
    .A2(_03337_),
    .B(_03341_),
    .Y(_03342_));
 AND2x2_ASAP7_75t_R _10140_ (.A(_03233_),
    .B(_03243_),
    .Y(_03343_));
 BUFx6f_ASAP7_75t_R _10141_ (.A(_03343_),
    .Y(_03344_));
 BUFx6f_ASAP7_75t_R _10142_ (.A(_03344_),
    .Y(_03345_));
 AO21x1_ASAP7_75t_R _10143_ (.A1(_03300_),
    .A2(_03342_),
    .B(_03345_),
    .Y(_03346_));
 BUFx10_ASAP7_75t_R _10144_ (.A(_03302_),
    .Y(_03347_));
 BUFx16f_ASAP7_75t_R _10145_ (.A(_03347_),
    .Y(_03348_));
 BUFx16f_ASAP7_75t_R _10146_ (.A(_03348_),
    .Y(_03349_));
 BUFx12f_ASAP7_75t_R _10147_ (.A(_03349_),
    .Y(_03350_));
 CKINVDCx11_ASAP7_75t_R _10148_ (.A(net24),
    .Y(_03351_));
 AND5x2_ASAP7_75t_R _10149_ (.A(_03016_),
    .B(net21),
    .C(_03252_),
    .D(net25),
    .E(_03239_),
    .Y(_03352_));
 AO21x1_ASAP7_75t_R _10150_ (.A1(_03351_),
    .A2(_03352_),
    .B(_03331_),
    .Y(_03353_));
 BUFx12_ASAP7_75t_R _10151_ (.A(_03353_),
    .Y(_03354_));
 BUFx16f_ASAP7_75t_R _10152_ (.A(_03354_),
    .Y(_03355_));
 BUFx16f_ASAP7_75t_R _10153_ (.A(_03355_),
    .Y(_03356_));
 BUFx16f_ASAP7_75t_R _10154_ (.A(_03356_),
    .Y(_03357_));
 OAI22x1_ASAP7_75t_R _10155_ (.A1(_00004_),
    .A2(_03350_),
    .B1(_03357_),
    .B2(_00005_),
    .Y(_03358_));
 AND2x6_ASAP7_75t_R _10156_ (.A(_03017_),
    .B(net8),
    .Y(_03359_));
 AND2x4_ASAP7_75t_R _10157_ (.A(_03338_),
    .B(_03359_),
    .Y(_03360_));
 BUFx6f_ASAP7_75t_R _10158_ (.A(_03360_),
    .Y(_03361_));
 BUFx10_ASAP7_75t_R _10159_ (.A(_03361_),
    .Y(_03362_));
 NAND2x1_ASAP7_75t_R _10160_ (.A(_03358_),
    .B(_03362_),
    .Y(_03363_));
 BUFx6f_ASAP7_75t_R _10161_ (.A(_03197_),
    .Y(_03364_));
 BUFx6f_ASAP7_75t_R _10162_ (.A(_03309_),
    .Y(_03365_));
 OA211x2_ASAP7_75t_R _10163_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03348_),
    .C(_00001_),
    .Y(_03366_));
 AO21x1_ASAP7_75t_R _10164_ (.A1(_00000_),
    .A2(_03356_),
    .B(_03366_),
    .Y(_03367_));
 INVx1_ASAP7_75t_R _10165_ (.A(_03188_),
    .Y(_03368_));
 INVx1_ASAP7_75t_R _10166_ (.A(_00032_),
    .Y(_03369_));
 OR4x1_ASAP7_75t_R _10167_ (.A(_03369_),
    .B(_00033_),
    .C(net65),
    .D(net95),
    .Y(_03370_));
 OR5x2_ASAP7_75t_R _10168_ (.A(_03181_),
    .B(_03184_),
    .C(_03187_),
    .D(_03368_),
    .E(_03370_),
    .Y(_03371_));
 AND2x2_ASAP7_75t_R _10169_ (.A(_03338_),
    .B(_03318_),
    .Y(_03372_));
 NAND2x2_ASAP7_75t_R _10170_ (.A(_03371_),
    .B(_03372_),
    .Y(_03373_));
 OR2x2_ASAP7_75t_R _10171_ (.A(_03367_),
    .B(_03373_),
    .Y(_03374_));
 OR3x1_ASAP7_75t_R _10172_ (.A(_03273_),
    .B(_03287_),
    .C(_03367_),
    .Y(_03375_));
 OA211x2_ASAP7_75t_R _10173_ (.A1(_03344_),
    .A2(_03363_),
    .B(_03374_),
    .C(_03375_),
    .Y(_03376_));
 BUFx12_ASAP7_75t_R _10174_ (.A(_03335_),
    .Y(_03377_));
 BUFx16f_ASAP7_75t_R _10175_ (.A(_03335_),
    .Y(_03378_));
 NAND2x1_ASAP7_75t_R _10176_ (.A(_00014_),
    .B(_03378_),
    .Y(_03379_));
 OA21x2_ASAP7_75t_R _10177_ (.A1(_03150_),
    .A2(_03377_),
    .B(_03379_),
    .Y(_03380_));
 AND2x6_ASAP7_75t_R _10178_ (.A(_03017_),
    .B(net7),
    .Y(_03381_));
 BUFx10_ASAP7_75t_R _10179_ (.A(_03381_),
    .Y(_03382_));
 BUFx10_ASAP7_75t_R _10180_ (.A(_03356_),
    .Y(_03383_));
 BUFx12f_ASAP7_75t_R _10181_ (.A(_03327_),
    .Y(_03384_));
 BUFx12f_ASAP7_75t_R _10182_ (.A(_03384_),
    .Y(_03385_));
 BUFx6f_ASAP7_75t_R _10183_ (.A(_03319_),
    .Y(_03386_));
 BUFx10_ASAP7_75t_R _10184_ (.A(_03386_),
    .Y(_03387_));
 BUFx12f_ASAP7_75t_R _10185_ (.A(_03387_),
    .Y(_03388_));
 OA21x2_ASAP7_75t_R _10186_ (.A1(_00010_),
    .A2(_03385_),
    .B(_03388_),
    .Y(_03389_));
 OAI21x1_ASAP7_75t_R _10187_ (.A1(_00011_),
    .A2(_03383_),
    .B(_03389_),
    .Y(_03390_));
 AO21x1_ASAP7_75t_R _10188_ (.A1(_03382_),
    .A2(_03390_),
    .B(_03278_),
    .Y(_03391_));
 AND2x2_ASAP7_75t_R _10189_ (.A(_03205_),
    .B(_03319_),
    .Y(_03392_));
 BUFx12_ASAP7_75t_R _10190_ (.A(_03392_),
    .Y(_03393_));
 BUFx6f_ASAP7_75t_R _10191_ (.A(_03393_),
    .Y(_03394_));
 BUFx12f_ASAP7_75t_R _10192_ (.A(_03333_),
    .Y(_03395_));
 BUFx12_ASAP7_75t_R _10193_ (.A(_03395_),
    .Y(_03396_));
 BUFx12f_ASAP7_75t_R _10194_ (.A(_03396_),
    .Y(_03397_));
 OA21x2_ASAP7_75t_R _10195_ (.A1(net24),
    .A2(_03308_),
    .B(_03302_),
    .Y(_03398_));
 BUFx6f_ASAP7_75t_R _10196_ (.A(_03398_),
    .Y(_03399_));
 BUFx12_ASAP7_75t_R _10197_ (.A(_03399_),
    .Y(_03400_));
 BUFx16f_ASAP7_75t_R _10198_ (.A(_03400_),
    .Y(_03401_));
 OAI22x1_ASAP7_75t_R _10199_ (.A1(_00013_),
    .A2(_03397_),
    .B1(_03401_),
    .B2(_00012_),
    .Y(_03402_));
 AO32x1_ASAP7_75t_R _10200_ (.A1(_03382_),
    .A2(_03394_),
    .A3(_03390_),
    .B1(_03402_),
    .B2(_03362_),
    .Y(_03403_));
 AO21x2_ASAP7_75t_R _10201_ (.A1(_03233_),
    .A2(_03243_),
    .B(_03298_),
    .Y(_03404_));
 BUFx10_ASAP7_75t_R _10202_ (.A(_03404_),
    .Y(_03405_));
 BUFx10_ASAP7_75t_R _10203_ (.A(_03405_),
    .Y(_03406_));
 AOI211x1_ASAP7_75t_R _10204_ (.A1(_03380_),
    .A2(_03391_),
    .B(_03403_),
    .C(_03406_),
    .Y(_03407_));
 BUFx16f_ASAP7_75t_R _10205_ (.A(_03399_),
    .Y(_03408_));
 BUFx12_ASAP7_75t_R _10206_ (.A(_03408_),
    .Y(_03409_));
 BUFx10_ASAP7_75t_R _10207_ (.A(_03409_),
    .Y(_03410_));
 BUFx6f_ASAP7_75t_R _10208_ (.A(_03373_),
    .Y(_03411_));
 BUFx12_ASAP7_75t_R _10209_ (.A(_03245_),
    .Y(_03412_));
 BUFx12f_ASAP7_75t_R _10210_ (.A(_03354_),
    .Y(_03413_));
 BUFx16f_ASAP7_75t_R _10211_ (.A(_03413_),
    .Y(_03414_));
 BUFx10_ASAP7_75t_R _10212_ (.A(_03414_),
    .Y(_03415_));
 AND2x2_ASAP7_75t_R _10213_ (.A(_00008_),
    .B(_03415_),
    .Y(_03416_));
 AO221x1_ASAP7_75t_R _10214_ (.A1(_00009_),
    .A2(_03410_),
    .B1(_03411_),
    .B2(_03412_),
    .C(_03416_),
    .Y(_03417_));
 BUFx16f_ASAP7_75t_R _10215_ (.A(_03355_),
    .Y(_03418_));
 AND2x2_ASAP7_75t_R _10216_ (.A(_03371_),
    .B(_03372_),
    .Y(_03419_));
 BUFx12f_ASAP7_75t_R _10217_ (.A(_03419_),
    .Y(_03420_));
 AO22x2_ASAP7_75t_R _10218_ (.A1(_03233_),
    .A2(_03243_),
    .B1(_03298_),
    .B2(_03420_),
    .Y(_03421_));
 AND2x6_ASAP7_75t_R _10219_ (.A(_03017_),
    .B(net10),
    .Y(_03422_));
 OA21x2_ASAP7_75t_R _10220_ (.A1(_03271_),
    .A2(_03285_),
    .B(_03422_),
    .Y(_03423_));
 BUFx6f_ASAP7_75t_R _10221_ (.A(_03423_),
    .Y(_03424_));
 AO21x2_ASAP7_75t_R _10222_ (.A1(_03418_),
    .A2(_03421_),
    .B(_03424_),
    .Y(_03425_));
 BUFx12_ASAP7_75t_R _10223_ (.A(_03425_),
    .Y(_03426_));
 AOI221x1_ASAP7_75t_R _10224_ (.A1(_03346_),
    .A2(_03376_),
    .B1(_03407_),
    .B2(_03417_),
    .C(_03426_),
    .Y(_03427_));
 BUFx12f_ASAP7_75t_R _10225_ (.A(_03348_),
    .Y(_03428_));
 BUFx12f_ASAP7_75t_R _10226_ (.A(_03428_),
    .Y(_03429_));
 BUFx12f_ASAP7_75t_R _10227_ (.A(_03354_),
    .Y(_03430_));
 BUFx12f_ASAP7_75t_R _10228_ (.A(_03430_),
    .Y(_03431_));
 BUFx12f_ASAP7_75t_R _10229_ (.A(_03431_),
    .Y(_03432_));
 OAI22x1_ASAP7_75t_R _10230_ (.A1(_00018_),
    .A2(_03429_),
    .B1(_03432_),
    .B2(_00019_),
    .Y(_03433_));
 AND2x2_ASAP7_75t_R _10231_ (.A(_03394_),
    .B(_03433_),
    .Y(_03434_));
 BUFx10_ASAP7_75t_R _10232_ (.A(_03332_),
    .Y(_03435_));
 BUFx12f_ASAP7_75t_R _10233_ (.A(_03435_),
    .Y(_03436_));
 BUFx12f_ASAP7_75t_R _10234_ (.A(_03436_),
    .Y(_03437_));
 NAND2x1_ASAP7_75t_R _10235_ (.A(_00022_),
    .B(_03437_),
    .Y(_03438_));
 NAND2x2_ASAP7_75t_R _10236_ (.A(_03206_),
    .B(_03319_),
    .Y(_03439_));
 BUFx12f_ASAP7_75t_R _10237_ (.A(_03439_),
    .Y(_03440_));
 BUFx12_ASAP7_75t_R _10238_ (.A(_03440_),
    .Y(_03441_));
 OA211x2_ASAP7_75t_R _10239_ (.A1(_03030_),
    .A2(_03397_),
    .B(_03438_),
    .C(_03441_),
    .Y(_03442_));
 OA21x2_ASAP7_75t_R _10240_ (.A1(_03272_),
    .A2(_03286_),
    .B(_03339_),
    .Y(_03443_));
 BUFx6f_ASAP7_75t_R _10241_ (.A(_03443_),
    .Y(_03444_));
 OA21x2_ASAP7_75t_R _10242_ (.A1(_03434_),
    .A2(_03442_),
    .B(_03444_),
    .Y(_03445_));
 AO21x2_ASAP7_75t_R _10243_ (.A1(_03232_),
    .A2(_03242_),
    .B(_03419_),
    .Y(_03446_));
 BUFx10_ASAP7_75t_R _10244_ (.A(_03446_),
    .Y(_03447_));
 BUFx10_ASAP7_75t_R _10245_ (.A(_03447_),
    .Y(_03448_));
 BUFx12_ASAP7_75t_R _10246_ (.A(_03354_),
    .Y(_03449_));
 BUFx12f_ASAP7_75t_R _10247_ (.A(_03449_),
    .Y(_03450_));
 BUFx12_ASAP7_75t_R _10248_ (.A(_03450_),
    .Y(_03451_));
 NAND2x1_ASAP7_75t_R _10249_ (.A(_00016_),
    .B(_03451_),
    .Y(_03452_));
 BUFx16f_ASAP7_75t_R _10250_ (.A(_03398_),
    .Y(_03453_));
 BUFx12f_ASAP7_75t_R _10251_ (.A(_03453_),
    .Y(_03454_));
 BUFx12f_ASAP7_75t_R _10252_ (.A(_03454_),
    .Y(_03455_));
 NAND2x1_ASAP7_75t_R _10253_ (.A(_00017_),
    .B(_03455_),
    .Y(_03456_));
 BUFx10_ASAP7_75t_R _10254_ (.A(_03361_),
    .Y(_03457_));
 OAI22x1_ASAP7_75t_R _10255_ (.A1(_00020_),
    .A2(_03429_),
    .B1(_03432_),
    .B2(_00021_),
    .Y(_03458_));
 AND2x4_ASAP7_75t_R _10256_ (.A(_03017_),
    .B(net9),
    .Y(_03459_));
 BUFx4f_ASAP7_75t_R _10257_ (.A(_03459_),
    .Y(_03460_));
 BUFx6f_ASAP7_75t_R _10258_ (.A(_03460_),
    .Y(_03461_));
 AO21x1_ASAP7_75t_R _10259_ (.A1(_03457_),
    .A2(_03458_),
    .B(_03461_),
    .Y(_03462_));
 AO32x1_ASAP7_75t_R _10260_ (.A1(_03448_),
    .A2(_03452_),
    .A3(_03456_),
    .B1(_03462_),
    .B2(_03412_),
    .Y(_03463_));
 INVx1_ASAP7_75t_R _10261_ (.A(_00026_),
    .Y(_03464_));
 BUFx10_ASAP7_75t_R _10262_ (.A(_03332_),
    .Y(_03465_));
 BUFx10_ASAP7_75t_R _10263_ (.A(_03465_),
    .Y(_03466_));
 BUFx16f_ASAP7_75t_R _10264_ (.A(_03399_),
    .Y(_03467_));
 BUFx10_ASAP7_75t_R _10265_ (.A(_03359_),
    .Y(_03468_));
 AO221x1_ASAP7_75t_R _10266_ (.A1(_03464_),
    .A2(_03466_),
    .B1(_03467_),
    .B2(_03164_),
    .C(_03468_),
    .Y(_03469_));
 BUFx6f_ASAP7_75t_R _10267_ (.A(_03277_),
    .Y(_03470_));
 AO21x1_ASAP7_75t_R _10268_ (.A1(_03382_),
    .A2(_03469_),
    .B(_03470_),
    .Y(_03471_));
 BUFx12f_ASAP7_75t_R _10269_ (.A(_03440_),
    .Y(_03472_));
 BUFx12f_ASAP7_75t_R _10270_ (.A(_03019_),
    .Y(_03473_));
 BUFx6f_ASAP7_75t_R _10271_ (.A(_03301_),
    .Y(_03474_));
 BUFx12f_ASAP7_75t_R _10272_ (.A(_03474_),
    .Y(_03475_));
 AND3x1_ASAP7_75t_R _10273_ (.A(_00031_),
    .B(_03473_),
    .C(_03475_),
    .Y(_03476_));
 AO21x1_ASAP7_75t_R _10274_ (.A1(_00030_),
    .A2(_03437_),
    .B(_03476_),
    .Y(_03477_));
 NAND2x1_ASAP7_75t_R _10275_ (.A(_03472_),
    .B(_03477_),
    .Y(_03478_));
 BUFx12f_ASAP7_75t_R _10276_ (.A(_03454_),
    .Y(_03479_));
 OAI22x1_ASAP7_75t_R _10277_ (.A1(_00029_),
    .A2(_03378_),
    .B1(_03479_),
    .B2(_00028_),
    .Y(_03480_));
 OA21x2_ASAP7_75t_R _10278_ (.A1(_03271_),
    .A2(_03286_),
    .B(_03360_),
    .Y(_03481_));
 BUFx6f_ASAP7_75t_R _10279_ (.A(_03481_),
    .Y(_03482_));
 BUFx6f_ASAP7_75t_R _10280_ (.A(_03482_),
    .Y(_03483_));
 BUFx12f_ASAP7_75t_R _10281_ (.A(_03420_),
    .Y(_03484_));
 BUFx16f_ASAP7_75t_R _10282_ (.A(_03354_),
    .Y(_03485_));
 BUFx12f_ASAP7_75t_R _10283_ (.A(_03485_),
    .Y(_03486_));
 BUFx6f_ASAP7_75t_R _10284_ (.A(_03197_),
    .Y(_03487_));
 BUFx6f_ASAP7_75t_R _10285_ (.A(_03487_),
    .Y(_03488_));
 BUFx6f_ASAP7_75t_R _10286_ (.A(_03309_),
    .Y(_03489_));
 BUFx10_ASAP7_75t_R _10287_ (.A(_03489_),
    .Y(_03490_));
 OA211x2_ASAP7_75t_R _10288_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03384_),
    .C(_03165_),
    .Y(_03491_));
 AO21x1_ASAP7_75t_R _10289_ (.A1(_03168_),
    .A2(_03486_),
    .B(_03491_),
    .Y(_03492_));
 AO21x1_ASAP7_75t_R _10290_ (.A1(_03484_),
    .A2(_03492_),
    .B(_03299_),
    .Y(_03493_));
 AO221x1_ASAP7_75t_R _10291_ (.A1(_03471_),
    .A2(_03478_),
    .B1(_03480_),
    .B2(_03483_),
    .C(_03493_),
    .Y(_03494_));
 BUFx10_ASAP7_75t_R _10292_ (.A(_03424_),
    .Y(_03495_));
 OA211x2_ASAP7_75t_R _10293_ (.A1(_03445_),
    .A2(_03463_),
    .B(_03494_),
    .C(_03495_),
    .Y(_03496_));
 OR2x2_ASAP7_75t_R _10294_ (.A(_03427_),
    .B(_03496_),
    .Y(_03497_));
 BUFx2_ASAP7_75t_R _10295_ (.A(_03497_),
    .Y(_09555_));
 INVx1_ASAP7_75t_R _10296_ (.A(_09555_),
    .Y(_09557_));
 AOI21x1_ASAP7_75t_R _10297_ (.A1(_03431_),
    .A2(_03421_),
    .B(_03424_),
    .Y(_03498_));
 BUFx10_ASAP7_75t_R _10298_ (.A(_03498_),
    .Y(_03499_));
 OAI22x1_ASAP7_75t_R _10299_ (.A1(_00048_),
    .A2(_03378_),
    .B1(_03479_),
    .B2(_00047_),
    .Y(_03500_));
 BUFx12f_ASAP7_75t_R _10300_ (.A(_03339_),
    .Y(_03501_));
 BUFx10_ASAP7_75t_R _10301_ (.A(_03501_),
    .Y(_03502_));
 BUFx10_ASAP7_75t_R _10302_ (.A(_03439_),
    .Y(_03503_));
 BUFx12f_ASAP7_75t_R _10303_ (.A(_03503_),
    .Y(_03504_));
 OA22x2_ASAP7_75t_R _10304_ (.A1(_00045_),
    .A2(_03384_),
    .B1(_03449_),
    .B2(_00046_),
    .Y(_03505_));
 BUFx12_ASAP7_75t_R _10305_ (.A(_03386_),
    .Y(_03506_));
 BUFx12f_ASAP7_75t_R _10306_ (.A(_03347_),
    .Y(_03507_));
 AND2x2_ASAP7_75t_R _10307_ (.A(_00049_),
    .B(_03333_),
    .Y(_03508_));
 AO221x1_ASAP7_75t_R _10308_ (.A1(_03324_),
    .A2(_03506_),
    .B1(_03507_),
    .B2(_00050_),
    .C(_03508_),
    .Y(_03509_));
 OAI21x1_ASAP7_75t_R _10309_ (.A1(_03504_),
    .A2(_03505_),
    .B(_03509_),
    .Y(_03510_));
 BUFx12f_ASAP7_75t_R _10310_ (.A(_03453_),
    .Y(_03511_));
 OR2x2_ASAP7_75t_R _10311_ (.A(_00044_),
    .B(_03413_),
    .Y(_03512_));
 OAI21x1_ASAP7_75t_R _10312_ (.A1(_00043_),
    .A2(_03511_),
    .B(_03512_),
    .Y(_03513_));
 AO221x1_ASAP7_75t_R _10313_ (.A1(_03502_),
    .A2(_03510_),
    .B1(_03513_),
    .B2(_03447_),
    .C(_03405_),
    .Y(_03514_));
 AO21x1_ASAP7_75t_R _10314_ (.A1(_03483_),
    .A2(_03500_),
    .B(_03514_),
    .Y(_03515_));
 BUFx6f_ASAP7_75t_R _10315_ (.A(_03482_),
    .Y(_03516_));
 OAI22x1_ASAP7_75t_R _10316_ (.A1(_00039_),
    .A2(_03429_),
    .B1(_03432_),
    .B2(_00040_),
    .Y(_03517_));
 INVx1_ASAP7_75t_R _10317_ (.A(_00035_),
    .Y(_01246_));
 NAND2x1_ASAP7_75t_R _10318_ (.A(_00036_),
    .B(_03400_),
    .Y(_03518_));
 OA21x2_ASAP7_75t_R _10319_ (.A1(_01246_),
    .A2(_03454_),
    .B(_03518_),
    .Y(_03519_));
 BUFx6f_ASAP7_75t_R _10320_ (.A(_03446_),
    .Y(_03520_));
 BUFx6f_ASAP7_75t_R _10321_ (.A(_03245_),
    .Y(_03521_));
 BUFx12f_ASAP7_75t_R _10322_ (.A(_03327_),
    .Y(_03522_));
 OA22x2_ASAP7_75t_R _10323_ (.A1(_00037_),
    .A2(_03522_),
    .B1(_03485_),
    .B2(_00038_),
    .Y(_03523_));
 AND2x2_ASAP7_75t_R _10324_ (.A(_00041_),
    .B(_03333_),
    .Y(_03524_));
 AO221x1_ASAP7_75t_R _10325_ (.A1(_03260_),
    .A2(_03506_),
    .B1(_03507_),
    .B2(_00042_),
    .C(_03524_),
    .Y(_03525_));
 OAI21x1_ASAP7_75t_R _10326_ (.A1(_03504_),
    .A2(_03523_),
    .B(_03525_),
    .Y(_03526_));
 AO21x1_ASAP7_75t_R _10327_ (.A1(_03502_),
    .A2(_03526_),
    .B(_03460_),
    .Y(_03527_));
 AO222x2_ASAP7_75t_R _10328_ (.A1(_03516_),
    .A2(_03517_),
    .B1(_03519_),
    .B2(_03520_),
    .C1(_03521_),
    .C2(_03527_),
    .Y(_03528_));
 BUFx16f_ASAP7_75t_R _10329_ (.A(_03431_),
    .Y(_03529_));
 OAI22x1_ASAP7_75t_R _10330_ (.A1(_00055_),
    .A2(_03429_),
    .B1(_03529_),
    .B2(_00056_),
    .Y(_03530_));
 OR2x2_ASAP7_75t_R _10331_ (.A(_00052_),
    .B(_03431_),
    .Y(_03531_));
 OAI21x1_ASAP7_75t_R _10332_ (.A1(_00051_),
    .A2(_03409_),
    .B(_03531_),
    .Y(_03532_));
 OA22x2_ASAP7_75t_R _10333_ (.A1(_00053_),
    .A2(_03522_),
    .B1(_03485_),
    .B2(_00054_),
    .Y(_03533_));
 AND3x1_ASAP7_75t_R _10334_ (.A(_03043_),
    .B(_03474_),
    .C(_00058_),
    .Y(_03534_));
 AO221x1_ASAP7_75t_R _10335_ (.A1(_03260_),
    .A2(_03506_),
    .B1(_03395_),
    .B2(_00057_),
    .C(_03534_),
    .Y(_03535_));
 OAI21x1_ASAP7_75t_R _10336_ (.A1(_03504_),
    .A2(_03533_),
    .B(_03535_),
    .Y(_03536_));
 AO21x1_ASAP7_75t_R _10337_ (.A1(_03502_),
    .A2(_03536_),
    .B(_03460_),
    .Y(_03537_));
 AO222x2_ASAP7_75t_R _10338_ (.A1(_03516_),
    .A2(_03530_),
    .B1(_03532_),
    .B2(_03520_),
    .C1(_03521_),
    .C2(_03537_),
    .Y(_03538_));
 BUFx10_ASAP7_75t_R _10339_ (.A(_03422_),
    .Y(_03539_));
 BUFx10_ASAP7_75t_R _10340_ (.A(_03482_),
    .Y(_03540_));
 BUFx12f_ASAP7_75t_R _10341_ (.A(_03408_),
    .Y(_03541_));
 OAI22x1_ASAP7_75t_R _10342_ (.A1(_00064_),
    .A2(_03397_),
    .B1(_03541_),
    .B2(_00063_),
    .Y(_03542_));
 NAND2x1_ASAP7_75t_R _10343_ (.A(_00066_),
    .B(_03328_),
    .Y(_03543_));
 NAND2x1_ASAP7_75t_R _10344_ (.A(_00065_),
    .B(_03395_),
    .Y(_03544_));
 OAI22x1_ASAP7_75t_R _10345_ (.A1(_00061_),
    .A2(_03507_),
    .B1(_03355_),
    .B2(_00062_),
    .Y(_03545_));
 AO32x1_ASAP7_75t_R _10346_ (.A1(_03359_),
    .A2(_03543_),
    .A3(_03544_),
    .B1(_03393_),
    .B2(_03545_),
    .Y(_03546_));
 INVx1_ASAP7_75t_R _10347_ (.A(_00060_),
    .Y(_03547_));
 NAND2x1_ASAP7_75t_R _10348_ (.A(_00059_),
    .B(_03355_),
    .Y(_03548_));
 OA211x2_ASAP7_75t_R _10349_ (.A1(_03547_),
    .A2(_03449_),
    .B(_03420_),
    .C(_03548_),
    .Y(_03549_));
 BUFx10_ASAP7_75t_R _10350_ (.A(_03298_),
    .Y(_03550_));
 AO211x2_ASAP7_75t_R _10351_ (.A1(_03382_),
    .A2(_03546_),
    .B(_03549_),
    .C(_03550_),
    .Y(_03551_));
 AO32x1_ASAP7_75t_R _10352_ (.A1(_03539_),
    .A2(_03540_),
    .A3(_03542_),
    .B1(_03551_),
    .B2(_03495_),
    .Y(_03552_));
 AO32x2_ASAP7_75t_R _10353_ (.A1(_03499_),
    .A2(_03515_),
    .A3(_03528_),
    .B1(_03538_),
    .B2(_03552_),
    .Y(_03553_));
 BUFx6f_ASAP7_75t_R _10354_ (.A(_03553_),
    .Y(_03554_));
 BUFx4f_ASAP7_75t_R _10355_ (.A(_03554_),
    .Y(_03555_));
 BUFx6f_ASAP7_75t_R _10356_ (.A(_03555_),
    .Y(_09561_));
 INVx1_ASAP7_75t_R _10357_ (.A(_09561_),
    .Y(_09563_));
 CKINVDCx10_ASAP7_75t_R _10358_ (.A(_03259_),
    .Y(_03556_));
 BUFx6f_ASAP7_75t_R _10359_ (.A(_03556_),
    .Y(_03557_));
 BUFx4f_ASAP7_75t_R _10360_ (.A(_03283_),
    .Y(_03558_));
 AND3x4_ASAP7_75t_R _10361_ (.A(_03037_),
    .B(_03026_),
    .C(_03017_),
    .Y(_03559_));
 BUFx10_ASAP7_75t_R _10362_ (.A(_03559_),
    .Y(_03560_));
 BUFx10_ASAP7_75t_R _10363_ (.A(_03560_),
    .Y(_03561_));
 AND2x2_ASAP7_75t_R _10364_ (.A(_03086_),
    .B(_00045_),
    .Y(_03562_));
 AO21x1_ASAP7_75t_R _10365_ (.A1(_03027_),
    .A2(_00043_),
    .B(_03562_),
    .Y(_03563_));
 BUFx6f_ASAP7_75t_R _10366_ (.A(_03053_),
    .Y(_03564_));
 BUFx6f_ASAP7_75t_R _10367_ (.A(_03564_),
    .Y(_03565_));
 BUFx10_ASAP7_75t_R _10368_ (.A(_03565_),
    .Y(_03566_));
 AND2x6_ASAP7_75t_R _10369_ (.A(_03038_),
    .B(_03085_),
    .Y(_03567_));
 BUFx6f_ASAP7_75t_R _10370_ (.A(_03567_),
    .Y(_03568_));
 AO21x1_ASAP7_75t_R _10371_ (.A1(_00046_),
    .A2(_03568_),
    .B(_03077_),
    .Y(_03569_));
 AO221x1_ASAP7_75t_R _10372_ (.A1(_00044_),
    .A2(_03561_),
    .B1(_03563_),
    .B2(_03566_),
    .C(_03569_),
    .Y(_03570_));
 BUFx10_ASAP7_75t_R _10373_ (.A(_03088_),
    .Y(_03571_));
 BUFx12f_ASAP7_75t_R _10374_ (.A(_03053_),
    .Y(_03572_));
 BUFx12f_ASAP7_75t_R _10375_ (.A(_03572_),
    .Y(_03573_));
 AND2x2_ASAP7_75t_R _10376_ (.A(_03091_),
    .B(_00050_),
    .Y(_03574_));
 AO21x1_ASAP7_75t_R _10377_ (.A1(_03573_),
    .A2(_00049_),
    .B(_03574_),
    .Y(_03575_));
 BUFx6f_ASAP7_75t_R _10378_ (.A(_03122_),
    .Y(_03576_));
 BUFx10_ASAP7_75t_R _10379_ (.A(_03576_),
    .Y(_03577_));
 BUFx12_ASAP7_75t_R _10380_ (.A(_03090_),
    .Y(_03578_));
 AND3x1_ASAP7_75t_R _10381_ (.A(_03578_),
    .B(_03063_),
    .C(_00048_),
    .Y(_03579_));
 AO21x1_ASAP7_75t_R _10382_ (.A1(_00047_),
    .A2(_03577_),
    .B(_03579_),
    .Y(_03580_));
 BUFx6f_ASAP7_75t_R _10383_ (.A(_03121_),
    .Y(_03581_));
 BUFx6f_ASAP7_75t_R _10384_ (.A(_03581_),
    .Y(_03582_));
 BUFx10_ASAP7_75t_R _10385_ (.A(_03125_),
    .Y(_03583_));
 AO221x1_ASAP7_75t_R _10386_ (.A1(_03571_),
    .A2(_03575_),
    .B1(_03580_),
    .B2(_03582_),
    .C(_03583_),
    .Y(_03584_));
 BUFx10_ASAP7_75t_R _10387_ (.A(_03120_),
    .Y(_03585_));
 BUFx10_ASAP7_75t_R _10388_ (.A(_03585_),
    .Y(_03586_));
 AO21x1_ASAP7_75t_R _10389_ (.A1(_03570_),
    .A2(_03584_),
    .B(_03586_),
    .Y(_03587_));
 BUFx12_ASAP7_75t_R _10390_ (.A(_03026_),
    .Y(_03588_));
 BUFx6f_ASAP7_75t_R _10391_ (.A(_03588_),
    .Y(_03589_));
 AND2x2_ASAP7_75t_R _10392_ (.A(_03037_),
    .B(_03017_),
    .Y(_03590_));
 BUFx10_ASAP7_75t_R _10393_ (.A(_03590_),
    .Y(_03591_));
 AO22x1_ASAP7_75t_R _10394_ (.A1(_03565_),
    .A2(_00035_),
    .B1(_00036_),
    .B2(_03591_),
    .Y(_03592_));
 BUFx12_ASAP7_75t_R _10395_ (.A(_03086_),
    .Y(_03593_));
 AND2x2_ASAP7_75t_R _10396_ (.A(_03039_),
    .B(_00038_),
    .Y(_03594_));
 AO21x1_ASAP7_75t_R _10397_ (.A1(_03080_),
    .A2(_00037_),
    .B(_03594_),
    .Y(_03595_));
 AO21x1_ASAP7_75t_R _10398_ (.A1(_03593_),
    .A2(_03595_),
    .B(_03077_),
    .Y(_03596_));
 BUFx10_ASAP7_75t_R _10399_ (.A(_03103_),
    .Y(_03597_));
 AND2x2_ASAP7_75t_R _10400_ (.A(_03597_),
    .B(_00035_),
    .Y(_03598_));
 AO221x1_ASAP7_75t_R _10401_ (.A1(_03589_),
    .A2(_03592_),
    .B1(_03596_),
    .B2(_03021_),
    .C(_03598_),
    .Y(_03599_));
 AND2x2_ASAP7_75t_R _10402_ (.A(_03091_),
    .B(_00042_),
    .Y(_03600_));
 AO21x1_ASAP7_75t_R _10403_ (.A1(_03573_),
    .A2(_00041_),
    .B(_03600_),
    .Y(_03601_));
 AND3x1_ASAP7_75t_R _10404_ (.A(_03578_),
    .B(_03063_),
    .C(_00040_),
    .Y(_03602_));
 AO21x1_ASAP7_75t_R _10405_ (.A1(_00039_),
    .A2(_03577_),
    .B(_03602_),
    .Y(_03603_));
 BUFx12_ASAP7_75t_R _10406_ (.A(_03121_),
    .Y(_03604_));
 AO221x2_ASAP7_75t_R _10407_ (.A1(_03571_),
    .A2(_03601_),
    .B1(_03603_),
    .B2(_03604_),
    .C(_03583_),
    .Y(_03605_));
 AO21x1_ASAP7_75t_R _10408_ (.A1(_03599_),
    .A2(_03605_),
    .B(_03119_),
    .Y(_03606_));
 AO21x1_ASAP7_75t_R _10409_ (.A1(_03587_),
    .A2(_03606_),
    .B(_03143_),
    .Y(_03607_));
 AND2x2_ASAP7_75t_R _10410_ (.A(_03072_),
    .B(_00061_),
    .Y(_03608_));
 AO21x1_ASAP7_75t_R _10411_ (.A1(_03588_),
    .A2(_00059_),
    .B(_03608_),
    .Y(_03609_));
 BUFx10_ASAP7_75t_R _10412_ (.A(net13),
    .Y(_03610_));
 AO21x1_ASAP7_75t_R _10413_ (.A1(_00062_),
    .A2(_03567_),
    .B(_03610_),
    .Y(_03611_));
 AO221x1_ASAP7_75t_R _10414_ (.A1(_00060_),
    .A2(_03560_),
    .B1(_03609_),
    .B2(_03062_),
    .C(_03611_),
    .Y(_03612_));
 AND2x2_ASAP7_75t_R _10415_ (.A(_03057_),
    .B(_00066_),
    .Y(_03613_));
 AO21x1_ASAP7_75t_R _10416_ (.A1(_03055_),
    .A2(_00065_),
    .B(_03613_),
    .Y(_03614_));
 AND3x1_ASAP7_75t_R _10417_ (.A(_03057_),
    .B(_03031_),
    .C(_00064_),
    .Y(_03615_));
 AO21x1_ASAP7_75t_R _10418_ (.A1(_00063_),
    .A2(_03123_),
    .B(_03615_),
    .Y(_03616_));
 BUFx10_ASAP7_75t_R _10419_ (.A(_03124_),
    .Y(_03617_));
 AO221x1_ASAP7_75t_R _10420_ (.A1(_03109_),
    .A2(_03614_),
    .B1(_03616_),
    .B2(_03581_),
    .C(_03617_),
    .Y(_03618_));
 AND2x2_ASAP7_75t_R _10421_ (.A(_03612_),
    .B(_03618_),
    .Y(_03619_));
 BUFx10_ASAP7_75t_R _10422_ (.A(_03572_),
    .Y(_03620_));
 AND2x2_ASAP7_75t_R _10423_ (.A(_03578_),
    .B(_00054_),
    .Y(_03621_));
 AO21x1_ASAP7_75t_R _10424_ (.A1(_03620_),
    .A2(_00053_),
    .B(_03621_),
    .Y(_03622_));
 BUFx6f_ASAP7_75t_R _10425_ (.A(_03610_),
    .Y(_03623_));
 AO21x1_ASAP7_75t_R _10426_ (.A1(_03107_),
    .A2(_03622_),
    .B(_03623_),
    .Y(_03624_));
 BUFx10_ASAP7_75t_R _10427_ (.A(_03564_),
    .Y(_03625_));
 BUFx12_ASAP7_75t_R _10428_ (.A(_03590_),
    .Y(_03626_));
 AO22x1_ASAP7_75t_R _10429_ (.A1(_03625_),
    .A2(_00051_),
    .B1(_00052_),
    .B2(_03626_),
    .Y(_03627_));
 AO22x1_ASAP7_75t_R _10430_ (.A1(_03130_),
    .A2(_00051_),
    .B1(_03627_),
    .B2(_03589_),
    .Y(_03628_));
 AO21x1_ASAP7_75t_R _10431_ (.A1(_03201_),
    .A2(_03624_),
    .B(_03628_),
    .Y(_03629_));
 BUFx10_ASAP7_75t_R _10432_ (.A(_03054_),
    .Y(_03630_));
 AND2x2_ASAP7_75t_R _10433_ (.A(_03047_),
    .B(_00058_),
    .Y(_03631_));
 AO21x1_ASAP7_75t_R _10434_ (.A1(_03630_),
    .A2(_00057_),
    .B(_03631_),
    .Y(_03632_));
 AND3x1_ASAP7_75t_R _10435_ (.A(_03047_),
    .B(_03019_),
    .C(_00056_),
    .Y(_03633_));
 AO21x1_ASAP7_75t_R _10436_ (.A1(_00055_),
    .A2(_03123_),
    .B(_03633_),
    .Y(_03634_));
 BUFx12_ASAP7_75t_R _10437_ (.A(_03121_),
    .Y(_03635_));
 BUFx6f_ASAP7_75t_R _10438_ (.A(_03125_),
    .Y(_03636_));
 AO221x1_ASAP7_75t_R _10439_ (.A1(_03109_),
    .A2(_03632_),
    .B1(_03634_),
    .B2(_03635_),
    .C(_03636_),
    .Y(_03637_));
 AND2x2_ASAP7_75t_R _10440_ (.A(_03586_),
    .B(_03637_),
    .Y(_03638_));
 AO221x1_ASAP7_75t_R _10441_ (.A1(_03119_),
    .A2(_03619_),
    .B1(_03629_),
    .B2(_03638_),
    .C(_03154_),
    .Y(_03639_));
 AO21x2_ASAP7_75t_R _10442_ (.A1(_03607_),
    .A2(_03639_),
    .B(_03127_),
    .Y(_03640_));
 INVx1_ASAP7_75t_R _10443_ (.A(net23),
    .Y(_03641_));
 OA21x2_ASAP7_75t_R _10444_ (.A1(_03099_),
    .A2(_03641_),
    .B(_03193_),
    .Y(_03642_));
 AND2x2_ASAP7_75t_R _10445_ (.A(_03270_),
    .B(_03642_),
    .Y(_03643_));
 AO21x1_ASAP7_75t_R _10446_ (.A1(_03558_),
    .A2(_03640_),
    .B(_03643_),
    .Y(_03644_));
 XNOR2x2_ASAP7_75t_R _10447_ (.A(_03557_),
    .B(_03644_),
    .Y(_09560_));
 INVx1_ASAP7_75t_R _10448_ (.A(_09560_),
    .Y(_09562_));
 BUFx6f_ASAP7_75t_R _10449_ (.A(_03270_),
    .Y(_03645_));
 AO22x1_ASAP7_75t_R _10450_ (.A1(_03061_),
    .A2(_00067_),
    .B1(_00068_),
    .B2(_03626_),
    .Y(_03646_));
 BUFx12_ASAP7_75t_R _10451_ (.A(_03085_),
    .Y(_03647_));
 AND2x2_ASAP7_75t_R _10452_ (.A(_03038_),
    .B(_00070_),
    .Y(_03648_));
 AO21x1_ASAP7_75t_R _10453_ (.A1(_03054_),
    .A2(_00069_),
    .B(_03648_),
    .Y(_03649_));
 BUFx4f_ASAP7_75t_R _10454_ (.A(net13),
    .Y(_03650_));
 AO21x1_ASAP7_75t_R _10455_ (.A1(_03647_),
    .A2(_03649_),
    .B(_03650_),
    .Y(_03651_));
 AND2x2_ASAP7_75t_R _10456_ (.A(_03096_),
    .B(_00067_),
    .Y(_03652_));
 AO221x1_ASAP7_75t_R _10457_ (.A1(_03027_),
    .A2(_03646_),
    .B1(_03651_),
    .B2(_03064_),
    .C(_03652_),
    .Y(_03653_));
 AND2x2_ASAP7_75t_R _10458_ (.A(_03039_),
    .B(_00074_),
    .Y(_03654_));
 AO21x1_ASAP7_75t_R _10459_ (.A1(_03080_),
    .A2(_00073_),
    .B(_03654_),
    .Y(_03655_));
 AND3x1_ASAP7_75t_R _10460_ (.A(_03057_),
    .B(_03031_),
    .C(_00072_),
    .Y(_03656_));
 AO21x1_ASAP7_75t_R _10461_ (.A1(_00071_),
    .A2(_03123_),
    .B(_03656_),
    .Y(_03657_));
 AO221x2_ASAP7_75t_R _10462_ (.A1(_03593_),
    .A2(_03655_),
    .B1(_03657_),
    .B2(_03581_),
    .C(_03617_),
    .Y(_03658_));
 AND3x1_ASAP7_75t_R _10463_ (.A(_03585_),
    .B(_03653_),
    .C(_03658_),
    .Y(_03659_));
 AND2x2_ASAP7_75t_R _10464_ (.A(_03039_),
    .B(_00082_),
    .Y(_03660_));
 AO21x1_ASAP7_75t_R _10465_ (.A1(_03080_),
    .A2(_00081_),
    .B(_03660_),
    .Y(_03661_));
 AND3x1_ASAP7_75t_R _10466_ (.A(_03039_),
    .B(_03031_),
    .C(_00080_),
    .Y(_03662_));
 AO21x1_ASAP7_75t_R _10467_ (.A1(_00079_),
    .A2(_03576_),
    .B(_03662_),
    .Y(_03663_));
 AO221x1_ASAP7_75t_R _10468_ (.A1(_03593_),
    .A2(_03661_),
    .B1(_03663_),
    .B2(_03581_),
    .C(_03617_),
    .Y(_03664_));
 BUFx10_ASAP7_75t_R _10469_ (.A(_03588_),
    .Y(_03665_));
 AO22x2_ASAP7_75t_R _10470_ (.A1(_03630_),
    .A2(_00075_),
    .B1(_00076_),
    .B2(_03626_),
    .Y(_03666_));
 BUFx6f_ASAP7_75t_R _10471_ (.A(_03037_),
    .Y(_03667_));
 AND2x2_ASAP7_75t_R _10472_ (.A(_03667_),
    .B(_00078_),
    .Y(_03668_));
 AO21x1_ASAP7_75t_R _10473_ (.A1(_03572_),
    .A2(_00077_),
    .B(_03668_),
    .Y(_03669_));
 AO21x1_ASAP7_75t_R _10474_ (.A1(_03073_),
    .A2(_03669_),
    .B(_03610_),
    .Y(_03670_));
 AO21x1_ASAP7_75t_R _10475_ (.A1(_03665_),
    .A2(_03666_),
    .B(_03670_),
    .Y(_03671_));
 AND3x1_ASAP7_75t_R _10476_ (.A(_03173_),
    .B(_03664_),
    .C(_03671_),
    .Y(_03672_));
 NOR3x1_ASAP7_75t_R _10477_ (.A(_03143_),
    .B(_03659_),
    .C(_03672_),
    .Y(_03673_));
 BUFx12f_ASAP7_75t_R _10478_ (.A(_03647_),
    .Y(_03674_));
 BUFx6f_ASAP7_75t_R _10479_ (.A(_03038_),
    .Y(_03675_));
 AND2x2_ASAP7_75t_R _10480_ (.A(_03675_),
    .B(_00098_),
    .Y(_03676_));
 AO21x1_ASAP7_75t_R _10481_ (.A1(_03625_),
    .A2(_00097_),
    .B(_03676_),
    .Y(_03677_));
 BUFx10_ASAP7_75t_R _10482_ (.A(_03667_),
    .Y(_03678_));
 AND3x1_ASAP7_75t_R _10483_ (.A(_03678_),
    .B(_03117_),
    .C(_00096_),
    .Y(_03679_));
 AO21x1_ASAP7_75t_R _10484_ (.A1(_00095_),
    .A2(_03289_),
    .B(_03679_),
    .Y(_03680_));
 BUFx6f_ASAP7_75t_R _10485_ (.A(_03121_),
    .Y(_03681_));
 AO221x1_ASAP7_75t_R _10486_ (.A1(_03674_),
    .A2(_03677_),
    .B1(_03680_),
    .B2(_03681_),
    .C(_03636_),
    .Y(_03682_));
 AND2x2_ASAP7_75t_R _10487_ (.A(_03072_),
    .B(_00093_),
    .Y(_03683_));
 AO21x1_ASAP7_75t_R _10488_ (.A1(_03027_),
    .A2(_00091_),
    .B(_03683_),
    .Y(_03684_));
 BUFx12_ASAP7_75t_R _10489_ (.A(_03630_),
    .Y(_03685_));
 AO21x1_ASAP7_75t_R _10490_ (.A1(_00092_),
    .A2(_03560_),
    .B(_03610_),
    .Y(_03686_));
 AO221x1_ASAP7_75t_R _10491_ (.A1(_00094_),
    .A2(_03568_),
    .B1(_03684_),
    .B2(_03685_),
    .C(_03686_),
    .Y(_03687_));
 AO21x2_ASAP7_75t_R _10492_ (.A1(_03682_),
    .A2(_03687_),
    .B(_03586_),
    .Y(_03688_));
 BUFx6f_ASAP7_75t_R _10493_ (.A(_03647_),
    .Y(_03689_));
 AND2x2_ASAP7_75t_R _10494_ (.A(_03678_),
    .B(_00090_),
    .Y(_03690_));
 AO21x1_ASAP7_75t_R _10495_ (.A1(_03625_),
    .A2(_00089_),
    .B(_03690_),
    .Y(_03691_));
 BUFx12_ASAP7_75t_R _10496_ (.A(_03667_),
    .Y(_03692_));
 AND3x1_ASAP7_75t_R _10497_ (.A(_03692_),
    .B(_03117_),
    .C(_00088_),
    .Y(_03693_));
 AO21x1_ASAP7_75t_R _10498_ (.A1(_00087_),
    .A2(_03289_),
    .B(_03693_),
    .Y(_03694_));
 BUFx10_ASAP7_75t_R _10499_ (.A(_03125_),
    .Y(_03695_));
 AO221x1_ASAP7_75t_R _10500_ (.A1(_03689_),
    .A2(_03691_),
    .B1(_03694_),
    .B2(_03681_),
    .C(_03695_),
    .Y(_03696_));
 BUFx10_ASAP7_75t_R _10501_ (.A(_03567_),
    .Y(_03697_));
 AND2x2_ASAP7_75t_R _10502_ (.A(_03086_),
    .B(_00085_),
    .Y(_03698_));
 AO21x1_ASAP7_75t_R _10503_ (.A1(_03027_),
    .A2(_00083_),
    .B(_03698_),
    .Y(_03699_));
 AO21x1_ASAP7_75t_R _10504_ (.A1(_00084_),
    .A2(_03560_),
    .B(_03610_),
    .Y(_03700_));
 AO221x1_ASAP7_75t_R _10505_ (.A1(_00086_),
    .A2(_03697_),
    .B1(_03699_),
    .B2(_03685_),
    .C(_03700_),
    .Y(_03701_));
 AO21x1_ASAP7_75t_R _10506_ (.A1(_03696_),
    .A2(_03701_),
    .B(_03173_),
    .Y(_03702_));
 BUFx6f_ASAP7_75t_R _10507_ (.A(_03154_),
    .Y(_03703_));
 AOI21x1_ASAP7_75t_R _10508_ (.A1(_03688_),
    .A2(_03702_),
    .B(_03703_),
    .Y(_03704_));
 INVx8_ASAP7_75t_R _10509_ (.A(_03126_),
    .Y(_03705_));
 OAI21x1_ASAP7_75t_R _10510_ (.A1(_03673_),
    .A2(_03704_),
    .B(_03705_),
    .Y(_03706_));
 BUFx4f_ASAP7_75t_R _10511_ (.A(_03270_),
    .Y(_03707_));
 AO21x2_ASAP7_75t_R _10512_ (.A1(_03209_),
    .A2(_03227_),
    .B(_03248_),
    .Y(_03708_));
 NAND2x1_ASAP7_75t_R _10513_ (.A(_03708_),
    .B(_03275_),
    .Y(_03709_));
 OA21x2_ASAP7_75t_R _10514_ (.A1(_03708_),
    .A2(_03642_),
    .B(_03709_),
    .Y(_03710_));
 OA21x2_ASAP7_75t_R _10515_ (.A1(_03265_),
    .A2(_03642_),
    .B(_03710_),
    .Y(_03711_));
 BUFx4f_ASAP7_75t_R _10516_ (.A(_03711_),
    .Y(_03712_));
 BUFx4f_ASAP7_75t_R _10517_ (.A(_03099_),
    .Y(_03713_));
 INVx3_ASAP7_75t_R _10518_ (.A(net22),
    .Y(_03714_));
 BUFx3_ASAP7_75t_R _10519_ (.A(_03247_),
    .Y(_03715_));
 OR3x1_ASAP7_75t_R _10520_ (.A(_03713_),
    .B(_03714_),
    .C(_03715_),
    .Y(_03716_));
 AND3x1_ASAP7_75t_R _10521_ (.A(_03708_),
    .B(_03275_),
    .C(_03642_),
    .Y(_03717_));
 BUFx4f_ASAP7_75t_R _10522_ (.A(_03717_),
    .Y(_03718_));
 AOI21x1_ASAP7_75t_R _10523_ (.A1(_03712_),
    .A2(_03716_),
    .B(_03718_),
    .Y(_09776_));
 NAND2x1_ASAP7_75t_R _10524_ (.A(_03707_),
    .B(_09776_),
    .Y(_03719_));
 OA21x2_ASAP7_75t_R _10525_ (.A1(_03645_),
    .A2(_03706_),
    .B(_03719_),
    .Y(_03720_));
 XNOR2x2_ASAP7_75t_R _10526_ (.A(_03557_),
    .B(_03720_),
    .Y(_09566_));
 INVx1_ASAP7_75t_R _10527_ (.A(_09566_),
    .Y(_09568_));
 INVx1_ASAP7_75t_R _10528_ (.A(_00092_),
    .Y(_03721_));
 BUFx12_ASAP7_75t_R _10529_ (.A(_03431_),
    .Y(_03722_));
 NAND2x1_ASAP7_75t_R _10530_ (.A(_00091_),
    .B(_03414_),
    .Y(_03723_));
 OA211x2_ASAP7_75t_R _10531_ (.A1(_03721_),
    .A2(_03722_),
    .B(_03447_),
    .C(_03723_),
    .Y(_03724_));
 OA22x2_ASAP7_75t_R _10532_ (.A1(_00093_),
    .A2(_03522_),
    .B1(_03485_),
    .B2(_00094_),
    .Y(_03725_));
 AND3x1_ASAP7_75t_R _10533_ (.A(_03043_),
    .B(_03474_),
    .C(_00098_),
    .Y(_03726_));
 AO221x1_ASAP7_75t_R _10534_ (.A1(_03260_),
    .A2(_03506_),
    .B1(_03465_),
    .B2(_00097_),
    .C(_03726_),
    .Y(_03727_));
 OAI21x1_ASAP7_75t_R _10535_ (.A1(_03440_),
    .A2(_03725_),
    .B(_03727_),
    .Y(_03728_));
 OAI22x1_ASAP7_75t_R _10536_ (.A1(_00096_),
    .A2(_03396_),
    .B1(_03511_),
    .B2(_00095_),
    .Y(_03729_));
 AO221x1_ASAP7_75t_R _10537_ (.A1(_03340_),
    .A2(_03728_),
    .B1(_03729_),
    .B2(_03482_),
    .C(_03404_),
    .Y(_03730_));
 AO21x2_ASAP7_75t_R _10538_ (.A1(_03371_),
    .A2(_03386_),
    .B(_03332_),
    .Y(_03731_));
 BUFx12f_ASAP7_75t_R _10539_ (.A(_03731_),
    .Y(_03732_));
 NAND2x2_ASAP7_75t_R _10540_ (.A(_03319_),
    .B(_03398_),
    .Y(_03733_));
 OAI22x1_ASAP7_75t_R _10541_ (.A1(_00090_),
    .A2(_03732_),
    .B1(_03733_),
    .B2(_00086_),
    .Y(_03734_));
 BUFx12_ASAP7_75t_R _10542_ (.A(_03522_),
    .Y(_03735_));
 BUFx12f_ASAP7_75t_R _10543_ (.A(_03386_),
    .Y(_03736_));
 AND3x1_ASAP7_75t_R _10544_ (.A(_00085_),
    .B(_03208_),
    .C(_03736_),
    .Y(_03737_));
 AOI211x1_ASAP7_75t_R _10545_ (.A1(_00089_),
    .A2(_03504_),
    .B(_03735_),
    .C(_03737_),
    .Y(_03738_));
 OA21x2_ASAP7_75t_R _10546_ (.A1(_03734_),
    .A2(_03738_),
    .B(_03443_),
    .Y(_03739_));
 BUFx12f_ASAP7_75t_R _10547_ (.A(_03485_),
    .Y(_03740_));
 NAND2x1_ASAP7_75t_R _10548_ (.A(_00083_),
    .B(_03740_),
    .Y(_03741_));
 NAND2x1_ASAP7_75t_R _10549_ (.A(_00084_),
    .B(_03454_),
    .Y(_03742_));
 OAI22x1_ASAP7_75t_R _10550_ (.A1(_00087_),
    .A2(_03313_),
    .B1(_03449_),
    .B2(_00088_),
    .Y(_03743_));
 AO21x1_ASAP7_75t_R _10551_ (.A1(_03361_),
    .A2(_03743_),
    .B(_03460_),
    .Y(_03744_));
 AO32x2_ASAP7_75t_R _10552_ (.A1(_03447_),
    .A2(_03741_),
    .A3(_03742_),
    .B1(_03744_),
    .B2(_03245_),
    .Y(_03745_));
 OA22x2_ASAP7_75t_R _10553_ (.A1(_03724_),
    .A2(_03730_),
    .B1(_03739_),
    .B2(_03745_),
    .Y(_03746_));
 BUFx12f_ASAP7_75t_R _10554_ (.A(_03503_),
    .Y(_03747_));
 AND2x6_ASAP7_75t_R _10555_ (.A(_03351_),
    .B(_03352_),
    .Y(_03748_));
 CKINVDCx12_ASAP7_75t_R _10556_ (.A(_03301_),
    .Y(_03749_));
 OR3x1_ASAP7_75t_R _10557_ (.A(_03103_),
    .B(_03749_),
    .C(_00070_),
    .Y(_03750_));
 OA22x2_ASAP7_75t_R _10558_ (.A1(_00069_),
    .A2(_03305_),
    .B1(_03748_),
    .B2(_03750_),
    .Y(_03751_));
 AND2x2_ASAP7_75t_R _10559_ (.A(_00073_),
    .B(_03435_),
    .Y(_03752_));
 AO221x2_ASAP7_75t_R _10560_ (.A1(_03324_),
    .A2(_03387_),
    .B1(_03522_),
    .B2(_00074_),
    .C(_03752_),
    .Y(_03753_));
 OAI21x1_ASAP7_75t_R _10561_ (.A1(_03747_),
    .A2(_03751_),
    .B(_03753_),
    .Y(_03754_));
 AND3x1_ASAP7_75t_R _10562_ (.A(_03245_),
    .B(_03502_),
    .C(_03754_),
    .Y(_03755_));
 NAND2x1_ASAP7_75t_R _10563_ (.A(_00067_),
    .B(_03740_),
    .Y(_03756_));
 NAND2x1_ASAP7_75t_R _10564_ (.A(_00068_),
    .B(_03511_),
    .Y(_03757_));
 INVx1_ASAP7_75t_R _10565_ (.A(_00071_),
    .Y(_03758_));
 NAND2x2_ASAP7_75t_R _10566_ (.A(_03351_),
    .B(_03352_),
    .Y(_03759_));
 NOR2x1_ASAP7_75t_R _10567_ (.A(_00072_),
    .B(_03435_),
    .Y(_03760_));
 AO22x1_ASAP7_75t_R _10568_ (.A1(_03758_),
    .A2(_03395_),
    .B1(_03759_),
    .B2(_03760_),
    .Y(_03761_));
 AO21x2_ASAP7_75t_R _10569_ (.A1(_03361_),
    .A2(_03761_),
    .B(_03460_),
    .Y(_03762_));
 AO32x1_ASAP7_75t_R _10570_ (.A1(_03447_),
    .A2(_03756_),
    .A3(_03757_),
    .B1(_03762_),
    .B2(_03245_),
    .Y(_03763_));
 INVx1_ASAP7_75t_R _10571_ (.A(_00076_),
    .Y(_03764_));
 BUFx12f_ASAP7_75t_R _10572_ (.A(_03413_),
    .Y(_03765_));
 NAND2x1_ASAP7_75t_R _10573_ (.A(_00075_),
    .B(_03765_),
    .Y(_03766_));
 OA211x2_ASAP7_75t_R _10574_ (.A1(_03764_),
    .A2(_03722_),
    .B(_03447_),
    .C(_03766_),
    .Y(_03767_));
 OA22x2_ASAP7_75t_R _10575_ (.A1(_00077_),
    .A2(_03522_),
    .B1(_03485_),
    .B2(_00078_),
    .Y(_03768_));
 AND2x2_ASAP7_75t_R _10576_ (.A(_00081_),
    .B(_03333_),
    .Y(_03769_));
 AO221x1_ASAP7_75t_R _10577_ (.A1(_03260_),
    .A2(_03506_),
    .B1(_03507_),
    .B2(_00082_),
    .C(_03769_),
    .Y(_03770_));
 OAI21x1_ASAP7_75t_R _10578_ (.A1(_03440_),
    .A2(_03768_),
    .B(_03770_),
    .Y(_03771_));
 OAI22x1_ASAP7_75t_R _10579_ (.A1(_00080_),
    .A2(_03396_),
    .B1(_03400_),
    .B2(_00079_),
    .Y(_03772_));
 AO221x1_ASAP7_75t_R _10580_ (.A1(_03340_),
    .A2(_03771_),
    .B1(_03772_),
    .B2(_03482_),
    .C(_03404_),
    .Y(_03773_));
 OA22x2_ASAP7_75t_R _10581_ (.A1(_03755_),
    .A2(_03763_),
    .B1(_03767_),
    .B2(_03773_),
    .Y(_03774_));
 AO32x1_ASAP7_75t_R _10582_ (.A1(_03247_),
    .A2(_03539_),
    .A3(_03746_),
    .B1(_03774_),
    .B2(_03499_),
    .Y(_03775_));
 BUFx6f_ASAP7_75t_R _10583_ (.A(_03775_),
    .Y(_09565_));
 INVx1_ASAP7_75t_R _10584_ (.A(_09565_),
    .Y(_09567_));
 INVx1_ASAP7_75t_R _10585_ (.A(net20),
    .Y(_03776_));
 BUFx3_ASAP7_75t_R _10586_ (.A(_03715_),
    .Y(_03777_));
 OR3x1_ASAP7_75t_R _10587_ (.A(_03713_),
    .B(_03776_),
    .C(_03777_),
    .Y(_03778_));
 BUFx6f_ASAP7_75t_R _10588_ (.A(_03718_),
    .Y(_03779_));
 AOI21x1_ASAP7_75t_R _10589_ (.A1(_03712_),
    .A2(_03778_),
    .B(_03779_),
    .Y(_09774_));
 BUFx4f_ASAP7_75t_R _10590_ (.A(_03270_),
    .Y(_03780_));
 BUFx10_ASAP7_75t_R _10591_ (.A(_03127_),
    .Y(_03781_));
 AO22x1_ASAP7_75t_R _10592_ (.A1(_03564_),
    .A2(_00101_),
    .B1(_00102_),
    .B2(_03590_),
    .Y(_03782_));
 AND2x2_ASAP7_75t_R _10593_ (.A(_03037_),
    .B(_00104_),
    .Y(_03783_));
 AO21x1_ASAP7_75t_R _10594_ (.A1(_03054_),
    .A2(_00103_),
    .B(_03783_),
    .Y(_03784_));
 AO21x1_ASAP7_75t_R _10595_ (.A1(_03086_),
    .A2(_03784_),
    .B(_03650_),
    .Y(_03785_));
 AND2x2_ASAP7_75t_R _10596_ (.A(_03103_),
    .B(_00101_),
    .Y(_03786_));
 AO221x1_ASAP7_75t_R _10597_ (.A1(_03588_),
    .A2(_03782_),
    .B1(_03785_),
    .B2(_03473_),
    .C(_03786_),
    .Y(_03787_));
 AND2x2_ASAP7_75t_R _10598_ (.A(_03667_),
    .B(_00108_),
    .Y(_03788_));
 AO21x1_ASAP7_75t_R _10599_ (.A1(_03564_),
    .A2(_00107_),
    .B(_03788_),
    .Y(_03789_));
 AND3x1_ASAP7_75t_R _10600_ (.A(_03090_),
    .B(_03116_),
    .C(_00106_),
    .Y(_03790_));
 AO21x1_ASAP7_75t_R _10601_ (.A1(_00105_),
    .A2(_03576_),
    .B(_03790_),
    .Y(_03791_));
 AO221x1_ASAP7_75t_R _10602_ (.A1(_03088_),
    .A2(_03789_),
    .B1(_03791_),
    .B2(_03581_),
    .C(_03125_),
    .Y(_03792_));
 AND3x1_ASAP7_75t_R _10603_ (.A(_03585_),
    .B(_03787_),
    .C(_03792_),
    .Y(_03793_));
 AND2x2_ASAP7_75t_R _10604_ (.A(_03667_),
    .B(_00116_),
    .Y(_03794_));
 AO21x1_ASAP7_75t_R _10605_ (.A1(_03564_),
    .A2(_00115_),
    .B(_03794_),
    .Y(_03795_));
 AND3x1_ASAP7_75t_R _10606_ (.A(_03667_),
    .B(_03116_),
    .C(_00114_),
    .Y(_03796_));
 AO21x1_ASAP7_75t_R _10607_ (.A1(_00113_),
    .A2(_03576_),
    .B(_03796_),
    .Y(_03797_));
 AO221x1_ASAP7_75t_R _10608_ (.A1(_03088_),
    .A2(_03795_),
    .B1(_03797_),
    .B2(_03121_),
    .C(_03125_),
    .Y(_03798_));
 AO22x1_ASAP7_75t_R _10609_ (.A1(_03061_),
    .A2(_00109_),
    .B1(_00110_),
    .B2(_03626_),
    .Y(_03799_));
 AND2x2_ASAP7_75t_R _10610_ (.A(_03038_),
    .B(_00112_),
    .Y(_03800_));
 AO21x1_ASAP7_75t_R _10611_ (.A1(_03054_),
    .A2(_00111_),
    .B(_03800_),
    .Y(_03801_));
 AO21x1_ASAP7_75t_R _10612_ (.A1(_03647_),
    .A2(_03801_),
    .B(_03650_),
    .Y(_03802_));
 AO21x1_ASAP7_75t_R _10613_ (.A1(_03160_),
    .A2(_03799_),
    .B(_03802_),
    .Y(_03803_));
 AND3x1_ASAP7_75t_R _10614_ (.A(_03118_),
    .B(_03798_),
    .C(_03803_),
    .Y(_03804_));
 OR3x1_ASAP7_75t_R _10615_ (.A(_03142_),
    .B(_03793_),
    .C(_03804_),
    .Y(_03805_));
 BUFx6f_ASAP7_75t_R _10616_ (.A(_03072_),
    .Y(_03806_));
 BUFx10_ASAP7_75t_R _10617_ (.A(_03037_),
    .Y(_03807_));
 AND2x2_ASAP7_75t_R _10618_ (.A(_03807_),
    .B(_00132_),
    .Y(_03808_));
 AO21x1_ASAP7_75t_R _10619_ (.A1(_03080_),
    .A2(_00131_),
    .B(_03808_),
    .Y(_03809_));
 AND3x1_ASAP7_75t_R _10620_ (.A(_03039_),
    .B(_03031_),
    .C(_00130_),
    .Y(_03810_));
 AO21x1_ASAP7_75t_R _10621_ (.A1(_00129_),
    .A2(_03576_),
    .B(_03810_),
    .Y(_03811_));
 AO221x1_ASAP7_75t_R _10622_ (.A1(_03806_),
    .A2(_03809_),
    .B1(_03811_),
    .B2(_03581_),
    .C(_03617_),
    .Y(_03812_));
 AND2x2_ASAP7_75t_R _10623_ (.A(_03085_),
    .B(_00127_),
    .Y(_03813_));
 AO21x1_ASAP7_75t_R _10624_ (.A1(_03026_),
    .A2(_00125_),
    .B(_03813_),
    .Y(_03814_));
 AO21x1_ASAP7_75t_R _10625_ (.A1(_00126_),
    .A2(_03559_),
    .B(_03650_),
    .Y(_03815_));
 AO221x1_ASAP7_75t_R _10626_ (.A1(_00128_),
    .A2(_03568_),
    .B1(_03814_),
    .B2(_03620_),
    .C(_03815_),
    .Y(_03816_));
 AO21x1_ASAP7_75t_R _10627_ (.A1(_03812_),
    .A2(_03816_),
    .B(_03585_),
    .Y(_03817_));
 AND2x2_ASAP7_75t_R _10628_ (.A(_03807_),
    .B(_00124_),
    .Y(_03818_));
 AO21x1_ASAP7_75t_R _10629_ (.A1(_03080_),
    .A2(_00123_),
    .B(_03818_),
    .Y(_03819_));
 AND3x1_ASAP7_75t_R _10630_ (.A(_03039_),
    .B(_03043_),
    .C(_00122_),
    .Y(_03820_));
 AO21x1_ASAP7_75t_R _10631_ (.A1(_00121_),
    .A2(_03576_),
    .B(_03820_),
    .Y(_03821_));
 AO221x1_ASAP7_75t_R _10632_ (.A1(_03806_),
    .A2(_03819_),
    .B1(_03821_),
    .B2(_03581_),
    .C(_03617_),
    .Y(_03822_));
 AND2x2_ASAP7_75t_R _10633_ (.A(_03085_),
    .B(_00119_),
    .Y(_03823_));
 AO21x1_ASAP7_75t_R _10634_ (.A1(_03026_),
    .A2(_00117_),
    .B(_03823_),
    .Y(_03824_));
 AO21x1_ASAP7_75t_R _10635_ (.A1(_00118_),
    .A2(_03559_),
    .B(_03650_),
    .Y(_03825_));
 AO221x1_ASAP7_75t_R _10636_ (.A1(_00120_),
    .A2(_03568_),
    .B1(_03824_),
    .B2(_03620_),
    .C(_03825_),
    .Y(_03826_));
 AO21x1_ASAP7_75t_R _10637_ (.A1(_03822_),
    .A2(_03826_),
    .B(_03173_),
    .Y(_03827_));
 AO21x1_ASAP7_75t_R _10638_ (.A1(_03817_),
    .A2(_03827_),
    .B(_03154_),
    .Y(_03828_));
 AND2x4_ASAP7_75t_R _10639_ (.A(_03805_),
    .B(_03828_),
    .Y(_03829_));
 OR2x4_ASAP7_75t_R _10640_ (.A(_03781_),
    .B(_03829_),
    .Y(_03830_));
 NOR2x1_ASAP7_75t_R _10641_ (.A(_03780_),
    .B(_03830_),
    .Y(_03831_));
 AOI21x1_ASAP7_75t_R _10642_ (.A1(_03645_),
    .A2(_09774_),
    .B(_03831_),
    .Y(_03832_));
 XNOR2x2_ASAP7_75t_R _10643_ (.A(_03557_),
    .B(_03832_),
    .Y(_09571_));
 INVx1_ASAP7_75t_R _10644_ (.A(_09571_),
    .Y(_09573_));
 OAI22x1_ASAP7_75t_R _10645_ (.A1(_00121_),
    .A2(_03349_),
    .B1(_03356_),
    .B2(_00122_),
    .Y(_03833_));
 AND2x2_ASAP7_75t_R _10646_ (.A(_03482_),
    .B(_03833_),
    .Y(_03834_));
 AND3x4_ASAP7_75t_R _10647_ (.A(_03260_),
    .B(_03298_),
    .C(_03338_),
    .Y(_03835_));
 AO21x2_ASAP7_75t_R _10648_ (.A1(_03233_),
    .A2(_03243_),
    .B(_03835_),
    .Y(_03836_));
 BUFx10_ASAP7_75t_R _10649_ (.A(_03303_),
    .Y(_03837_));
 OA22x2_ASAP7_75t_R _10650_ (.A1(_00119_),
    .A2(_03837_),
    .B1(_03355_),
    .B2(_00120_),
    .Y(_03838_));
 AND2x2_ASAP7_75t_R _10651_ (.A(_00123_),
    .B(_03332_),
    .Y(_03839_));
 AO221x1_ASAP7_75t_R _10652_ (.A1(_03207_),
    .A2(_03320_),
    .B1(_03304_),
    .B2(_00124_),
    .C(_03839_),
    .Y(_03840_));
 OA211x2_ASAP7_75t_R _10653_ (.A1(_03440_),
    .A2(_03838_),
    .B(_03840_),
    .C(_03298_),
    .Y(_03841_));
 AND2x2_ASAP7_75t_R _10654_ (.A(_00118_),
    .B(_03453_),
    .Y(_03842_));
 AO21x1_ASAP7_75t_R _10655_ (.A1(_00117_),
    .A2(_03356_),
    .B(_03842_),
    .Y(_03843_));
 OA21x2_ASAP7_75t_R _10656_ (.A1(_03272_),
    .A2(_03286_),
    .B(_03373_),
    .Y(_03844_));
 BUFx6f_ASAP7_75t_R _10657_ (.A(_03844_),
    .Y(_03845_));
 OAI22x1_ASAP7_75t_R _10658_ (.A1(_03836_),
    .A2(_03841_),
    .B1(_03843_),
    .B2(_03845_),
    .Y(_03846_));
 BUFx12f_ASAP7_75t_R _10659_ (.A(_03465_),
    .Y(_03847_));
 OAI22x1_ASAP7_75t_R _10660_ (.A1(_00130_),
    .A2(_03847_),
    .B1(_03467_),
    .B2(_00129_),
    .Y(_03848_));
 AND3x1_ASAP7_75t_R _10661_ (.A(_03422_),
    .B(_03482_),
    .C(_03848_),
    .Y(_03849_));
 AND3x1_ASAP7_75t_R _10662_ (.A(_03116_),
    .B(_03474_),
    .C(_00132_),
    .Y(_03850_));
 AO21x1_ASAP7_75t_R _10663_ (.A1(_00131_),
    .A2(_03465_),
    .B(_03850_),
    .Y(_03851_));
 OA21x2_ASAP7_75t_R _10664_ (.A1(_00127_),
    .A2(_03327_),
    .B(_03386_),
    .Y(_03852_));
 OA21x2_ASAP7_75t_R _10665_ (.A1(_00128_),
    .A2(_03355_),
    .B(_03852_),
    .Y(_03853_));
 AND2x2_ASAP7_75t_R _10666_ (.A(_03206_),
    .B(_03338_),
    .Y(_03854_));
 BUFx10_ASAP7_75t_R _10667_ (.A(_03854_),
    .Y(_03855_));
 AO221x1_ASAP7_75t_R _10668_ (.A1(_03440_),
    .A2(_03851_),
    .B1(_03853_),
    .B2(_03371_),
    .C(_03855_),
    .Y(_03856_));
 OA211x2_ASAP7_75t_R _10669_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03327_),
    .C(_00126_),
    .Y(_03857_));
 AO21x1_ASAP7_75t_R _10670_ (.A1(_00125_),
    .A2(_03485_),
    .B(_03857_),
    .Y(_03858_));
 OA21x2_ASAP7_75t_R _10671_ (.A1(_03373_),
    .A2(_03858_),
    .B(_03460_),
    .Y(_03859_));
 BUFx10_ASAP7_75t_R _10672_ (.A(_03116_),
    .Y(_03860_));
 NAND2x2_ASAP7_75t_R _10673_ (.A(_03860_),
    .B(net10),
    .Y(_03861_));
 AO21x2_ASAP7_75t_R _10674_ (.A1(_03233_),
    .A2(_03243_),
    .B(_03861_),
    .Y(_03862_));
 AOI21x1_ASAP7_75t_R _10675_ (.A1(_03856_),
    .A2(_03859_),
    .B(_03862_),
    .Y(_03863_));
 OA22x2_ASAP7_75t_R _10676_ (.A1(_03834_),
    .A2(_03846_),
    .B1(_03849_),
    .B2(_03863_),
    .Y(_03864_));
 NAND2x2_ASAP7_75t_R _10677_ (.A(_03338_),
    .B(_03359_),
    .Y(_03865_));
 OA22x2_ASAP7_75t_R _10678_ (.A1(_00105_),
    .A2(_03328_),
    .B1(_03413_),
    .B2(_00106_),
    .Y(_03866_));
 AND2x2_ASAP7_75t_R _10679_ (.A(_00101_),
    .B(_03413_),
    .Y(_03867_));
 AND2x2_ASAP7_75t_R _10680_ (.A(_00102_),
    .B(_03453_),
    .Y(_03868_));
 OA33x2_ASAP7_75t_R _10681_ (.A1(_03344_),
    .A2(_03865_),
    .A3(_03866_),
    .B1(_03867_),
    .B2(_03868_),
    .B3(_03845_),
    .Y(_03869_));
 AND3x1_ASAP7_75t_R _10682_ (.A(_03043_),
    .B(_03474_),
    .C(_00108_),
    .Y(_03870_));
 AOI221x1_ASAP7_75t_R _10683_ (.A1(_03250_),
    .A2(_03387_),
    .B1(_03334_),
    .B2(_00107_),
    .C(_03870_),
    .Y(_03871_));
 INVx1_ASAP7_75t_R _10684_ (.A(_00104_),
    .Y(_03872_));
 OA211x2_ASAP7_75t_R _10685_ (.A1(_03197_),
    .A2(_03309_),
    .B(_03347_),
    .C(_03872_),
    .Y(_03873_));
 NOR2x1_ASAP7_75t_R _10686_ (.A(_00103_),
    .B(_03304_),
    .Y(_03874_));
 OA211x2_ASAP7_75t_R _10687_ (.A1(_03873_),
    .A2(_03874_),
    .B(_03260_),
    .C(_03320_),
    .Y(_03875_));
 OAI21x1_ASAP7_75t_R _10688_ (.A1(_03871_),
    .A2(_03875_),
    .B(_03501_),
    .Y(_03876_));
 AO21x1_ASAP7_75t_R _10689_ (.A1(_03550_),
    .A2(_03876_),
    .B(_03344_),
    .Y(_03877_));
 OAI22x1_ASAP7_75t_R _10690_ (.A1(_00114_),
    .A2(_03396_),
    .B1(_03511_),
    .B2(_00113_),
    .Y(_03878_));
 NAND2x1_ASAP7_75t_R _10691_ (.A(_03516_),
    .B(_03878_),
    .Y(_03879_));
 OR3x1_ASAP7_75t_R _10692_ (.A(_03095_),
    .B(_03749_),
    .C(_00112_),
    .Y(_03880_));
 OA22x2_ASAP7_75t_R _10693_ (.A1(_00111_),
    .A2(_03312_),
    .B1(_03748_),
    .B2(_03880_),
    .Y(_03881_));
 AND3x1_ASAP7_75t_R _10694_ (.A(_03018_),
    .B(_03301_),
    .C(_00116_),
    .Y(_03882_));
 AO221x1_ASAP7_75t_R _10695_ (.A1(_03207_),
    .A2(_03386_),
    .B1(_03333_),
    .B2(_00115_),
    .C(_03882_),
    .Y(_03883_));
 OA21x2_ASAP7_75t_R _10696_ (.A1(_03503_),
    .A2(_03881_),
    .B(_03883_),
    .Y(_03884_));
 AND2x2_ASAP7_75t_R _10697_ (.A(_00109_),
    .B(_03430_),
    .Y(_03885_));
 AND2x2_ASAP7_75t_R _10698_ (.A(_00110_),
    .B(_03399_),
    .Y(_03886_));
 OR3x1_ASAP7_75t_R _10699_ (.A(_03373_),
    .B(_03885_),
    .C(_03886_),
    .Y(_03887_));
 OA21x2_ASAP7_75t_R _10700_ (.A1(_03272_),
    .A2(_03286_),
    .B(_03459_),
    .Y(_03888_));
 OA211x2_ASAP7_75t_R _10701_ (.A1(_03855_),
    .A2(_03884_),
    .B(_03887_),
    .C(_03888_),
    .Y(_03889_));
 AOI221x1_ASAP7_75t_R _10702_ (.A1(_03869_),
    .A2(_03877_),
    .B1(_03879_),
    .B2(_03889_),
    .C(_03425_),
    .Y(_03890_));
 OR2x2_ASAP7_75t_R _10703_ (.A(_03864_),
    .B(_03890_),
    .Y(_03891_));
 BUFx6f_ASAP7_75t_R _10704_ (.A(_03891_),
    .Y(_09570_));
 INVx1_ASAP7_75t_R _10705_ (.A(_09570_),
    .Y(_09572_));
 OR2x2_ASAP7_75t_R _10706_ (.A(_03119_),
    .B(_03127_),
    .Y(_03892_));
 BUFx6f_ASAP7_75t_R _10707_ (.A(_03109_),
    .Y(_03893_));
 BUFx10_ASAP7_75t_R _10708_ (.A(_03047_),
    .Y(_03894_));
 AND2x2_ASAP7_75t_R _10709_ (.A(_03894_),
    .B(_00157_),
    .Y(_03895_));
 AO21x1_ASAP7_75t_R _10710_ (.A1(_03685_),
    .A2(_00156_),
    .B(_03895_),
    .Y(_03896_));
 BUFx10_ASAP7_75t_R _10711_ (.A(_03123_),
    .Y(_03897_));
 BUFx10_ASAP7_75t_R _10712_ (.A(_03047_),
    .Y(_03898_));
 AND3x1_ASAP7_75t_R _10713_ (.A(_03898_),
    .B(_03473_),
    .C(_00155_),
    .Y(_03899_));
 AO21x1_ASAP7_75t_R _10714_ (.A1(_00154_),
    .A2(_03897_),
    .B(_03899_),
    .Y(_03900_));
 BUFx6f_ASAP7_75t_R _10715_ (.A(_03635_),
    .Y(_03901_));
 BUFx6f_ASAP7_75t_R _10716_ (.A(_03636_),
    .Y(_03902_));
 AO221x1_ASAP7_75t_R _10717_ (.A1(_03893_),
    .A2(_03896_),
    .B1(_03900_),
    .B2(_03901_),
    .C(_03902_),
    .Y(_03903_));
 BUFx6f_ASAP7_75t_R _10718_ (.A(_03589_),
    .Y(_03904_));
 BUFx10_ASAP7_75t_R _10719_ (.A(_03630_),
    .Y(_03905_));
 BUFx10_ASAP7_75t_R _10720_ (.A(_03626_),
    .Y(_03906_));
 AO22x1_ASAP7_75t_R _10721_ (.A1(_03905_),
    .A2(_00150_),
    .B1(_00151_),
    .B2(_03906_),
    .Y(_03907_));
 AND2x6_ASAP7_75t_R _10722_ (.A(_03085_),
    .B(_03116_),
    .Y(_03908_));
 BUFx12f_ASAP7_75t_R _10723_ (.A(_03908_),
    .Y(_03909_));
 BUFx12f_ASAP7_75t_R _10724_ (.A(_03564_),
    .Y(_03910_));
 AND2x2_ASAP7_75t_R _10725_ (.A(_03692_),
    .B(_00153_),
    .Y(_03911_));
 AO21x1_ASAP7_75t_R _10726_ (.A1(_03910_),
    .A2(_00152_),
    .B(_03911_),
    .Y(_03912_));
 AND2x2_ASAP7_75t_R _10727_ (.A(net13),
    .B(_03116_),
    .Y(_03913_));
 BUFx6f_ASAP7_75t_R _10728_ (.A(_03913_),
    .Y(_03914_));
 AO221x1_ASAP7_75t_R _10729_ (.A1(_03097_),
    .A2(_00150_),
    .B1(_03909_),
    .B2(_03912_),
    .C(_03914_),
    .Y(_03915_));
 AO21x1_ASAP7_75t_R _10730_ (.A1(_03904_),
    .A2(_03907_),
    .B(_03915_),
    .Y(_03916_));
 AND3x1_ASAP7_75t_R _10731_ (.A(_03143_),
    .B(_03903_),
    .C(_03916_),
    .Y(_03917_));
 AND2x2_ASAP7_75t_R _10732_ (.A(_03894_),
    .B(_00141_),
    .Y(_03918_));
 AO21x1_ASAP7_75t_R _10733_ (.A1(_03685_),
    .A2(_00140_),
    .B(_03918_),
    .Y(_03919_));
 AND3x1_ASAP7_75t_R _10734_ (.A(_03898_),
    .B(_03473_),
    .C(_00139_),
    .Y(_03920_));
 AO21x1_ASAP7_75t_R _10735_ (.A1(_00138_),
    .A2(_03897_),
    .B(_03920_),
    .Y(_03921_));
 BUFx6f_ASAP7_75t_R _10736_ (.A(_03635_),
    .Y(_03922_));
 AO221x2_ASAP7_75t_R _10737_ (.A1(_03893_),
    .A2(_03919_),
    .B1(_03921_),
    .B2(_03922_),
    .C(_03902_),
    .Y(_03923_));
 AO22x1_ASAP7_75t_R _10738_ (.A1(_03566_),
    .A2(_00134_),
    .B1(_00135_),
    .B2(_03906_),
    .Y(_03924_));
 BUFx10_ASAP7_75t_R _10739_ (.A(_03908_),
    .Y(_03925_));
 BUFx10_ASAP7_75t_R _10740_ (.A(_03667_),
    .Y(_03926_));
 AND2x2_ASAP7_75t_R _10741_ (.A(_03926_),
    .B(_00137_),
    .Y(_03927_));
 AO21x2_ASAP7_75t_R _10742_ (.A1(_03910_),
    .A2(_00136_),
    .B(_03927_),
    .Y(_03928_));
 AO221x1_ASAP7_75t_R _10743_ (.A1(_03130_),
    .A2(_00134_),
    .B1(_03925_),
    .B2(_03928_),
    .C(_03914_),
    .Y(_03929_));
 AO21x1_ASAP7_75t_R _10744_ (.A1(_03904_),
    .A2(_03924_),
    .B(_03929_),
    .Y(_03930_));
 AND3x1_ASAP7_75t_R _10745_ (.A(_03703_),
    .B(_03923_),
    .C(_03930_),
    .Y(_03931_));
 BUFx10_ASAP7_75t_R _10746_ (.A(_03572_),
    .Y(_03932_));
 AO22x1_ASAP7_75t_R _10747_ (.A1(_03932_),
    .A2(_00158_),
    .B1(_00159_),
    .B2(_03591_),
    .Y(_03933_));
 AND2x2_ASAP7_75t_R _10748_ (.A(_03090_),
    .B(_00161_),
    .Y(_03934_));
 AO21x1_ASAP7_75t_R _10749_ (.A1(_03572_),
    .A2(_00160_),
    .B(_03934_),
    .Y(_03935_));
 BUFx10_ASAP7_75t_R _10750_ (.A(_03913_),
    .Y(_03936_));
 AO221x1_ASAP7_75t_R _10751_ (.A1(_03104_),
    .A2(_00158_),
    .B1(_03908_),
    .B2(_03935_),
    .C(_03936_),
    .Y(_03937_));
 AO21x1_ASAP7_75t_R _10752_ (.A1(_03132_),
    .A2(_03933_),
    .B(_03937_),
    .Y(_03938_));
 AND2x2_ASAP7_75t_R _10753_ (.A(_03675_),
    .B(_00165_),
    .Y(_03939_));
 AO21x1_ASAP7_75t_R _10754_ (.A1(_03111_),
    .A2(_00164_),
    .B(_03939_),
    .Y(_03940_));
 AND3x1_ASAP7_75t_R _10755_ (.A(_03678_),
    .B(_03117_),
    .C(_00163_),
    .Y(_03941_));
 AO21x1_ASAP7_75t_R _10756_ (.A1(_00162_),
    .A2(_03123_),
    .B(_03941_),
    .Y(_03942_));
 AO221x1_ASAP7_75t_R _10757_ (.A1(_03674_),
    .A2(_03940_),
    .B1(_03942_),
    .B2(_03635_),
    .C(_03636_),
    .Y(_03943_));
 AND2x2_ASAP7_75t_R _10758_ (.A(_03938_),
    .B(_03943_),
    .Y(_03944_));
 BUFx10_ASAP7_75t_R _10759_ (.A(_03061_),
    .Y(_03945_));
 BUFx12f_ASAP7_75t_R _10760_ (.A(_03626_),
    .Y(_03946_));
 AO22x1_ASAP7_75t_R _10761_ (.A1(_03945_),
    .A2(_00142_),
    .B1(_00143_),
    .B2(_03946_),
    .Y(_03947_));
 AND2x2_ASAP7_75t_R _10762_ (.A(_03039_),
    .B(_00145_),
    .Y(_03948_));
 AO21x1_ASAP7_75t_R _10763_ (.A1(_03080_),
    .A2(_00144_),
    .B(_03948_),
    .Y(_03949_));
 AO221x1_ASAP7_75t_R _10764_ (.A1(_03597_),
    .A2(_00142_),
    .B1(_03909_),
    .B2(_03949_),
    .C(_03936_),
    .Y(_03950_));
 AO21x1_ASAP7_75t_R _10765_ (.A1(_03068_),
    .A2(_03947_),
    .B(_03950_),
    .Y(_03951_));
 AND2x2_ASAP7_75t_R _10766_ (.A(_03926_),
    .B(_00149_),
    .Y(_03952_));
 AO21x1_ASAP7_75t_R _10767_ (.A1(_03910_),
    .A2(_00148_),
    .B(_03952_),
    .Y(_03953_));
 AND3x1_ASAP7_75t_R _10768_ (.A(_03578_),
    .B(_03860_),
    .C(_00147_),
    .Y(_03954_));
 AO21x1_ASAP7_75t_R _10769_ (.A1(_00146_),
    .A2(_03289_),
    .B(_03954_),
    .Y(_03955_));
 AO221x1_ASAP7_75t_R _10770_ (.A1(_03571_),
    .A2(_03953_),
    .B1(_03955_),
    .B2(_03604_),
    .C(_03695_),
    .Y(_03956_));
 AO21x1_ASAP7_75t_R _10771_ (.A1(_03951_),
    .A2(_03956_),
    .B(_03142_),
    .Y(_03957_));
 OA21x2_ASAP7_75t_R _10772_ (.A1(_03703_),
    .A2(_03944_),
    .B(_03957_),
    .Y(_03958_));
 INVx3_ASAP7_75t_R _10773_ (.A(net14),
    .Y(_03959_));
 OA33x2_ASAP7_75t_R _10774_ (.A1(_03892_),
    .A2(_03917_),
    .A3(_03931_),
    .B1(_03958_),
    .B2(_03959_),
    .B3(_03099_),
    .Y(_03960_));
 INVx1_ASAP7_75t_R _10775_ (.A(net19),
    .Y(_03961_));
 OR3x1_ASAP7_75t_R _10776_ (.A(_03713_),
    .B(_03961_),
    .C(_03715_),
    .Y(_03962_));
 AOI21x1_ASAP7_75t_R _10777_ (.A1(_03712_),
    .A2(_03962_),
    .B(_03718_),
    .Y(_09772_));
 NAND2x1_ASAP7_75t_R _10778_ (.A(_03707_),
    .B(_09772_),
    .Y(_03963_));
 OA21x2_ASAP7_75t_R _10779_ (.A1(_03645_),
    .A2(_03960_),
    .B(_03963_),
    .Y(_03964_));
 XNOR2x2_ASAP7_75t_R _10780_ (.A(_03557_),
    .B(_03964_),
    .Y(_09576_));
 INVx1_ASAP7_75t_R _10781_ (.A(_09576_),
    .Y(_09578_));
 INVx5_ASAP7_75t_R _10782_ (.A(net9),
    .Y(_03965_));
 INVx2_ASAP7_75t_R _10783_ (.A(_00152_),
    .Y(_03966_));
 INVx1_ASAP7_75t_R _10784_ (.A(_00153_),
    .Y(_03967_));
 OA211x2_ASAP7_75t_R _10785_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03837_),
    .C(_03967_),
    .Y(_03968_));
 AOI21x1_ASAP7_75t_R _10786_ (.A1(_03966_),
    .A2(_03847_),
    .B(_03968_),
    .Y(_03969_));
 BUFx10_ASAP7_75t_R _10787_ (.A(_03474_),
    .Y(_03970_));
 AND3x1_ASAP7_75t_R _10788_ (.A(_03019_),
    .B(_03970_),
    .C(_00157_),
    .Y(_03971_));
 AO221x1_ASAP7_75t_R _10789_ (.A1(_03250_),
    .A2(_03736_),
    .B1(_03334_),
    .B2(_00156_),
    .C(_03971_),
    .Y(_03972_));
 OA21x2_ASAP7_75t_R _10790_ (.A1(_03747_),
    .A2(_03969_),
    .B(_03972_),
    .Y(_03973_));
 INVx1_ASAP7_75t_R _10791_ (.A(_00154_),
    .Y(_03974_));
 BUFx12f_ASAP7_75t_R _10792_ (.A(_03435_),
    .Y(_03975_));
 BUFx12f_ASAP7_75t_R _10793_ (.A(_03975_),
    .Y(_03976_));
 INVx1_ASAP7_75t_R _10794_ (.A(_00155_),
    .Y(_03977_));
 AOI22x1_ASAP7_75t_R _10795_ (.A1(_03974_),
    .A2(_03976_),
    .B1(_03409_),
    .B2(_03977_),
    .Y(_03978_));
 BUFx12f_ASAP7_75t_R _10796_ (.A(_03865_),
    .Y(_03979_));
 OA222x2_ASAP7_75t_R _10797_ (.A1(_03098_),
    .A2(_03965_),
    .B1(_03855_),
    .B2(_03973_),
    .C1(_03978_),
    .C2(_03979_),
    .Y(_03980_));
 AND2x2_ASAP7_75t_R _10798_ (.A(_00151_),
    .B(_03467_),
    .Y(_03981_));
 AO21x1_ASAP7_75t_R _10799_ (.A1(_00150_),
    .A2(_03529_),
    .B(_03981_),
    .Y(_03982_));
 AO21x2_ASAP7_75t_R _10800_ (.A1(_03405_),
    .A2(_03982_),
    .B(_03845_),
    .Y(_03983_));
 OA21x2_ASAP7_75t_R _10801_ (.A1(_03345_),
    .A2(_03980_),
    .B(_03983_),
    .Y(_03984_));
 OR3x1_ASAP7_75t_R _10802_ (.A(_03095_),
    .B(_03749_),
    .C(_00161_),
    .Y(_03985_));
 AO21x1_ASAP7_75t_R _10803_ (.A1(_03351_),
    .A2(_03352_),
    .B(_03985_),
    .Y(_03986_));
 OA21x2_ASAP7_75t_R _10804_ (.A1(_00160_),
    .A2(_03348_),
    .B(_03506_),
    .Y(_03987_));
 BUFx12f_ASAP7_75t_R _10805_ (.A(_03338_),
    .Y(_03988_));
 AO21x1_ASAP7_75t_R _10806_ (.A1(_03986_),
    .A2(_03987_),
    .B(_03988_),
    .Y(_03989_));
 AND3x1_ASAP7_75t_R _10807_ (.A(_03860_),
    .B(_03970_),
    .C(_00165_),
    .Y(_03990_));
 AO21x1_ASAP7_75t_R _10808_ (.A1(_00164_),
    .A2(_03975_),
    .B(_03990_),
    .Y(_03991_));
 AO22x1_ASAP7_75t_R _10809_ (.A1(_03209_),
    .A2(_03989_),
    .B1(_03991_),
    .B2(_03747_),
    .Y(_03992_));
 INVx1_ASAP7_75t_R _10810_ (.A(_00163_),
    .Y(_03993_));
 BUFx12_ASAP7_75t_R _10811_ (.A(_03507_),
    .Y(_03994_));
 INVx1_ASAP7_75t_R _10812_ (.A(_00162_),
    .Y(_03995_));
 AOI22x1_ASAP7_75t_R _10813_ (.A1(_03993_),
    .A2(_03994_),
    .B1(_03418_),
    .B2(_03995_),
    .Y(_03996_));
 BUFx12_ASAP7_75t_R _10814_ (.A(_03460_),
    .Y(_03997_));
 OA21x2_ASAP7_75t_R _10815_ (.A1(_03979_),
    .A2(_03996_),
    .B(_03997_),
    .Y(_03998_));
 AND2x2_ASAP7_75t_R _10816_ (.A(_03992_),
    .B(_03998_),
    .Y(_03999_));
 AND2x2_ASAP7_75t_R _10817_ (.A(_00159_),
    .B(_03467_),
    .Y(_04000_));
 AO21x1_ASAP7_75t_R _10818_ (.A1(_00158_),
    .A2(_03529_),
    .B(_04000_),
    .Y(_04001_));
 AND3x4_ASAP7_75t_R _10819_ (.A(_03992_),
    .B(_03998_),
    .C(_04001_),
    .Y(_04002_));
 BUFx16f_ASAP7_75t_R _10820_ (.A(_03862_),
    .Y(_04003_));
 AO211x2_ASAP7_75t_R _10821_ (.A1(_03983_),
    .A2(_03999_),
    .B(_04002_),
    .C(_04003_),
    .Y(_04004_));
 BUFx12f_ASAP7_75t_R _10822_ (.A(_03449_),
    .Y(_04005_));
 AND2x2_ASAP7_75t_R _10823_ (.A(_00134_),
    .B(_04005_),
    .Y(_04006_));
 AO221x2_ASAP7_75t_R _10824_ (.A1(_00135_),
    .A2(_03455_),
    .B1(_03411_),
    .B2(_03521_),
    .C(_04006_),
    .Y(_04007_));
 INVx1_ASAP7_75t_R _10825_ (.A(_00138_),
    .Y(_04008_));
 BUFx6f_ASAP7_75t_R _10826_ (.A(_03031_),
    .Y(_04009_));
 INVx1_ASAP7_75t_R _10827_ (.A(_00139_),
    .Y(_04010_));
 AND3x1_ASAP7_75t_R _10828_ (.A(_04009_),
    .B(_03475_),
    .C(_04010_),
    .Y(_04011_));
 AO22x1_ASAP7_75t_R _10829_ (.A1(_04008_),
    .A2(_03335_),
    .B1(_03759_),
    .B2(_04011_),
    .Y(_04012_));
 AO21x1_ASAP7_75t_R _10830_ (.A1(_03457_),
    .A2(_04012_),
    .B(_03461_),
    .Y(_04013_));
 INVx1_ASAP7_75t_R _10831_ (.A(_00136_),
    .Y(_04014_));
 AND2x2_ASAP7_75t_R _10832_ (.A(_04014_),
    .B(_03334_),
    .Y(_04015_));
 INVx1_ASAP7_75t_R _10833_ (.A(_00137_),
    .Y(_04016_));
 OA211x2_ASAP7_75t_R _10834_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03507_),
    .C(_04016_),
    .Y(_04017_));
 BUFx12f_ASAP7_75t_R _10835_ (.A(_03506_),
    .Y(_04018_));
 OA211x2_ASAP7_75t_R _10836_ (.A1(_04015_),
    .A2(_04017_),
    .B(_03325_),
    .C(_04018_),
    .Y(_04019_));
 BUFx10_ASAP7_75t_R _10837_ (.A(_03736_),
    .Y(_04020_));
 BUFx6f_ASAP7_75t_R _10838_ (.A(_03303_),
    .Y(_04021_));
 BUFx16f_ASAP7_75t_R _10839_ (.A(_04021_),
    .Y(_04022_));
 BUFx12f_ASAP7_75t_R _10840_ (.A(_04022_),
    .Y(_04023_));
 AND2x2_ASAP7_75t_R _10841_ (.A(_00140_),
    .B(_03975_),
    .Y(_04024_));
 AOI221x1_ASAP7_75t_R _10842_ (.A1(_03209_),
    .A2(_04020_),
    .B1(_04023_),
    .B2(_00141_),
    .C(_04024_),
    .Y(_04025_));
 BUFx12_ASAP7_75t_R _10843_ (.A(_03501_),
    .Y(_04026_));
 OA21x2_ASAP7_75t_R _10844_ (.A1(_04019_),
    .A2(_04025_),
    .B(_04026_),
    .Y(_04027_));
 OAI21x1_ASAP7_75t_R _10845_ (.A1(_04013_),
    .A2(_04027_),
    .B(_03412_),
    .Y(_04028_));
 AND2x2_ASAP7_75t_R _10846_ (.A(_00143_),
    .B(_03467_),
    .Y(_04029_));
 AO21x1_ASAP7_75t_R _10847_ (.A1(_00142_),
    .A2(_03432_),
    .B(_04029_),
    .Y(_04030_));
 INVx1_ASAP7_75t_R _10848_ (.A(_00147_),
    .Y(_04031_));
 INVx1_ASAP7_75t_R _10849_ (.A(_00146_),
    .Y(_04032_));
 AOI22x1_ASAP7_75t_R _10850_ (.A1(_04031_),
    .A2(_03428_),
    .B1(_03356_),
    .B2(_04032_),
    .Y(_04033_));
 AND3x1_ASAP7_75t_R _10851_ (.A(_03018_),
    .B(_03301_),
    .C(_00149_),
    .Y(_04034_));
 AO21x1_ASAP7_75t_R _10852_ (.A1(_00148_),
    .A2(_03333_),
    .B(_04034_),
    .Y(_04035_));
 OR2x2_ASAP7_75t_R _10853_ (.A(_03324_),
    .B(_04035_),
    .Y(_04036_));
 AO211x2_ASAP7_75t_R _10854_ (.A1(_03351_),
    .A2(_03352_),
    .B(_03333_),
    .C(_00145_),
    .Y(_04037_));
 OA21x2_ASAP7_75t_R _10855_ (.A1(_00144_),
    .A2(_03312_),
    .B(_03320_),
    .Y(_04038_));
 AO221x1_ASAP7_75t_R _10856_ (.A1(_03359_),
    .A2(_04035_),
    .B1(_04037_),
    .B2(_04038_),
    .C(_03988_),
    .Y(_04039_));
 OA211x2_ASAP7_75t_R _10857_ (.A1(_03979_),
    .A2(_04033_),
    .B(_04036_),
    .C(_04039_),
    .Y(_04040_));
 OA211x2_ASAP7_75t_R _10858_ (.A1(_03845_),
    .A2(_04030_),
    .B(_04040_),
    .C(_03888_),
    .Y(_04041_));
 AO211x2_ASAP7_75t_R _10859_ (.A1(_04007_),
    .A2(_04028_),
    .B(_04041_),
    .C(_03426_),
    .Y(_04042_));
 OAI21x1_ASAP7_75t_R _10860_ (.A1(_03984_),
    .A2(_04004_),
    .B(_04042_),
    .Y(_09575_));
 INVx2_ASAP7_75t_R _10861_ (.A(_09575_),
    .Y(_09577_));
 BUFx12f_ASAP7_75t_R _10862_ (.A(_03142_),
    .Y(_04043_));
 AO22x1_ASAP7_75t_R _10863_ (.A1(_03565_),
    .A2(_00168_),
    .B1(_00169_),
    .B2(_03591_),
    .Y(_04044_));
 AND2x2_ASAP7_75t_R _10864_ (.A(_03807_),
    .B(_00171_),
    .Y(_04045_));
 AO21x1_ASAP7_75t_R _10865_ (.A1(_03061_),
    .A2(_00170_),
    .B(_04045_),
    .Y(_04046_));
 AO21x1_ASAP7_75t_R _10866_ (.A1(_03593_),
    .A2(_04046_),
    .B(_03077_),
    .Y(_04047_));
 AND2x2_ASAP7_75t_R _10867_ (.A(_03597_),
    .B(_00168_),
    .Y(_04048_));
 AO221x1_ASAP7_75t_R _10868_ (.A1(_03589_),
    .A2(_04044_),
    .B1(_04047_),
    .B2(_03021_),
    .C(_04048_),
    .Y(_04049_));
 AND2x2_ASAP7_75t_R _10869_ (.A(_03926_),
    .B(_00175_),
    .Y(_04050_));
 AO21x1_ASAP7_75t_R _10870_ (.A1(_03932_),
    .A2(_00174_),
    .B(_04050_),
    .Y(_04051_));
 AND3x1_ASAP7_75t_R _10871_ (.A(_03578_),
    .B(_03063_),
    .C(_00173_),
    .Y(_04052_));
 AO21x1_ASAP7_75t_R _10872_ (.A1(_00172_),
    .A2(_03577_),
    .B(_04052_),
    .Y(_04053_));
 AO221x1_ASAP7_75t_R _10873_ (.A1(_03571_),
    .A2(_04051_),
    .B1(_04053_),
    .B2(_03604_),
    .C(_03583_),
    .Y(_04054_));
 AND3x2_ASAP7_75t_R _10874_ (.A(_03586_),
    .B(_04049_),
    .C(_04054_),
    .Y(_04055_));
 AND2x2_ASAP7_75t_R _10875_ (.A(_03926_),
    .B(_00183_),
    .Y(_04056_));
 AO21x1_ASAP7_75t_R _10876_ (.A1(_03910_),
    .A2(_00182_),
    .B(_04056_),
    .Y(_04057_));
 AND3x1_ASAP7_75t_R _10877_ (.A(_03091_),
    .B(_03860_),
    .C(_00181_),
    .Y(_04058_));
 AO21x1_ASAP7_75t_R _10878_ (.A1(_00180_),
    .A2(_03289_),
    .B(_04058_),
    .Y(_04059_));
 AO221x1_ASAP7_75t_R _10879_ (.A1(_03571_),
    .A2(_04057_),
    .B1(_04059_),
    .B2(_03604_),
    .C(_03695_),
    .Y(_04060_));
 AO22x1_ASAP7_75t_R _10880_ (.A1(_03945_),
    .A2(_00176_),
    .B1(_00177_),
    .B2(_03946_),
    .Y(_04061_));
 AND2x2_ASAP7_75t_R _10881_ (.A(_03047_),
    .B(_00179_),
    .Y(_04062_));
 AO21x1_ASAP7_75t_R _10882_ (.A1(_03630_),
    .A2(_00178_),
    .B(_04062_),
    .Y(_04063_));
 AO21x1_ASAP7_75t_R _10883_ (.A1(_03087_),
    .A2(_04063_),
    .B(_03077_),
    .Y(_04064_));
 AO21x1_ASAP7_75t_R _10884_ (.A1(_03068_),
    .A2(_04061_),
    .B(_04064_),
    .Y(_04065_));
 AND3x1_ASAP7_75t_R _10885_ (.A(_03173_),
    .B(_04060_),
    .C(_04065_),
    .Y(_04066_));
 NOR3x1_ASAP7_75t_R _10886_ (.A(_04043_),
    .B(_04055_),
    .C(_04066_),
    .Y(_04067_));
 BUFx4f_ASAP7_75t_R _10887_ (.A(_03806_),
    .Y(_04068_));
 AND2x2_ASAP7_75t_R _10888_ (.A(_03065_),
    .B(_00199_),
    .Y(_04069_));
 AO21x1_ASAP7_75t_R _10889_ (.A1(_03138_),
    .A2(_00198_),
    .B(_04069_),
    .Y(_04070_));
 BUFx6f_ASAP7_75t_R _10890_ (.A(_03576_),
    .Y(_04071_));
 AND3x1_ASAP7_75t_R _10891_ (.A(_03058_),
    .B(_04009_),
    .C(_00197_),
    .Y(_04072_));
 AO21x1_ASAP7_75t_R _10892_ (.A1(_00196_),
    .A2(_04071_),
    .B(_04072_),
    .Y(_04073_));
 BUFx6f_ASAP7_75t_R _10893_ (.A(_03581_),
    .Y(_04074_));
 BUFx6f_ASAP7_75t_R _10894_ (.A(_03617_),
    .Y(_04075_));
 AO221x1_ASAP7_75t_R _10895_ (.A1(_04068_),
    .A2(_04070_),
    .B1(_04073_),
    .B2(_04074_),
    .C(_04075_),
    .Y(_04076_));
 BUFx6f_ASAP7_75t_R _10896_ (.A(_03568_),
    .Y(_04077_));
 AND2x2_ASAP7_75t_R _10897_ (.A(_03088_),
    .B(_00194_),
    .Y(_04078_));
 AO21x1_ASAP7_75t_R _10898_ (.A1(_03665_),
    .A2(_00192_),
    .B(_04078_),
    .Y(_04079_));
 BUFx12_ASAP7_75t_R _10899_ (.A(_03945_),
    .Y(_04080_));
 BUFx6f_ASAP7_75t_R _10900_ (.A(_03559_),
    .Y(_04081_));
 BUFx10_ASAP7_75t_R _10901_ (.A(_03650_),
    .Y(_04082_));
 AO21x1_ASAP7_75t_R _10902_ (.A1(_00193_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_04083_));
 AO221x1_ASAP7_75t_R _10903_ (.A1(_00195_),
    .A2(_04077_),
    .B1(_04079_),
    .B2(_04080_),
    .C(_04083_),
    .Y(_04084_));
 BUFx10_ASAP7_75t_R _10904_ (.A(_03585_),
    .Y(_04085_));
 AO21x1_ASAP7_75t_R _10905_ (.A1(_04076_),
    .A2(_04084_),
    .B(_04085_),
    .Y(_04086_));
 BUFx10_ASAP7_75t_R _10906_ (.A(_03057_),
    .Y(_04087_));
 AND2x2_ASAP7_75t_R _10907_ (.A(_04087_),
    .B(_00191_),
    .Y(_04088_));
 AO21x1_ASAP7_75t_R _10908_ (.A1(_03138_),
    .A2(_00190_),
    .B(_04088_),
    .Y(_04089_));
 AND3x1_ASAP7_75t_R _10909_ (.A(_03155_),
    .B(_04009_),
    .C(_00189_),
    .Y(_04090_));
 AO21x1_ASAP7_75t_R _10910_ (.A1(_00188_),
    .A2(_04071_),
    .B(_04090_),
    .Y(_04091_));
 AO221x1_ASAP7_75t_R _10911_ (.A1(_04068_),
    .A2(_04089_),
    .B1(_04091_),
    .B2(_04074_),
    .C(_04075_),
    .Y(_04092_));
 AND2x2_ASAP7_75t_R _10912_ (.A(_03088_),
    .B(_00186_),
    .Y(_04093_));
 AO21x1_ASAP7_75t_R _10913_ (.A1(_03665_),
    .A2(_00184_),
    .B(_04093_),
    .Y(_04094_));
 BUFx10_ASAP7_75t_R _10914_ (.A(_03945_),
    .Y(_04095_));
 AO21x1_ASAP7_75t_R _10915_ (.A1(_00185_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_04096_));
 AO221x1_ASAP7_75t_R _10916_ (.A1(_00187_),
    .A2(_04077_),
    .B1(_04094_),
    .B2(_04095_),
    .C(_04096_),
    .Y(_04097_));
 BUFx6f_ASAP7_75t_R _10917_ (.A(_03173_),
    .Y(_04098_));
 AO21x1_ASAP7_75t_R _10918_ (.A1(_04092_),
    .A2(_04097_),
    .B(_04098_),
    .Y(_04099_));
 BUFx10_ASAP7_75t_R _10919_ (.A(_03154_),
    .Y(_04100_));
 AOI21x1_ASAP7_75t_R _10920_ (.A1(_04086_),
    .A2(_04099_),
    .B(_04100_),
    .Y(_04101_));
 OAI21x1_ASAP7_75t_R _10921_ (.A1(_04067_),
    .A2(_04101_),
    .B(_03705_),
    .Y(_04102_));
 INVx1_ASAP7_75t_R _10922_ (.A(net18),
    .Y(_04103_));
 OR3x1_ASAP7_75t_R _10923_ (.A(_03713_),
    .B(_04103_),
    .C(_03715_),
    .Y(_04104_));
 AOI21x1_ASAP7_75t_R _10924_ (.A1(_03712_),
    .A2(_04104_),
    .B(_03718_),
    .Y(_09770_));
 NAND2x1_ASAP7_75t_R _10925_ (.A(_03707_),
    .B(_09770_),
    .Y(_04105_));
 OA21x2_ASAP7_75t_R _10926_ (.A1(_03645_),
    .A2(_04102_),
    .B(_04105_),
    .Y(_04106_));
 XNOR2x1_ASAP7_75t_R _10927_ (.B(_04106_),
    .Y(_09581_),
    .A(_03557_));
 INVx1_ASAP7_75t_R _10928_ (.A(_09581_),
    .Y(_09583_));
 AO21x2_ASAP7_75t_R _10929_ (.A1(_03233_),
    .A2(_03243_),
    .B(_03865_),
    .Y(_04107_));
 OA22x2_ASAP7_75t_R _10930_ (.A1(_00181_),
    .A2(_03396_),
    .B1(_03511_),
    .B2(_00180_),
    .Y(_04108_));
 OR3x1_ASAP7_75t_R _10931_ (.A(_03095_),
    .B(_03749_),
    .C(_00179_),
    .Y(_04109_));
 OA22x2_ASAP7_75t_R _10932_ (.A1(_00178_),
    .A2(_03312_),
    .B1(_03748_),
    .B2(_04109_),
    .Y(_04110_));
 AND2x2_ASAP7_75t_R _10933_ (.A(_00182_),
    .B(_03332_),
    .Y(_04111_));
 AO221x1_ASAP7_75t_R _10934_ (.A1(_03207_),
    .A2(_03386_),
    .B1(_03312_),
    .B2(_00183_),
    .C(_04111_),
    .Y(_04112_));
 OA21x2_ASAP7_75t_R _10935_ (.A1(_03503_),
    .A2(_04110_),
    .B(_04112_),
    .Y(_04113_));
 AND2x2_ASAP7_75t_R _10936_ (.A(_00177_),
    .B(_03399_),
    .Y(_04114_));
 AO21x1_ASAP7_75t_R _10937_ (.A1(_00176_),
    .A2(_03449_),
    .B(_04114_),
    .Y(_04115_));
 OA22x2_ASAP7_75t_R _10938_ (.A1(_03855_),
    .A2(_04113_),
    .B1(_04115_),
    .B2(_03373_),
    .Y(_04116_));
 OA211x2_ASAP7_75t_R _10939_ (.A1(_04107_),
    .A2(_04108_),
    .B(_04116_),
    .C(_03888_),
    .Y(_04117_));
 NAND2x1_ASAP7_75t_R _10940_ (.A(_00168_),
    .B(_03740_),
    .Y(_04118_));
 NAND2x1_ASAP7_75t_R _10941_ (.A(_00169_),
    .B(_03511_),
    .Y(_04119_));
 OAI22x1_ASAP7_75t_R _10942_ (.A1(_00172_),
    .A2(_03385_),
    .B1(_03414_),
    .B2(_00173_),
    .Y(_04120_));
 AO32x2_ASAP7_75t_R _10943_ (.A1(_03447_),
    .A2(_04118_),
    .A3(_04119_),
    .B1(_03482_),
    .B2(_04120_),
    .Y(_04121_));
 INVx1_ASAP7_75t_R _10944_ (.A(_00171_),
    .Y(_04122_));
 OA211x2_ASAP7_75t_R _10945_ (.A1(_03197_),
    .A2(_03309_),
    .B(_03347_),
    .C(_04122_),
    .Y(_04123_));
 NOR2x1_ASAP7_75t_R _10946_ (.A(_00170_),
    .B(_03304_),
    .Y(_04124_));
 OA211x2_ASAP7_75t_R _10947_ (.A1(_04123_),
    .A2(_04124_),
    .B(_03260_),
    .C(_03320_),
    .Y(_04125_));
 AND2x2_ASAP7_75t_R _10948_ (.A(_00174_),
    .B(_03435_),
    .Y(_04126_));
 AOI221x1_ASAP7_75t_R _10949_ (.A1(_03250_),
    .A2(_03736_),
    .B1(_03305_),
    .B2(_00175_),
    .C(_04126_),
    .Y(_04127_));
 OA21x2_ASAP7_75t_R _10950_ (.A1(_04125_),
    .A2(_04127_),
    .B(_03501_),
    .Y(_04128_));
 OA21x2_ASAP7_75t_R _10951_ (.A1(_03997_),
    .A2(_04128_),
    .B(_03521_),
    .Y(_04129_));
 OAI21x1_ASAP7_75t_R _10952_ (.A1(_04121_),
    .A2(_04129_),
    .B(_03498_),
    .Y(_04130_));
 NAND2x1_ASAP7_75t_R _10953_ (.A(_00184_),
    .B(_03450_),
    .Y(_04131_));
 BUFx12f_ASAP7_75t_R _10954_ (.A(_03408_),
    .Y(_04132_));
 NAND2x1_ASAP7_75t_R _10955_ (.A(_00185_),
    .B(_04132_),
    .Y(_04133_));
 OAI22x1_ASAP7_75t_R _10956_ (.A1(_00188_),
    .A2(_03306_),
    .B1(_03486_),
    .B2(_00189_),
    .Y(_04134_));
 AO32x1_ASAP7_75t_R _10957_ (.A1(_03447_),
    .A2(_04131_),
    .A3(_04133_),
    .B1(_03516_),
    .B2(_04134_),
    .Y(_04135_));
 AND3x1_ASAP7_75t_R _10958_ (.A(_03019_),
    .B(_03970_),
    .C(_00191_),
    .Y(_04136_));
 AOI221x1_ASAP7_75t_R _10959_ (.A1(_03316_),
    .A2(_03321_),
    .B1(_03975_),
    .B2(_00190_),
    .C(_04136_),
    .Y(_04137_));
 INVx1_ASAP7_75t_R _10960_ (.A(_00187_),
    .Y(_04138_));
 OA211x2_ASAP7_75t_R _10961_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03327_),
    .C(_04138_),
    .Y(_04139_));
 NOR2x1_ASAP7_75t_R _10962_ (.A(_00186_),
    .B(_04021_),
    .Y(_04140_));
 OA211x2_ASAP7_75t_R _10963_ (.A1(_04139_),
    .A2(_04140_),
    .B(_03324_),
    .C(_03387_),
    .Y(_04141_));
 OA21x2_ASAP7_75t_R _10964_ (.A1(_04137_),
    .A2(_04141_),
    .B(_03340_),
    .Y(_04142_));
 OA21x2_ASAP7_75t_R _10965_ (.A1(_03997_),
    .A2(_04142_),
    .B(_03521_),
    .Y(_04143_));
 OAI22x1_ASAP7_75t_R _10966_ (.A1(_00197_),
    .A2(_03437_),
    .B1(_04132_),
    .B2(_00196_),
    .Y(_04144_));
 AND3x1_ASAP7_75t_R _10967_ (.A(_03422_),
    .B(_03516_),
    .C(_04144_),
    .Y(_04145_));
 INVx1_ASAP7_75t_R _10968_ (.A(_00195_),
    .Y(_04146_));
 OA211x2_ASAP7_75t_R _10969_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03327_),
    .C(_04146_),
    .Y(_04147_));
 NOR2x1_ASAP7_75t_R _10970_ (.A(_00194_),
    .B(_04021_),
    .Y(_04148_));
 OA211x2_ASAP7_75t_R _10971_ (.A1(_04147_),
    .A2(_04148_),
    .B(_03324_),
    .C(_03387_),
    .Y(_04149_));
 AND2x2_ASAP7_75t_R _10972_ (.A(_00198_),
    .B(_03435_),
    .Y(_04150_));
 AOI221x1_ASAP7_75t_R _10973_ (.A1(_03208_),
    .A2(_03321_),
    .B1(_03313_),
    .B2(_00199_),
    .C(_04150_),
    .Y(_04151_));
 OA21x2_ASAP7_75t_R _10974_ (.A1(_04149_),
    .A2(_04151_),
    .B(_03340_),
    .Y(_04152_));
 BUFx12f_ASAP7_75t_R _10975_ (.A(_03430_),
    .Y(_04153_));
 OA211x2_ASAP7_75t_R _10976_ (.A1(_03225_),
    .A2(_03310_),
    .B(_04021_),
    .C(_00193_),
    .Y(_04154_));
 AOI21x1_ASAP7_75t_R _10977_ (.A1(_00192_),
    .A2(_04153_),
    .B(_04154_),
    .Y(_04155_));
 AO21x1_ASAP7_75t_R _10978_ (.A1(_03420_),
    .A2(_04155_),
    .B(_03550_),
    .Y(_04156_));
 OA21x2_ASAP7_75t_R _10979_ (.A1(_04152_),
    .A2(_04156_),
    .B(_03424_),
    .Y(_04157_));
 OAI22x1_ASAP7_75t_R _10980_ (.A1(_04135_),
    .A2(_04143_),
    .B1(_04145_),
    .B2(_04157_),
    .Y(_04158_));
 OAI21x1_ASAP7_75t_R _10981_ (.A1(_04117_),
    .A2(_04130_),
    .B(_04158_),
    .Y(_09580_));
 INVx2_ASAP7_75t_R _10982_ (.A(_09580_),
    .Y(_09582_));
 BUFx4f_ASAP7_75t_R _10983_ (.A(_03558_),
    .Y(_04159_));
 INVx1_ASAP7_75t_R _10984_ (.A(net17),
    .Y(_04160_));
 OR3x1_ASAP7_75t_R _10985_ (.A(_03713_),
    .B(_04160_),
    .C(_03777_),
    .Y(_04161_));
 AO21x1_ASAP7_75t_R _10986_ (.A1(_03712_),
    .A2(_04161_),
    .B(_03779_),
    .Y(_04162_));
 BUFx6f_ASAP7_75t_R _10987_ (.A(_03127_),
    .Y(_04163_));
 AO22x1_ASAP7_75t_R _10988_ (.A1(_03564_),
    .A2(_00201_),
    .B1(_00202_),
    .B2(_03590_),
    .Y(_04164_));
 AND2x2_ASAP7_75t_R _10989_ (.A(_03038_),
    .B(_00204_),
    .Y(_04165_));
 AO21x1_ASAP7_75t_R _10990_ (.A1(_03054_),
    .A2(_00203_),
    .B(_04165_),
    .Y(_04166_));
 AO21x1_ASAP7_75t_R _10991_ (.A1(_03086_),
    .A2(_04166_),
    .B(_03650_),
    .Y(_04167_));
 AND2x2_ASAP7_75t_R _10992_ (.A(_03096_),
    .B(_00201_),
    .Y(_04168_));
 AO221x1_ASAP7_75t_R _10993_ (.A1(_03027_),
    .A2(_04164_),
    .B1(_04167_),
    .B2(_03149_),
    .C(_04168_),
    .Y(_04169_));
 AND2x2_ASAP7_75t_R _10994_ (.A(_03090_),
    .B(_00208_),
    .Y(_04170_));
 AO21x1_ASAP7_75t_R _10995_ (.A1(_03061_),
    .A2(_00207_),
    .B(_04170_),
    .Y(_04171_));
 AND3x1_ASAP7_75t_R _10996_ (.A(_03807_),
    .B(_03043_),
    .C(_00206_),
    .Y(_04172_));
 AO21x1_ASAP7_75t_R _10997_ (.A1(_00205_),
    .A2(_03576_),
    .B(_04172_),
    .Y(_04173_));
 AO221x1_ASAP7_75t_R _10998_ (.A1(_03806_),
    .A2(_04171_),
    .B1(_04173_),
    .B2(_03581_),
    .C(_03125_),
    .Y(_04174_));
 AND3x1_ASAP7_75t_R _10999_ (.A(_03585_),
    .B(_04169_),
    .C(_04174_),
    .Y(_04175_));
 AND2x2_ASAP7_75t_R _11000_ (.A(_03090_),
    .B(_00216_),
    .Y(_04176_));
 AO21x1_ASAP7_75t_R _11001_ (.A1(_03572_),
    .A2(_00215_),
    .B(_04176_),
    .Y(_04177_));
 AND3x1_ASAP7_75t_R _11002_ (.A(_03807_),
    .B(_03043_),
    .C(_00214_),
    .Y(_04178_));
 AO21x1_ASAP7_75t_R _11003_ (.A1(_00213_),
    .A2(_03576_),
    .B(_04178_),
    .Y(_04179_));
 AO221x1_ASAP7_75t_R _11004_ (.A1(_03806_),
    .A2(_04177_),
    .B1(_04179_),
    .B2(_03581_),
    .C(_03125_),
    .Y(_04180_));
 AO22x1_ASAP7_75t_R _11005_ (.A1(_03055_),
    .A2(_00209_),
    .B1(_00210_),
    .B2(_03626_),
    .Y(_04181_));
 AND2x2_ASAP7_75t_R _11006_ (.A(_03667_),
    .B(_00212_),
    .Y(_04182_));
 AO21x1_ASAP7_75t_R _11007_ (.A1(_03564_),
    .A2(_00211_),
    .B(_04182_),
    .Y(_04183_));
 AO21x1_ASAP7_75t_R _11008_ (.A1(_03088_),
    .A2(_04183_),
    .B(_03610_),
    .Y(_04184_));
 AO21x1_ASAP7_75t_R _11009_ (.A1(_03160_),
    .A2(_04181_),
    .B(_04184_),
    .Y(_04185_));
 AND3x1_ASAP7_75t_R _11010_ (.A(_03173_),
    .B(_04180_),
    .C(_04185_),
    .Y(_04186_));
 AND2x2_ASAP7_75t_R _11011_ (.A(_03038_),
    .B(_00232_),
    .Y(_04187_));
 AO21x1_ASAP7_75t_R _11012_ (.A1(_03054_),
    .A2(_00231_),
    .B(_04187_),
    .Y(_04188_));
 AO21x1_ASAP7_75t_R _11013_ (.A1(_03647_),
    .A2(_04188_),
    .B(_03125_),
    .Y(_04189_));
 AND3x1_ASAP7_75t_R _11014_ (.A(_03807_),
    .B(_03043_),
    .C(_00230_),
    .Y(_04190_));
 OA21x2_ASAP7_75t_R _11015_ (.A1(_03054_),
    .A2(_03103_),
    .B(_00229_),
    .Y(_04191_));
 OA21x2_ASAP7_75t_R _11016_ (.A1(_04190_),
    .A2(_04191_),
    .B(_03121_),
    .Y(_04192_));
 AND2x2_ASAP7_75t_R _11017_ (.A(net12),
    .B(_00227_),
    .Y(_04193_));
 AO21x1_ASAP7_75t_R _11018_ (.A1(_03026_),
    .A2(_00225_),
    .B(_04193_),
    .Y(_04194_));
 AO22x1_ASAP7_75t_R _11019_ (.A1(_00228_),
    .A2(_03567_),
    .B1(_04194_),
    .B2(_03061_),
    .Y(_04195_));
 AO21x1_ASAP7_75t_R _11020_ (.A1(_00226_),
    .A2(_03559_),
    .B(_03650_),
    .Y(_04196_));
 OA22x2_ASAP7_75t_R _11021_ (.A1(_04189_),
    .A2(_04192_),
    .B1(_04195_),
    .B2(_04196_),
    .Y(_04197_));
 AND2x2_ASAP7_75t_R _11022_ (.A(_03038_),
    .B(_00224_),
    .Y(_04198_));
 AO21x1_ASAP7_75t_R _11023_ (.A1(_03054_),
    .A2(_00223_),
    .B(_04198_),
    .Y(_04199_));
 AO21x1_ASAP7_75t_R _11024_ (.A1(_03086_),
    .A2(_04199_),
    .B(_03125_),
    .Y(_04200_));
 AND3x1_ASAP7_75t_R _11025_ (.A(_03667_),
    .B(_03116_),
    .C(_00222_),
    .Y(_04201_));
 OA21x2_ASAP7_75t_R _11026_ (.A1(_03053_),
    .A2(_03095_),
    .B(_00221_),
    .Y(_04202_));
 OA21x2_ASAP7_75t_R _11027_ (.A1(_04201_),
    .A2(_04202_),
    .B(_03121_),
    .Y(_04203_));
 AND2x2_ASAP7_75t_R _11028_ (.A(net12),
    .B(_00219_),
    .Y(_04204_));
 AO21x1_ASAP7_75t_R _11029_ (.A1(_03026_),
    .A2(_00217_),
    .B(_04204_),
    .Y(_04205_));
 AO22x1_ASAP7_75t_R _11030_ (.A1(_00220_),
    .A2(_03567_),
    .B1(_04205_),
    .B2(_03564_),
    .Y(_04206_));
 AO21x1_ASAP7_75t_R _11031_ (.A1(_00218_),
    .A2(_03559_),
    .B(_03650_),
    .Y(_04207_));
 OA222x2_ASAP7_75t_R _11032_ (.A1(_03959_),
    .A2(_03597_),
    .B1(_04200_),
    .B2(_04203_),
    .C1(_04206_),
    .C2(_04207_),
    .Y(_04208_));
 AO211x2_ASAP7_75t_R _11033_ (.A1(_03118_),
    .A2(_04197_),
    .B(_04208_),
    .C(_03032_),
    .Y(_04209_));
 OA31x2_ASAP7_75t_R _11034_ (.A1(_03142_),
    .A2(_04175_),
    .A3(_04186_),
    .B1(_04209_),
    .Y(_04210_));
 OR3x1_ASAP7_75t_R _11035_ (.A(_04163_),
    .B(_03270_),
    .C(_04210_),
    .Y(_04211_));
 OA21x2_ASAP7_75t_R _11036_ (.A1(_04159_),
    .A2(_04162_),
    .B(_04211_),
    .Y(_04212_));
 XNOR2x1_ASAP7_75t_R _11037_ (.B(_04212_),
    .Y(_09586_),
    .A(_03557_));
 INVx1_ASAP7_75t_R _11038_ (.A(_09586_),
    .Y(_09588_));
 AO21x1_ASAP7_75t_R _11039_ (.A1(_03233_),
    .A2(_03243_),
    .B(_03854_),
    .Y(_04213_));
 BUFx12_ASAP7_75t_R _11040_ (.A(_04213_),
    .Y(_04214_));
 OA22x2_ASAP7_75t_R _11041_ (.A1(_00203_),
    .A2(_04021_),
    .B1(_03430_),
    .B2(_00204_),
    .Y(_04215_));
 AND2x2_ASAP7_75t_R _11042_ (.A(_00207_),
    .B(_03332_),
    .Y(_04216_));
 AO221x1_ASAP7_75t_R _11043_ (.A1(_03207_),
    .A2(_03320_),
    .B1(_03304_),
    .B2(_00208_),
    .C(_04216_),
    .Y(_04217_));
 OA21x2_ASAP7_75t_R _11044_ (.A1(_03503_),
    .A2(_04215_),
    .B(_04217_),
    .Y(_04218_));
 NOR2x1_ASAP7_75t_R _11045_ (.A(_04214_),
    .B(_04218_),
    .Y(_04219_));
 NAND2x1_ASAP7_75t_R _11046_ (.A(_00201_),
    .B(_03431_),
    .Y(_04220_));
 NAND2x1_ASAP7_75t_R _11047_ (.A(_00202_),
    .B(_03408_),
    .Y(_04221_));
 OAI22x1_ASAP7_75t_R _11048_ (.A1(_00205_),
    .A2(_04021_),
    .B1(_03430_),
    .B2(_00206_),
    .Y(_04222_));
 AO21x1_ASAP7_75t_R _11049_ (.A1(_03361_),
    .A2(_04222_),
    .B(_03460_),
    .Y(_04223_));
 AO32x1_ASAP7_75t_R _11050_ (.A1(_03447_),
    .A2(_04220_),
    .A3(_04221_),
    .B1(_04223_),
    .B2(_03245_),
    .Y(_04224_));
 OAI22x1_ASAP7_75t_R _11051_ (.A1(_00214_),
    .A2(_03333_),
    .B1(_03399_),
    .B2(_00213_),
    .Y(_04225_));
 OA211x2_ASAP7_75t_R _11052_ (.A1(_03272_),
    .A2(_03286_),
    .B(_03360_),
    .C(_04225_),
    .Y(_04226_));
 OA211x2_ASAP7_75t_R _11053_ (.A1(_03197_),
    .A2(_03309_),
    .B(_03302_),
    .C(_00210_),
    .Y(_04227_));
 AOI21x1_ASAP7_75t_R _11054_ (.A1(_00209_),
    .A2(_03354_),
    .B(_04227_),
    .Y(_04228_));
 INVx1_ASAP7_75t_R _11055_ (.A(_00211_),
    .Y(_04229_));
 INVx1_ASAP7_75t_R _11056_ (.A(_00212_),
    .Y(_04230_));
 OA211x2_ASAP7_75t_R _11057_ (.A1(net24),
    .A2(_03309_),
    .B(_03302_),
    .C(_04230_),
    .Y(_04231_));
 AO221x1_ASAP7_75t_R _11058_ (.A1(_03206_),
    .A2(_03338_),
    .B1(_03332_),
    .B2(_04229_),
    .C(_04231_),
    .Y(_04232_));
 OA211x2_ASAP7_75t_R _11059_ (.A1(_03339_),
    .A2(_04228_),
    .B(_04232_),
    .C(_03393_),
    .Y(_04233_));
 OR3x1_ASAP7_75t_R _11060_ (.A(_03095_),
    .B(_03749_),
    .C(_00216_),
    .Y(_04234_));
 OAI21x1_ASAP7_75t_R _11061_ (.A1(_00215_),
    .A2(_03312_),
    .B(_04234_),
    .Y(_04235_));
 AND3x1_ASAP7_75t_R _11062_ (.A(_03339_),
    .B(_03439_),
    .C(_04235_),
    .Y(_04236_));
 OR4x1_ASAP7_75t_R _11063_ (.A(_03404_),
    .B(_04226_),
    .C(_04233_),
    .D(_04236_),
    .Y(_04237_));
 OA211x2_ASAP7_75t_R _11064_ (.A1(_04219_),
    .A2(_04224_),
    .B(_04237_),
    .C(_03498_),
    .Y(_04238_));
 BUFx3_ASAP7_75t_R _11065_ (.A(_04238_),
    .Y(_04239_));
 NAND2x1_ASAP7_75t_R _11066_ (.A(_00217_),
    .B(_03450_),
    .Y(_04240_));
 NAND2x1_ASAP7_75t_R _11067_ (.A(_00218_),
    .B(_04132_),
    .Y(_04241_));
 OAI22x1_ASAP7_75t_R _11068_ (.A1(_00221_),
    .A2(_03306_),
    .B1(_03450_),
    .B2(_00222_),
    .Y(_04242_));
 AO32x1_ASAP7_75t_R _11069_ (.A1(_03520_),
    .A2(_04240_),
    .A3(_04241_),
    .B1(_03516_),
    .B2(_04242_),
    .Y(_04243_));
 AND3x1_ASAP7_75t_R _11070_ (.A(_03019_),
    .B(_03970_),
    .C(_00224_),
    .Y(_04244_));
 AOI221x1_ASAP7_75t_R _11071_ (.A1(_03208_),
    .A2(_03321_),
    .B1(_03975_),
    .B2(_00223_),
    .C(_04244_),
    .Y(_04245_));
 INVx1_ASAP7_75t_R _11072_ (.A(_00220_),
    .Y(_04246_));
 OA211x2_ASAP7_75t_R _11073_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03347_),
    .C(_04246_),
    .Y(_04247_));
 NOR2x1_ASAP7_75t_R _11074_ (.A(_00219_),
    .B(_04021_),
    .Y(_04248_));
 OA211x2_ASAP7_75t_R _11075_ (.A1(_04247_),
    .A2(_04248_),
    .B(_03324_),
    .C(_03506_),
    .Y(_04249_));
 OA21x2_ASAP7_75t_R _11076_ (.A1(_04245_),
    .A2(_04249_),
    .B(_03501_),
    .Y(_04250_));
 OA21x2_ASAP7_75t_R _11077_ (.A1(_03997_),
    .A2(_04250_),
    .B(_03521_),
    .Y(_04251_));
 OAI22x1_ASAP7_75t_R _11078_ (.A1(_00230_),
    .A2(_03437_),
    .B1(_04132_),
    .B2(_00229_),
    .Y(_04252_));
 AND3x1_ASAP7_75t_R _11079_ (.A(_03539_),
    .B(_03516_),
    .C(_04252_),
    .Y(_04253_));
 INVx1_ASAP7_75t_R _11080_ (.A(_00228_),
    .Y(_04254_));
 OA211x2_ASAP7_75t_R _11081_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03347_),
    .C(_04254_),
    .Y(_04255_));
 NOR2x1_ASAP7_75t_R _11082_ (.A(_00227_),
    .B(_04021_),
    .Y(_04256_));
 OA211x2_ASAP7_75t_R _11083_ (.A1(_04255_),
    .A2(_04256_),
    .B(_03324_),
    .C(_03506_),
    .Y(_04257_));
 AND2x2_ASAP7_75t_R _11084_ (.A(_00231_),
    .B(_03435_),
    .Y(_04258_));
 AOI221x1_ASAP7_75t_R _11085_ (.A1(_03208_),
    .A2(_03321_),
    .B1(_03313_),
    .B2(_00232_),
    .C(_04258_),
    .Y(_04259_));
 OA21x2_ASAP7_75t_R _11086_ (.A1(_04257_),
    .A2(_04259_),
    .B(_03340_),
    .Y(_04260_));
 OA211x2_ASAP7_75t_R _11087_ (.A1(_03225_),
    .A2(_03310_),
    .B(_04021_),
    .C(_00226_),
    .Y(_04261_));
 AOI21x1_ASAP7_75t_R _11088_ (.A1(_00225_),
    .A2(_04153_),
    .B(_04261_),
    .Y(_04262_));
 AO21x1_ASAP7_75t_R _11089_ (.A1(_03420_),
    .A2(_04262_),
    .B(_03550_),
    .Y(_04263_));
 OA21x2_ASAP7_75t_R _11090_ (.A1(_04260_),
    .A2(_04263_),
    .B(_03424_),
    .Y(_04264_));
 OA22x2_ASAP7_75t_R _11091_ (.A1(_04243_),
    .A2(_04251_),
    .B1(_04253_),
    .B2(_04264_),
    .Y(_04265_));
 OR2x2_ASAP7_75t_R _11092_ (.A(_04239_),
    .B(_04265_),
    .Y(_04266_));
 BUFx3_ASAP7_75t_R _11093_ (.A(_04266_),
    .Y(_09585_));
 INVx1_ASAP7_75t_R _11094_ (.A(_09585_),
    .Y(_09587_));
 BUFx6f_ASAP7_75t_R _11095_ (.A(_03807_),
    .Y(_04267_));
 AND2x2_ASAP7_75t_R _11096_ (.A(_04267_),
    .B(_00238_),
    .Y(_04268_));
 AO21x1_ASAP7_75t_R _11097_ (.A1(_03620_),
    .A2(_00237_),
    .B(_04268_),
    .Y(_04269_));
 AO21x1_ASAP7_75t_R _11098_ (.A1(_03074_),
    .A2(_04269_),
    .B(_03623_),
    .Y(_04270_));
 AO22x1_ASAP7_75t_R _11099_ (.A1(_03565_),
    .A2(_00235_),
    .B1(_00236_),
    .B2(_03591_),
    .Y(_04271_));
 AO22x1_ASAP7_75t_R _11100_ (.A1(_03130_),
    .A2(_00235_),
    .B1(_04271_),
    .B2(_03589_),
    .Y(_04272_));
 AO21x1_ASAP7_75t_R _11101_ (.A1(_03201_),
    .A2(_04270_),
    .B(_04272_),
    .Y(_04273_));
 AND2x2_ASAP7_75t_R _11102_ (.A(_03058_),
    .B(_00242_),
    .Y(_04274_));
 AO21x1_ASAP7_75t_R _11103_ (.A1(_03138_),
    .A2(_00241_),
    .B(_04274_),
    .Y(_04275_));
 AND3x1_ASAP7_75t_R _11104_ (.A(_03155_),
    .B(_03020_),
    .C(_00240_),
    .Y(_04276_));
 AO21x1_ASAP7_75t_R _11105_ (.A1(_00239_),
    .A2(_04071_),
    .B(_04276_),
    .Y(_04277_));
 AO221x1_ASAP7_75t_R _11106_ (.A1(_04068_),
    .A2(_04275_),
    .B1(_04277_),
    .B2(_03901_),
    .C(_04075_),
    .Y(_04278_));
 AND3x1_ASAP7_75t_R _11107_ (.A(_04085_),
    .B(_04273_),
    .C(_04278_),
    .Y(_04279_));
 AND2x2_ASAP7_75t_R _11108_ (.A(_04087_),
    .B(_00250_),
    .Y(_04280_));
 AO21x1_ASAP7_75t_R _11109_ (.A1(_03138_),
    .A2(_00249_),
    .B(_04280_),
    .Y(_04281_));
 AND3x1_ASAP7_75t_R _11110_ (.A(_03155_),
    .B(_04009_),
    .C(_00248_),
    .Y(_04282_));
 AO21x1_ASAP7_75t_R _11111_ (.A1(_00247_),
    .A2(_04071_),
    .B(_04282_),
    .Y(_04283_));
 AO221x1_ASAP7_75t_R _11112_ (.A1(_04068_),
    .A2(_04281_),
    .B1(_04283_),
    .B2(_04074_),
    .C(_04075_),
    .Y(_04284_));
 AO22x1_ASAP7_75t_R _11113_ (.A1(_03905_),
    .A2(_00243_),
    .B1(_00244_),
    .B2(_03906_),
    .Y(_04285_));
 AND2x2_ASAP7_75t_R _11114_ (.A(_04267_),
    .B(_00246_),
    .Y(_04286_));
 AO21x1_ASAP7_75t_R _11115_ (.A1(_03620_),
    .A2(_00245_),
    .B(_04286_),
    .Y(_04287_));
 AO21x1_ASAP7_75t_R _11116_ (.A1(_03074_),
    .A2(_04287_),
    .B(_03623_),
    .Y(_04288_));
 AO21x1_ASAP7_75t_R _11117_ (.A1(_03904_),
    .A2(_04285_),
    .B(_04288_),
    .Y(_04289_));
 AND3x1_ASAP7_75t_R _11118_ (.A(_04098_),
    .B(_04284_),
    .C(_04289_),
    .Y(_04290_));
 AND2x2_ASAP7_75t_R _11119_ (.A(_03057_),
    .B(_00266_),
    .Y(_04291_));
 AO21x1_ASAP7_75t_R _11120_ (.A1(_03055_),
    .A2(_00265_),
    .B(_04291_),
    .Y(_04292_));
 AND3x1_ASAP7_75t_R _11121_ (.A(_03047_),
    .B(_03031_),
    .C(_00264_),
    .Y(_04293_));
 AO21x1_ASAP7_75t_R _11122_ (.A1(_00263_),
    .A2(_03123_),
    .B(_04293_),
    .Y(_04294_));
 AO221x1_ASAP7_75t_R _11123_ (.A1(_03109_),
    .A2(_04292_),
    .B1(_04294_),
    .B2(_03635_),
    .C(_03617_),
    .Y(_04295_));
 AND2x2_ASAP7_75t_R _11124_ (.A(_03072_),
    .B(_00261_),
    .Y(_04296_));
 AO21x1_ASAP7_75t_R _11125_ (.A1(_03588_),
    .A2(_00259_),
    .B(_04296_),
    .Y(_04297_));
 AO21x1_ASAP7_75t_R _11126_ (.A1(_00260_),
    .A2(_03560_),
    .B(_03610_),
    .Y(_04298_));
 AO221x1_ASAP7_75t_R _11127_ (.A1(_00262_),
    .A2(_03568_),
    .B1(_04297_),
    .B2(_03062_),
    .C(_04298_),
    .Y(_04299_));
 AND3x1_ASAP7_75t_R _11128_ (.A(_03173_),
    .B(_04295_),
    .C(_04299_),
    .Y(_04300_));
 AND2x2_ASAP7_75t_R _11129_ (.A(_03057_),
    .B(_00258_),
    .Y(_04301_));
 AO21x1_ASAP7_75t_R _11130_ (.A1(_03055_),
    .A2(_00257_),
    .B(_04301_),
    .Y(_04302_));
 AND3x1_ASAP7_75t_R _11131_ (.A(_03047_),
    .B(_03031_),
    .C(_00256_),
    .Y(_04303_));
 AO21x1_ASAP7_75t_R _11132_ (.A1(_00255_),
    .A2(_03123_),
    .B(_04303_),
    .Y(_04304_));
 AO221x1_ASAP7_75t_R _11133_ (.A1(_03109_),
    .A2(_04302_),
    .B1(_04304_),
    .B2(_03635_),
    .C(_03617_),
    .Y(_04305_));
 AND2x2_ASAP7_75t_R _11134_ (.A(_03072_),
    .B(_00253_),
    .Y(_04306_));
 AO21x1_ASAP7_75t_R _11135_ (.A1(_03588_),
    .A2(_00251_),
    .B(_04306_),
    .Y(_04307_));
 AO21x1_ASAP7_75t_R _11136_ (.A1(_00252_),
    .A2(_03560_),
    .B(_03610_),
    .Y(_04308_));
 AO221x1_ASAP7_75t_R _11137_ (.A1(_00254_),
    .A2(_03568_),
    .B1(_04307_),
    .B2(_03062_),
    .C(_04308_),
    .Y(_04309_));
 AND3x1_ASAP7_75t_R _11138_ (.A(_03586_),
    .B(_04305_),
    .C(_04309_),
    .Y(_04310_));
 OR3x1_ASAP7_75t_R _11139_ (.A(_03154_),
    .B(_04300_),
    .C(_04310_),
    .Y(_04311_));
 OA31x2_ASAP7_75t_R _11140_ (.A1(_04043_),
    .A2(_04279_),
    .A3(_04290_),
    .B1(_04311_),
    .Y(_04312_));
 OR2x4_ASAP7_75t_R _11141_ (.A(_03781_),
    .B(_04312_),
    .Y(_04313_));
 INVx1_ASAP7_75t_R _11142_ (.A(net16),
    .Y(_04314_));
 OR3x1_ASAP7_75t_R _11143_ (.A(_03713_),
    .B(_04314_),
    .C(_03715_),
    .Y(_04315_));
 AOI21x1_ASAP7_75t_R _11144_ (.A1(_03712_),
    .A2(_04315_),
    .B(_03718_),
    .Y(_09766_));
 NAND2x1_ASAP7_75t_R _11145_ (.A(_03707_),
    .B(_09766_),
    .Y(_04316_));
 OA21x2_ASAP7_75t_R _11146_ (.A1(_03645_),
    .A2(_04313_),
    .B(_04316_),
    .Y(_04317_));
 XNOR2x1_ASAP7_75t_R _11147_ (.B(_04317_),
    .Y(_09591_),
    .A(_03557_));
 INVx1_ASAP7_75t_R _11148_ (.A(_09591_),
    .Y(_09593_));
 OAI22x1_ASAP7_75t_R _11149_ (.A1(_00258_),
    .A2(_03731_),
    .B1(_03733_),
    .B2(_00254_),
    .Y(_04318_));
 AND3x1_ASAP7_75t_R _11150_ (.A(_00253_),
    .B(_03207_),
    .C(_03386_),
    .Y(_04319_));
 AOI211x1_ASAP7_75t_R _11151_ (.A1(_00257_),
    .A2(_03503_),
    .B(_03328_),
    .C(_04319_),
    .Y(_04320_));
 OA21x2_ASAP7_75t_R _11152_ (.A1(_04318_),
    .A2(_04320_),
    .B(_03443_),
    .Y(_04321_));
 OAI22x1_ASAP7_75t_R _11153_ (.A1(_00255_),
    .A2(_03312_),
    .B1(_03430_),
    .B2(_00256_),
    .Y(_04322_));
 AO21x1_ASAP7_75t_R _11154_ (.A1(_03360_),
    .A2(_04322_),
    .B(_03459_),
    .Y(_04323_));
 AND2x2_ASAP7_75t_R _11155_ (.A(_03244_),
    .B(_04323_),
    .Y(_04324_));
 INVx1_ASAP7_75t_R _11156_ (.A(_00252_),
    .Y(_04325_));
 NAND2x1_ASAP7_75t_R _11157_ (.A(_00251_),
    .B(_03355_),
    .Y(_04326_));
 OA211x2_ASAP7_75t_R _11158_ (.A1(_04325_),
    .A2(_03449_),
    .B(_03446_),
    .C(_04326_),
    .Y(_04327_));
 OAI22x1_ASAP7_75t_R _11159_ (.A1(_00264_),
    .A2(_03395_),
    .B1(_03453_),
    .B2(_00263_),
    .Y(_04328_));
 OR2x2_ASAP7_75t_R _11160_ (.A(_00259_),
    .B(_03398_),
    .Y(_04329_));
 OAI21x1_ASAP7_75t_R _11161_ (.A1(_00260_),
    .A2(_03413_),
    .B(_04329_),
    .Y(_04330_));
 OA211x2_ASAP7_75t_R _11162_ (.A1(_03272_),
    .A2(_03286_),
    .B(_03420_),
    .C(_03422_),
    .Y(_04331_));
 AO32x1_ASAP7_75t_R _11163_ (.A1(_03422_),
    .A2(_03482_),
    .A3(_04328_),
    .B1(_04330_),
    .B2(_04331_),
    .Y(_04332_));
 OAI22x1_ASAP7_75t_R _11164_ (.A1(_00266_),
    .A2(_03731_),
    .B1(_03733_),
    .B2(_00262_),
    .Y(_04333_));
 AND3x1_ASAP7_75t_R _11165_ (.A(_00261_),
    .B(_03207_),
    .C(_03386_),
    .Y(_04334_));
 AOI211x1_ASAP7_75t_R _11166_ (.A1(_00265_),
    .A2(_03503_),
    .B(_03507_),
    .C(_04334_),
    .Y(_04335_));
 OA211x2_ASAP7_75t_R _11167_ (.A1(_04333_),
    .A2(_04335_),
    .B(_03339_),
    .C(_03424_),
    .Y(_04336_));
 AND2x2_ASAP7_75t_R _11168_ (.A(_03424_),
    .B(_03404_),
    .Y(_04337_));
 OA33x2_ASAP7_75t_R _11169_ (.A1(_04321_),
    .A2(_04324_),
    .A3(_04327_),
    .B1(_04332_),
    .B2(_04336_),
    .B3(_04337_),
    .Y(_04338_));
 INVx1_ASAP7_75t_R _11170_ (.A(_00244_),
    .Y(_04339_));
 NAND2x1_ASAP7_75t_R _11171_ (.A(_00243_),
    .B(_03413_),
    .Y(_04340_));
 OA211x2_ASAP7_75t_R _11172_ (.A1(_04339_),
    .A2(_03431_),
    .B(_03446_),
    .C(_04340_),
    .Y(_04341_));
 OAI22x1_ASAP7_75t_R _11173_ (.A1(_00248_),
    .A2(_03465_),
    .B1(_03453_),
    .B2(_00247_),
    .Y(_04342_));
 OA22x2_ASAP7_75t_R _11174_ (.A1(_00245_),
    .A2(_03327_),
    .B1(_03354_),
    .B2(_00246_),
    .Y(_04343_));
 AND2x2_ASAP7_75t_R _11175_ (.A(_00249_),
    .B(_03332_),
    .Y(_04344_));
 AO221x1_ASAP7_75t_R _11176_ (.A1(_03206_),
    .A2(_03319_),
    .B1(_03347_),
    .B2(_00250_),
    .C(_04344_),
    .Y(_04345_));
 OAI21x1_ASAP7_75t_R _11177_ (.A1(_03503_),
    .A2(_04343_),
    .B(_04345_),
    .Y(_04346_));
 AO221x1_ASAP7_75t_R _11178_ (.A1(_03481_),
    .A2(_04342_),
    .B1(_04346_),
    .B2(_03501_),
    .C(_03404_),
    .Y(_04347_));
 OR3x4_ASAP7_75t_R _11179_ (.A(_03276_),
    .B(_03459_),
    .C(_03381_),
    .Y(_04348_));
 OA21x2_ASAP7_75t_R _11180_ (.A1(_03272_),
    .A2(_03286_),
    .B(_04348_),
    .Y(_04349_));
 OAI22x1_ASAP7_75t_R _11181_ (.A1(_00237_),
    .A2(_03347_),
    .B1(_03354_),
    .B2(_00238_),
    .Y(_04350_));
 AND3x1_ASAP7_75t_R _11182_ (.A(_03017_),
    .B(_03301_),
    .C(_00242_),
    .Y(_04351_));
 AOI221x1_ASAP7_75t_R _11183_ (.A1(_03206_),
    .A2(_03319_),
    .B1(_03332_),
    .B2(_00241_),
    .C(_04351_),
    .Y(_04352_));
 AO211x2_ASAP7_75t_R _11184_ (.A1(_03392_),
    .A2(_04350_),
    .B(_04352_),
    .C(_03459_),
    .Y(_04353_));
 INVx1_ASAP7_75t_R _11185_ (.A(_00235_),
    .Y(_01239_));
 NAND2x1_ASAP7_75t_R _11186_ (.A(_00236_),
    .B(_03399_),
    .Y(_04354_));
 OA21x2_ASAP7_75t_R _11187_ (.A1(_01239_),
    .A2(_03399_),
    .B(_04354_),
    .Y(_04355_));
 OAI22x1_ASAP7_75t_R _11188_ (.A1(_00239_),
    .A2(_03347_),
    .B1(_03354_),
    .B2(_00240_),
    .Y(_04356_));
 OA211x2_ASAP7_75t_R _11189_ (.A1(_03272_),
    .A2(_03286_),
    .B(_03360_),
    .C(_04356_),
    .Y(_04357_));
 AO221x1_ASAP7_75t_R _11190_ (.A1(_04349_),
    .A2(_04353_),
    .B1(_04355_),
    .B2(_03446_),
    .C(_04357_),
    .Y(_04358_));
 OA211x2_ASAP7_75t_R _11191_ (.A1(_04341_),
    .A2(_04347_),
    .B(_03498_),
    .C(_04358_),
    .Y(_04359_));
 OR2x2_ASAP7_75t_R _11192_ (.A(_04338_),
    .B(_04359_),
    .Y(_04360_));
 BUFx4f_ASAP7_75t_R _11193_ (.A(_04360_),
    .Y(_09590_));
 INVx2_ASAP7_75t_R _11194_ (.A(_09590_),
    .Y(_09592_));
 BUFx10_ASAP7_75t_R _11195_ (.A(_03626_),
    .Y(_04361_));
 AO22x1_ASAP7_75t_R _11196_ (.A1(_03062_),
    .A2(_00268_),
    .B1(_00269_),
    .B2(_04361_),
    .Y(_04362_));
 AND2x2_ASAP7_75t_R _11197_ (.A(_03675_),
    .B(_00271_),
    .Y(_04363_));
 AO21x2_ASAP7_75t_R _11198_ (.A1(_03111_),
    .A2(_00270_),
    .B(_04363_),
    .Y(_04364_));
 AO21x1_ASAP7_75t_R _11199_ (.A1(_03674_),
    .A2(_04364_),
    .B(_04082_),
    .Y(_04365_));
 AND2x2_ASAP7_75t_R _11200_ (.A(_03097_),
    .B(_00268_),
    .Y(_04366_));
 AO221x1_ASAP7_75t_R _11201_ (.A1(_03068_),
    .A2(_04362_),
    .B1(_04365_),
    .B2(_03215_),
    .C(_04366_),
    .Y(_04367_));
 AND2x2_ASAP7_75t_R _11202_ (.A(_04087_),
    .B(_00275_),
    .Y(_04368_));
 AO21x1_ASAP7_75t_R _11203_ (.A1(_03138_),
    .A2(_00274_),
    .B(_04368_),
    .Y(_04369_));
 AND3x1_ASAP7_75t_R _11204_ (.A(_03058_),
    .B(_04009_),
    .C(_00273_),
    .Y(_04370_));
 AO21x1_ASAP7_75t_R _11205_ (.A1(_00272_),
    .A2(_04071_),
    .B(_04370_),
    .Y(_04371_));
 AO221x1_ASAP7_75t_R _11206_ (.A1(_04068_),
    .A2(_04369_),
    .B1(_04371_),
    .B2(_04074_),
    .C(_04075_),
    .Y(_04372_));
 AND3x1_ASAP7_75t_R _11207_ (.A(_04085_),
    .B(_04367_),
    .C(_04372_),
    .Y(_04373_));
 AND2x2_ASAP7_75t_R _11208_ (.A(_03065_),
    .B(_00283_),
    .Y(_04374_));
 AO21x1_ASAP7_75t_R _11209_ (.A1(_03138_),
    .A2(_00282_),
    .B(_04374_),
    .Y(_04375_));
 BUFx10_ASAP7_75t_R _11210_ (.A(_03576_),
    .Y(_04376_));
 AND3x1_ASAP7_75t_R _11211_ (.A(_03058_),
    .B(_04009_),
    .C(_00281_),
    .Y(_04377_));
 AO21x1_ASAP7_75t_R _11212_ (.A1(_00280_),
    .A2(_04376_),
    .B(_04377_),
    .Y(_04378_));
 BUFx6f_ASAP7_75t_R _11213_ (.A(_03617_),
    .Y(_04379_));
 AO221x1_ASAP7_75t_R _11214_ (.A1(_04068_),
    .A2(_04375_),
    .B1(_04378_),
    .B2(_04074_),
    .C(_04379_),
    .Y(_04380_));
 BUFx10_ASAP7_75t_R _11215_ (.A(_03160_),
    .Y(_04381_));
 AO22x1_ASAP7_75t_R _11216_ (.A1(_03112_),
    .A2(_00276_),
    .B1(_00277_),
    .B2(_04361_),
    .Y(_04382_));
 AND2x2_ASAP7_75t_R _11217_ (.A(_03578_),
    .B(_00279_),
    .Y(_04383_));
 AO21x1_ASAP7_75t_R _11218_ (.A1(_03620_),
    .A2(_00278_),
    .B(_04383_),
    .Y(_04384_));
 AO21x1_ASAP7_75t_R _11219_ (.A1(_03074_),
    .A2(_04384_),
    .B(_03623_),
    .Y(_04385_));
 AO21x1_ASAP7_75t_R _11220_ (.A1(_04381_),
    .A2(_04382_),
    .B(_04385_),
    .Y(_04386_));
 AND3x1_ASAP7_75t_R _11221_ (.A(_04098_),
    .B(_04380_),
    .C(_04386_),
    .Y(_04387_));
 NOR3x1_ASAP7_75t_R _11222_ (.A(_04043_),
    .B(_04373_),
    .C(_04387_),
    .Y(_04388_));
 BUFx6f_ASAP7_75t_R _11223_ (.A(_03674_),
    .Y(_04389_));
 BUFx10_ASAP7_75t_R _11224_ (.A(_03692_),
    .Y(_04390_));
 AND2x2_ASAP7_75t_R _11225_ (.A(_04390_),
    .B(_00299_),
    .Y(_04391_));
 AO21x1_ASAP7_75t_R _11226_ (.A1(_03566_),
    .A2(_00298_),
    .B(_04391_),
    .Y(_04392_));
 BUFx6f_ASAP7_75t_R _11227_ (.A(_03123_),
    .Y(_04393_));
 AND3x1_ASAP7_75t_R _11228_ (.A(_04390_),
    .B(_03149_),
    .C(_00297_),
    .Y(_04394_));
 AO21x1_ASAP7_75t_R _11229_ (.A1(_00296_),
    .A2(_04393_),
    .B(_04394_),
    .Y(_04395_));
 BUFx6f_ASAP7_75t_R _11230_ (.A(_03635_),
    .Y(_04396_));
 BUFx10_ASAP7_75t_R _11231_ (.A(_03636_),
    .Y(_04397_));
 AO221x1_ASAP7_75t_R _11232_ (.A1(_04389_),
    .A2(_04392_),
    .B1(_04395_),
    .B2(_04396_),
    .C(_04397_),
    .Y(_04398_));
 AND2x2_ASAP7_75t_R _11233_ (.A(_03806_),
    .B(_00294_),
    .Y(_04399_));
 AO21x1_ASAP7_75t_R _11234_ (.A1(_03028_),
    .A2(_00292_),
    .B(_04399_),
    .Y(_04400_));
 BUFx12f_ASAP7_75t_R _11235_ (.A(_03112_),
    .Y(_04401_));
 AO21x1_ASAP7_75t_R _11236_ (.A1(_00293_),
    .A2(_03561_),
    .B(_03623_),
    .Y(_04402_));
 AO221x1_ASAP7_75t_R _11237_ (.A1(_00295_),
    .A2(_04077_),
    .B1(_04400_),
    .B2(_04401_),
    .C(_04402_),
    .Y(_04403_));
 BUFx10_ASAP7_75t_R _11238_ (.A(_03585_),
    .Y(_04404_));
 AO21x1_ASAP7_75t_R _11239_ (.A1(_04398_),
    .A2(_04403_),
    .B(_04404_),
    .Y(_04405_));
 AND2x2_ASAP7_75t_R _11240_ (.A(_04390_),
    .B(_00291_),
    .Y(_04406_));
 AO21x1_ASAP7_75t_R _11241_ (.A1(_03566_),
    .A2(_00290_),
    .B(_04406_),
    .Y(_04407_));
 BUFx10_ASAP7_75t_R _11242_ (.A(_03926_),
    .Y(_04408_));
 AND3x1_ASAP7_75t_R _11243_ (.A(_04408_),
    .B(_03149_),
    .C(_00289_),
    .Y(_04409_));
 AO21x1_ASAP7_75t_R _11244_ (.A1(_00288_),
    .A2(_03290_),
    .B(_04409_),
    .Y(_04410_));
 BUFx6f_ASAP7_75t_R _11245_ (.A(_03695_),
    .Y(_04411_));
 AO221x1_ASAP7_75t_R _11246_ (.A1(_04389_),
    .A2(_04407_),
    .B1(_04410_),
    .B2(_04396_),
    .C(_04411_),
    .Y(_04412_));
 BUFx10_ASAP7_75t_R _11247_ (.A(_03568_),
    .Y(_04413_));
 AND2x2_ASAP7_75t_R _11248_ (.A(_03806_),
    .B(_00286_),
    .Y(_04414_));
 AO21x1_ASAP7_75t_R _11249_ (.A1(_03028_),
    .A2(_00284_),
    .B(_04414_),
    .Y(_04415_));
 BUFx10_ASAP7_75t_R _11250_ (.A(_03610_),
    .Y(_04416_));
 AO21x1_ASAP7_75t_R _11251_ (.A1(_00285_),
    .A2(_03561_),
    .B(_04416_),
    .Y(_04417_));
 AO221x1_ASAP7_75t_R _11252_ (.A1(_00287_),
    .A2(_04413_),
    .B1(_04415_),
    .B2(_04401_),
    .C(_04417_),
    .Y(_04418_));
 AO21x1_ASAP7_75t_R _11253_ (.A1(_04412_),
    .A2(_04418_),
    .B(_03174_),
    .Y(_04419_));
 AOI21x1_ASAP7_75t_R _11254_ (.A1(_04405_),
    .A2(_04419_),
    .B(_04100_),
    .Y(_04420_));
 OAI21x1_ASAP7_75t_R _11255_ (.A1(_04388_),
    .A2(_04420_),
    .B(_03705_),
    .Y(_04421_));
 BUFx3_ASAP7_75t_R _11256_ (.A(_03558_),
    .Y(_04422_));
 BUFx6f_ASAP7_75t_R _11257_ (.A(_03703_),
    .Y(_04423_));
 OA21x2_ASAP7_75t_R _11258_ (.A1(_04423_),
    .A2(_03777_),
    .B(_03712_),
    .Y(_04424_));
 OR3x1_ASAP7_75t_R _11259_ (.A(_04422_),
    .B(_03779_),
    .C(_04424_),
    .Y(_04425_));
 OA21x2_ASAP7_75t_R _11260_ (.A1(_03645_),
    .A2(_04421_),
    .B(_04425_),
    .Y(_04426_));
 XNOR2x1_ASAP7_75t_R _11261_ (.B(_04426_),
    .Y(_09596_),
    .A(_03557_));
 INVx1_ASAP7_75t_R _11262_ (.A(_09596_),
    .Y(_09598_));
 OAI22x1_ASAP7_75t_R _11263_ (.A1(_00297_),
    .A2(_03976_),
    .B1(_03409_),
    .B2(_00296_),
    .Y(_04427_));
 AND3x1_ASAP7_75t_R _11264_ (.A(_03539_),
    .B(_03540_),
    .C(_04427_),
    .Y(_04428_));
 INVx1_ASAP7_75t_R _11265_ (.A(_00293_),
    .Y(_04429_));
 NAND2x1_ASAP7_75t_R _11266_ (.A(_00292_),
    .B(_04005_),
    .Y(_04430_));
 OA211x2_ASAP7_75t_R _11267_ (.A1(_04429_),
    .A2(_03357_),
    .B(_04331_),
    .C(_04430_),
    .Y(_04431_));
 BUFx6f_ASAP7_75t_R _11268_ (.A(_03501_),
    .Y(_04432_));
 OAI22x1_ASAP7_75t_R _11269_ (.A1(_00294_),
    .A2(_03428_),
    .B1(_04153_),
    .B2(_00295_),
    .Y(_04433_));
 INVx1_ASAP7_75t_R _11270_ (.A(_00299_),
    .Y(_04434_));
 NOR2x1_ASAP7_75t_R _11271_ (.A(_00298_),
    .B(_03507_),
    .Y(_04435_));
 AO221x1_ASAP7_75t_R _11272_ (.A1(_03250_),
    .A2(_03736_),
    .B1(_03384_),
    .B2(_04434_),
    .C(_04435_),
    .Y(_04436_));
 OA21x2_ASAP7_75t_R _11273_ (.A1(_03747_),
    .A2(_04433_),
    .B(_04436_),
    .Y(_04437_));
 AND3x1_ASAP7_75t_R _11274_ (.A(_04432_),
    .B(_03424_),
    .C(_04437_),
    .Y(_04438_));
 OR4x2_ASAP7_75t_R _11275_ (.A(_04337_),
    .B(_04428_),
    .C(_04431_),
    .D(_04438_),
    .Y(_04439_));
 BUFx12_ASAP7_75t_R _11276_ (.A(_03429_),
    .Y(_04440_));
 BUFx12f_ASAP7_75t_R _11277_ (.A(_03387_),
    .Y(_04441_));
 AND3x1_ASAP7_75t_R _11278_ (.A(_00286_),
    .B(_03251_),
    .C(_04441_),
    .Y(_04442_));
 AO21x1_ASAP7_75t_R _11279_ (.A1(_00290_),
    .A2(_03472_),
    .B(_04442_),
    .Y(_04443_));
 BUFx10_ASAP7_75t_R _11280_ (.A(_03440_),
    .Y(_04444_));
 BUFx6f_ASAP7_75t_R _11281_ (.A(_04153_),
    .Y(_04445_));
 OR3x1_ASAP7_75t_R _11282_ (.A(_00287_),
    .B(_04444_),
    .C(_04445_),
    .Y(_04446_));
 BUFx10_ASAP7_75t_R _11283_ (.A(_03393_),
    .Y(_04447_));
 OR3x1_ASAP7_75t_R _11284_ (.A(_00291_),
    .B(_04447_),
    .C(_03976_),
    .Y(_04448_));
 OA211x2_ASAP7_75t_R _11285_ (.A1(_04440_),
    .A2(_04443_),
    .B(_04446_),
    .C(_04448_),
    .Y(_04449_));
 BUFx6f_ASAP7_75t_R _11286_ (.A(_03845_),
    .Y(_04450_));
 BUFx12_ASAP7_75t_R _11287_ (.A(_03414_),
    .Y(_04451_));
 AND2x2_ASAP7_75t_R _11288_ (.A(_00285_),
    .B(_03454_),
    .Y(_04452_));
 AO21x1_ASAP7_75t_R _11289_ (.A1(_00284_),
    .A2(_04451_),
    .B(_04452_),
    .Y(_04453_));
 OA22x2_ASAP7_75t_R _11290_ (.A1(_00288_),
    .A2(_03385_),
    .B1(_03740_),
    .B2(_00289_),
    .Y(_04454_));
 OA21x2_ASAP7_75t_R _11291_ (.A1(_03979_),
    .A2(_04454_),
    .B(_03299_),
    .Y(_04455_));
 OA22x2_ASAP7_75t_R _11292_ (.A1(_04450_),
    .A2(_04453_),
    .B1(_04455_),
    .B2(_03344_),
    .Y(_04456_));
 OAI21x1_ASAP7_75t_R _11293_ (.A1(_04214_),
    .A2(_04449_),
    .B(_04456_),
    .Y(_04457_));
 BUFx12_ASAP7_75t_R _11294_ (.A(_03836_),
    .Y(_04458_));
 OA22x2_ASAP7_75t_R _11295_ (.A1(_00270_),
    .A2(_03994_),
    .B1(_03765_),
    .B2(_00271_),
    .Y(_04459_));
 BUFx6f_ASAP7_75t_R _11296_ (.A(_03320_),
    .Y(_04460_));
 AND2x2_ASAP7_75t_R _11297_ (.A(_00274_),
    .B(_03465_),
    .Y(_04461_));
 AO221x1_ASAP7_75t_R _11298_ (.A1(_03316_),
    .A2(_04460_),
    .B1(_04022_),
    .B2(_00275_),
    .C(_04461_),
    .Y(_04462_));
 OA211x2_ASAP7_75t_R _11299_ (.A1(_03441_),
    .A2(_04459_),
    .B(_04462_),
    .C(_03550_),
    .Y(_04463_));
 NOR2x1_ASAP7_75t_R _11300_ (.A(_04458_),
    .B(_04463_),
    .Y(_04464_));
 OAI22x1_ASAP7_75t_R _11301_ (.A1(_00272_),
    .A2(_03350_),
    .B1(_03357_),
    .B2(_00273_),
    .Y(_04465_));
 INVx1_ASAP7_75t_R _11302_ (.A(_00268_),
    .Y(_01238_));
 BUFx12f_ASAP7_75t_R _11303_ (.A(_03408_),
    .Y(_04466_));
 NAND2x1_ASAP7_75t_R _11304_ (.A(_00269_),
    .B(_03454_),
    .Y(_04467_));
 OA21x2_ASAP7_75t_R _11305_ (.A1(_01238_),
    .A2(_04466_),
    .B(_04467_),
    .Y(_04468_));
 BUFx10_ASAP7_75t_R _11306_ (.A(_03447_),
    .Y(_04469_));
 AO32x1_ASAP7_75t_R _11307_ (.A1(_03246_),
    .A2(_03362_),
    .A3(_04465_),
    .B1(_04468_),
    .B2(_04469_),
    .Y(_04470_));
 INVx1_ASAP7_75t_R _11308_ (.A(_00277_),
    .Y(_04471_));
 BUFx10_ASAP7_75t_R _11309_ (.A(_03486_),
    .Y(_04472_));
 BUFx12f_ASAP7_75t_R _11310_ (.A(_03356_),
    .Y(_04473_));
 NAND2x1_ASAP7_75t_R _11311_ (.A(_00276_),
    .B(_04473_),
    .Y(_04474_));
 OA211x2_ASAP7_75t_R _11312_ (.A1(_04471_),
    .A2(_04472_),
    .B(_03520_),
    .C(_04474_),
    .Y(_04475_));
 OA22x2_ASAP7_75t_R _11313_ (.A1(_00278_),
    .A2(_03349_),
    .B1(_03418_),
    .B2(_00279_),
    .Y(_04476_));
 AND2x2_ASAP7_75t_R _11314_ (.A(_00282_),
    .B(_03465_),
    .Y(_04477_));
 AO221x1_ASAP7_75t_R _11315_ (.A1(_03316_),
    .A2(_04460_),
    .B1(_04022_),
    .B2(_00283_),
    .C(_04477_),
    .Y(_04478_));
 OAI21x1_ASAP7_75t_R _11316_ (.A1(_04444_),
    .A2(_04476_),
    .B(_04478_),
    .Y(_04479_));
 BUFx10_ASAP7_75t_R _11317_ (.A(_03466_),
    .Y(_04480_));
 OAI22x1_ASAP7_75t_R _11318_ (.A1(_00281_),
    .A2(_04480_),
    .B1(_03541_),
    .B2(_00280_),
    .Y(_04481_));
 AO221x1_ASAP7_75t_R _11319_ (.A1(_04026_),
    .A2(_04479_),
    .B1(_04481_),
    .B2(_03540_),
    .C(_03405_),
    .Y(_04482_));
 OA22x2_ASAP7_75t_R _11320_ (.A1(_04464_),
    .A2(_04470_),
    .B1(_04475_),
    .B2(_04482_),
    .Y(_04483_));
 BUFx6f_ASAP7_75t_R _11321_ (.A(_03499_),
    .Y(_04484_));
 AO22x1_ASAP7_75t_R _11322_ (.A1(_04439_),
    .A2(_04457_),
    .B1(_04483_),
    .B2(_04484_),
    .Y(_04485_));
 BUFx6f_ASAP7_75t_R _11323_ (.A(_04485_),
    .Y(_09595_));
 INVx1_ASAP7_75t_R _11324_ (.A(_09595_),
    .Y(_09597_));
 BUFx6f_ASAP7_75t_R _11325_ (.A(_03143_),
    .Y(_04486_));
 BUFx6f_ASAP7_75t_R _11326_ (.A(_03593_),
    .Y(_04487_));
 BUFx10_ASAP7_75t_R _11327_ (.A(_03807_),
    .Y(_04488_));
 AND2x2_ASAP7_75t_R _11328_ (.A(_04488_),
    .B(_00304_),
    .Y(_04489_));
 AO21x1_ASAP7_75t_R _11329_ (.A1(_03081_),
    .A2(_00303_),
    .B(_04489_),
    .Y(_04490_));
 AO21x1_ASAP7_75t_R _11330_ (.A1(_04487_),
    .A2(_04490_),
    .B(_04416_),
    .Y(_04491_));
 BUFx6f_ASAP7_75t_R _11331_ (.A(_03103_),
    .Y(_04492_));
 BUFx10_ASAP7_75t_R _11332_ (.A(_04492_),
    .Y(_04493_));
 AO22x1_ASAP7_75t_R _11333_ (.A1(_03573_),
    .A2(_00301_),
    .B1(_00302_),
    .B2(_03946_),
    .Y(_04494_));
 AO22x1_ASAP7_75t_R _11334_ (.A1(_04493_),
    .A2(_00301_),
    .B1(_04494_),
    .B2(_03028_),
    .Y(_04495_));
 AO21x1_ASAP7_75t_R _11335_ (.A1(_03201_),
    .A2(_04491_),
    .B(_04495_),
    .Y(_04496_));
 BUFx6f_ASAP7_75t_R _11336_ (.A(_03109_),
    .Y(_04497_));
 BUFx10_ASAP7_75t_R _11337_ (.A(_03630_),
    .Y(_04498_));
 BUFx10_ASAP7_75t_R _11338_ (.A(_03675_),
    .Y(_04499_));
 AND2x2_ASAP7_75t_R _11339_ (.A(_04499_),
    .B(_00308_),
    .Y(_04500_));
 AO21x1_ASAP7_75t_R _11340_ (.A1(_04498_),
    .A2(_00307_),
    .B(_04500_),
    .Y(_04501_));
 BUFx6f_ASAP7_75t_R _11341_ (.A(_03675_),
    .Y(_04502_));
 BUFx10_ASAP7_75t_R _11342_ (.A(_03019_),
    .Y(_04503_));
 AND3x1_ASAP7_75t_R _11343_ (.A(_04502_),
    .B(_04503_),
    .C(_00306_),
    .Y(_04504_));
 AO21x1_ASAP7_75t_R _11344_ (.A1(_00305_),
    .A2(_04393_),
    .B(_04504_),
    .Y(_04505_));
 AO221x1_ASAP7_75t_R _11345_ (.A1(_04497_),
    .A2(_04501_),
    .B1(_04505_),
    .B2(_03922_),
    .C(_04397_),
    .Y(_04506_));
 AND3x1_ASAP7_75t_R _11346_ (.A(_04404_),
    .B(_04496_),
    .C(_04506_),
    .Y(_04507_));
 AND2x2_ASAP7_75t_R _11347_ (.A(_04499_),
    .B(_00316_),
    .Y(_04508_));
 AO21x1_ASAP7_75t_R _11348_ (.A1(_04498_),
    .A2(_00315_),
    .B(_04508_),
    .Y(_04509_));
 AND3x1_ASAP7_75t_R _11349_ (.A(_04502_),
    .B(_04503_),
    .C(_00314_),
    .Y(_04510_));
 AO21x1_ASAP7_75t_R _11350_ (.A1(_00313_),
    .A2(_03897_),
    .B(_04510_),
    .Y(_04511_));
 AO221x1_ASAP7_75t_R _11351_ (.A1(_04497_),
    .A2(_04509_),
    .B1(_04511_),
    .B2(_03922_),
    .C(_03902_),
    .Y(_04512_));
 BUFx10_ASAP7_75t_R _11352_ (.A(_03591_),
    .Y(_04513_));
 AO22x1_ASAP7_75t_R _11353_ (.A1(_03566_),
    .A2(_00309_),
    .B1(_00310_),
    .B2(_04513_),
    .Y(_04514_));
 AND2x2_ASAP7_75t_R _11354_ (.A(_04488_),
    .B(_00312_),
    .Y(_04515_));
 AO21x1_ASAP7_75t_R _11355_ (.A1(_03081_),
    .A2(_00311_),
    .B(_04515_),
    .Y(_04516_));
 AO21x1_ASAP7_75t_R _11356_ (.A1(_04487_),
    .A2(_04516_),
    .B(_04416_),
    .Y(_04517_));
 AO21x1_ASAP7_75t_R _11357_ (.A1(_03029_),
    .A2(_04514_),
    .B(_04517_),
    .Y(_04518_));
 AND3x1_ASAP7_75t_R _11358_ (.A(_04098_),
    .B(_04512_),
    .C(_04518_),
    .Y(_04519_));
 OR3x1_ASAP7_75t_R _11359_ (.A(_04486_),
    .B(_04507_),
    .C(_04519_),
    .Y(_04520_));
 AND2x2_ASAP7_75t_R _11360_ (.A(_04499_),
    .B(_00332_),
    .Y(_04521_));
 AO21x1_ASAP7_75t_R _11361_ (.A1(_04498_),
    .A2(_00331_),
    .B(_04521_),
    .Y(_04522_));
 AND3x1_ASAP7_75t_R _11362_ (.A(_04502_),
    .B(_04503_),
    .C(_00330_),
    .Y(_04523_));
 AO21x1_ASAP7_75t_R _11363_ (.A1(_00329_),
    .A2(_03897_),
    .B(_04523_),
    .Y(_04524_));
 AO221x1_ASAP7_75t_R _11364_ (.A1(_04497_),
    .A2(_04522_),
    .B1(_04524_),
    .B2(_03922_),
    .C(_03902_),
    .Y(_04525_));
 AND2x2_ASAP7_75t_R _11365_ (.A(_03073_),
    .B(_00327_),
    .Y(_04526_));
 AO21x1_ASAP7_75t_R _11366_ (.A1(_03589_),
    .A2(_00325_),
    .B(_04526_),
    .Y(_04527_));
 BUFx10_ASAP7_75t_R _11367_ (.A(_03138_),
    .Y(_04528_));
 BUFx6f_ASAP7_75t_R _11368_ (.A(_03610_),
    .Y(_04529_));
 AO21x1_ASAP7_75t_R _11369_ (.A1(_00326_),
    .A2(_03561_),
    .B(_04529_),
    .Y(_04530_));
 AO221x1_ASAP7_75t_R _11370_ (.A1(_00328_),
    .A2(_04077_),
    .B1(_04527_),
    .B2(_04528_),
    .C(_04530_),
    .Y(_04531_));
 AND3x1_ASAP7_75t_R _11371_ (.A(_03174_),
    .B(_04525_),
    .C(_04531_),
    .Y(_04532_));
 AND2x2_ASAP7_75t_R _11372_ (.A(_04499_),
    .B(_00324_),
    .Y(_04533_));
 AO21x1_ASAP7_75t_R _11373_ (.A1(_04498_),
    .A2(_00323_),
    .B(_04533_),
    .Y(_04534_));
 AND3x1_ASAP7_75t_R _11374_ (.A(_03898_),
    .B(_03473_),
    .C(_00322_),
    .Y(_04535_));
 AO21x1_ASAP7_75t_R _11375_ (.A1(_00321_),
    .A2(_03897_),
    .B(_04535_),
    .Y(_04536_));
 AO221x1_ASAP7_75t_R _11376_ (.A1(_03893_),
    .A2(_04534_),
    .B1(_04536_),
    .B2(_03922_),
    .C(_03902_),
    .Y(_04537_));
 AND2x2_ASAP7_75t_R _11377_ (.A(_03073_),
    .B(_00319_),
    .Y(_04538_));
 AO21x1_ASAP7_75t_R _11378_ (.A1(_03665_),
    .A2(_00317_),
    .B(_04538_),
    .Y(_04539_));
 AO21x1_ASAP7_75t_R _11379_ (.A1(_00318_),
    .A2(_03561_),
    .B(_04529_),
    .Y(_04540_));
 AO221x1_ASAP7_75t_R _11380_ (.A1(_00320_),
    .A2(_04077_),
    .B1(_04539_),
    .B2(_04528_),
    .C(_04540_),
    .Y(_04541_));
 AND3x1_ASAP7_75t_R _11381_ (.A(_04404_),
    .B(_04537_),
    .C(_04541_),
    .Y(_04542_));
 OR3x1_ASAP7_75t_R _11382_ (.A(_04100_),
    .B(_04532_),
    .C(_04542_),
    .Y(_04543_));
 AO21x2_ASAP7_75t_R _11383_ (.A1(_04520_),
    .A2(_04543_),
    .B(_03781_),
    .Y(_04544_));
 BUFx6f_ASAP7_75t_R _11384_ (.A(_04085_),
    .Y(_04545_));
 OA21x2_ASAP7_75t_R _11385_ (.A1(_04545_),
    .A2(_03777_),
    .B(_03712_),
    .Y(_04546_));
 OR3x1_ASAP7_75t_R _11386_ (.A(_04422_),
    .B(_03779_),
    .C(_04546_),
    .Y(_04547_));
 OA21x2_ASAP7_75t_R _11387_ (.A1(_03780_),
    .A2(_04544_),
    .B(_04547_),
    .Y(_04548_));
 XNOR2x2_ASAP7_75t_R _11388_ (.A(_03557_),
    .B(_04548_),
    .Y(_09601_));
 INVx1_ASAP7_75t_R _11389_ (.A(_09601_),
    .Y(_09603_));
 BUFx10_ASAP7_75t_R _11390_ (.A(_03483_),
    .Y(_04549_));
 BUFx12f_ASAP7_75t_R _11391_ (.A(_04480_),
    .Y(_04550_));
 OAI22x1_ASAP7_75t_R _11392_ (.A1(_00314_),
    .A2(_04550_),
    .B1(_03410_),
    .B2(_00313_),
    .Y(_04551_));
 BUFx6f_ASAP7_75t_R _11393_ (.A(_03404_),
    .Y(_04552_));
 OA211x2_ASAP7_75t_R _11394_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03328_),
    .C(_00310_),
    .Y(_04553_));
 AOI21x1_ASAP7_75t_R _11395_ (.A1(_00309_),
    .A2(_03486_),
    .B(_04553_),
    .Y(_04554_));
 INVx1_ASAP7_75t_R _11396_ (.A(_00311_),
    .Y(_04555_));
 INVx1_ASAP7_75t_R _11397_ (.A(_00312_),
    .Y(_04556_));
 OA211x2_ASAP7_75t_R _11398_ (.A1(_03225_),
    .A2(_03310_),
    .B(_03304_),
    .C(_04556_),
    .Y(_04557_));
 AO221x1_ASAP7_75t_R _11399_ (.A1(_03208_),
    .A2(_03988_),
    .B1(_03975_),
    .B2(_04555_),
    .C(_04557_),
    .Y(_04558_));
 OA211x2_ASAP7_75t_R _11400_ (.A1(_03502_),
    .A2(_04554_),
    .B(_04558_),
    .C(_04447_),
    .Y(_04559_));
 BUFx12_ASAP7_75t_R _11401_ (.A(_03384_),
    .Y(_04560_));
 BUFx10_ASAP7_75t_R _11402_ (.A(_03749_),
    .Y(_04561_));
 OR3x1_ASAP7_75t_R _11403_ (.A(_04492_),
    .B(_04561_),
    .C(_00316_),
    .Y(_04562_));
 OAI21x1_ASAP7_75t_R _11404_ (.A1(_00315_),
    .A2(_04560_),
    .B(_04562_),
    .Y(_04563_));
 AND3x1_ASAP7_75t_R _11405_ (.A(_04432_),
    .B(_04444_),
    .C(_04563_),
    .Y(_04564_));
 OR3x1_ASAP7_75t_R _11406_ (.A(_04552_),
    .B(_04559_),
    .C(_04564_),
    .Y(_04565_));
 AO21x2_ASAP7_75t_R _11407_ (.A1(_04549_),
    .A2(_04551_),
    .B(_04565_),
    .Y(_04566_));
 NAND2x1_ASAP7_75t_R _11408_ (.A(_00301_),
    .B(_04451_),
    .Y(_04567_));
 NAND2x1_ASAP7_75t_R _11409_ (.A(_00302_),
    .B(_03479_),
    .Y(_04568_));
 OAI22x1_ASAP7_75t_R _11410_ (.A1(_00305_),
    .A2(_03330_),
    .B1(_03415_),
    .B2(_00306_),
    .Y(_04569_));
 AO32x1_ASAP7_75t_R _11411_ (.A1(_03448_),
    .A2(_04567_),
    .A3(_04568_),
    .B1(_03483_),
    .B2(_04569_),
    .Y(_04570_));
 INVx1_ASAP7_75t_R _11412_ (.A(_00304_),
    .Y(_04571_));
 OA211x2_ASAP7_75t_R _11413_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03837_),
    .C(_04571_),
    .Y(_04572_));
 NOR2x1_ASAP7_75t_R _11414_ (.A(_00303_),
    .B(_03305_),
    .Y(_04573_));
 BUFx6f_ASAP7_75t_R _11415_ (.A(_03260_),
    .Y(_04574_));
 BUFx10_ASAP7_75t_R _11416_ (.A(_03320_),
    .Y(_04575_));
 OA211x2_ASAP7_75t_R _11417_ (.A1(_04572_),
    .A2(_04573_),
    .B(_04574_),
    .C(_04575_),
    .Y(_04576_));
 AND2x2_ASAP7_75t_R _11418_ (.A(_00307_),
    .B(_03436_),
    .Y(_04577_));
 AOI221x1_ASAP7_75t_R _11419_ (.A1(_03251_),
    .A2(_03388_),
    .B1(_03735_),
    .B2(_00308_),
    .C(_04577_),
    .Y(_04578_));
 OA21x2_ASAP7_75t_R _11420_ (.A1(_04576_),
    .A2(_04578_),
    .B(_04432_),
    .Y(_04579_));
 OA21x2_ASAP7_75t_R _11421_ (.A1(_03461_),
    .A2(_04579_),
    .B(_03412_),
    .Y(_04580_));
 OA21x2_ASAP7_75t_R _11422_ (.A1(_04570_),
    .A2(_04580_),
    .B(_03499_),
    .Y(_04581_));
 NAND2x1_ASAP7_75t_R _11423_ (.A(_00317_),
    .B(_03415_),
    .Y(_04582_));
 NAND2x1_ASAP7_75t_R _11424_ (.A(_00318_),
    .B(_03479_),
    .Y(_04583_));
 OAI22x1_ASAP7_75t_R _11425_ (.A1(_00321_),
    .A2(_03330_),
    .B1(_03415_),
    .B2(_00322_),
    .Y(_04584_));
 AO32x1_ASAP7_75t_R _11426_ (.A1(_04469_),
    .A2(_04582_),
    .A3(_04583_),
    .B1(_03483_),
    .B2(_04584_),
    .Y(_04585_));
 BUFx12_ASAP7_75t_R _11427_ (.A(_03474_),
    .Y(_04586_));
 AND3x1_ASAP7_75t_R _11428_ (.A(_04009_),
    .B(_04586_),
    .C(_00324_),
    .Y(_04587_));
 AOI221x1_ASAP7_75t_R _11429_ (.A1(_03251_),
    .A2(_03388_),
    .B1(_03335_),
    .B2(_00323_),
    .C(_04587_),
    .Y(_04588_));
 INVx1_ASAP7_75t_R _11430_ (.A(_00320_),
    .Y(_04589_));
 OA211x2_ASAP7_75t_R _11431_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03837_),
    .C(_04589_),
    .Y(_04590_));
 NOR2x1_ASAP7_75t_R _11432_ (.A(_00319_),
    .B(_03305_),
    .Y(_04591_));
 OA211x2_ASAP7_75t_R _11433_ (.A1(_04590_),
    .A2(_04591_),
    .B(_04574_),
    .C(_04460_),
    .Y(_04592_));
 OA21x2_ASAP7_75t_R _11434_ (.A1(_04588_),
    .A2(_04592_),
    .B(_04432_),
    .Y(_04593_));
 OA21x2_ASAP7_75t_R _11435_ (.A1(_03461_),
    .A2(_04593_),
    .B(_03246_),
    .Y(_04594_));
 OAI22x1_ASAP7_75t_R _11436_ (.A1(_00330_),
    .A2(_03378_),
    .B1(_03479_),
    .B2(_00329_),
    .Y(_04595_));
 AND3x1_ASAP7_75t_R _11437_ (.A(_03539_),
    .B(_03483_),
    .C(_04595_),
    .Y(_04596_));
 INVx1_ASAP7_75t_R _11438_ (.A(_00328_),
    .Y(_04597_));
 OA211x2_ASAP7_75t_R _11439_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03837_),
    .C(_04597_),
    .Y(_04598_));
 NOR2x1_ASAP7_75t_R _11440_ (.A(_00327_),
    .B(_03305_),
    .Y(_04599_));
 OA211x2_ASAP7_75t_R _11441_ (.A1(_04598_),
    .A2(_04599_),
    .B(_04574_),
    .C(_04575_),
    .Y(_04600_));
 AND2x2_ASAP7_75t_R _11442_ (.A(_00331_),
    .B(_03436_),
    .Y(_04601_));
 AOI221x1_ASAP7_75t_R _11443_ (.A1(_03251_),
    .A2(_03388_),
    .B1(_03735_),
    .B2(_00332_),
    .C(_04601_),
    .Y(_04602_));
 OA21x2_ASAP7_75t_R _11444_ (.A1(_04600_),
    .A2(_04602_),
    .B(_04432_),
    .Y(_04603_));
 OA211x2_ASAP7_75t_R _11445_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03305_),
    .C(_00326_),
    .Y(_04604_));
 AOI21x1_ASAP7_75t_R _11446_ (.A1(_00325_),
    .A2(_03722_),
    .B(_04604_),
    .Y(_04605_));
 AO21x1_ASAP7_75t_R _11447_ (.A1(_03484_),
    .A2(_04605_),
    .B(_03299_),
    .Y(_04606_));
 OA21x2_ASAP7_75t_R _11448_ (.A1(_04603_),
    .A2(_04606_),
    .B(_03495_),
    .Y(_04607_));
 OA22x2_ASAP7_75t_R _11449_ (.A1(_04585_),
    .A2(_04594_),
    .B1(_04596_),
    .B2(_04607_),
    .Y(_04608_));
 AO21x1_ASAP7_75t_R _11450_ (.A1(_04566_),
    .A2(_04581_),
    .B(_04608_),
    .Y(_04609_));
 BUFx6f_ASAP7_75t_R _11451_ (.A(_04609_),
    .Y(_09600_));
 INVx1_ASAP7_75t_R _11452_ (.A(_09600_),
    .Y(_09602_));
 BUFx10_ASAP7_75t_R _11453_ (.A(_03556_),
    .Y(_04610_));
 AND2x2_ASAP7_75t_R _11454_ (.A(_04267_),
    .B(_00338_),
    .Y(_04611_));
 AO21x1_ASAP7_75t_R _11455_ (.A1(_03945_),
    .A2(_00337_),
    .B(_04611_),
    .Y(_04612_));
 AO21x1_ASAP7_75t_R _11456_ (.A1(_03074_),
    .A2(_04612_),
    .B(_03623_),
    .Y(_04613_));
 AO22x1_ASAP7_75t_R _11457_ (.A1(_03565_),
    .A2(_00335_),
    .B1(_00336_),
    .B2(_03591_),
    .Y(_04614_));
 AO22x1_ASAP7_75t_R _11458_ (.A1(_04493_),
    .A2(_00335_),
    .B1(_04614_),
    .B2(_03028_),
    .Y(_04615_));
 AO21x1_ASAP7_75t_R _11459_ (.A1(_03201_),
    .A2(_04613_),
    .B(_04615_),
    .Y(_04616_));
 AND2x2_ASAP7_75t_R _11460_ (.A(_03155_),
    .B(_00342_),
    .Y(_04617_));
 AO21x1_ASAP7_75t_R _11461_ (.A1(_03056_),
    .A2(_00341_),
    .B(_04617_),
    .Y(_04618_));
 AND3x1_ASAP7_75t_R _11462_ (.A(_03894_),
    .B(_03020_),
    .C(_00340_),
    .Y(_04619_));
 AO21x1_ASAP7_75t_R _11463_ (.A1(_00339_),
    .A2(_04071_),
    .B(_04619_),
    .Y(_04620_));
 AO221x1_ASAP7_75t_R _11464_ (.A1(_03893_),
    .A2(_04618_),
    .B1(_04620_),
    .B2(_03901_),
    .C(_04075_),
    .Y(_04621_));
 AND3x1_ASAP7_75t_R _11465_ (.A(_04404_),
    .B(_04616_),
    .C(_04621_),
    .Y(_04622_));
 AND2x2_ASAP7_75t_R _11466_ (.A(_03058_),
    .B(_00350_),
    .Y(_04623_));
 AO21x1_ASAP7_75t_R _11467_ (.A1(_03056_),
    .A2(_00349_),
    .B(_04623_),
    .Y(_04624_));
 AND3x1_ASAP7_75t_R _11468_ (.A(_03894_),
    .B(_03020_),
    .C(_00348_),
    .Y(_04625_));
 AO21x1_ASAP7_75t_R _11469_ (.A1(_00347_),
    .A2(_04071_),
    .B(_04625_),
    .Y(_04626_));
 AO221x1_ASAP7_75t_R _11470_ (.A1(_04068_),
    .A2(_04624_),
    .B1(_04626_),
    .B2(_03901_),
    .C(_04075_),
    .Y(_04627_));
 AO22x1_ASAP7_75t_R _11471_ (.A1(_03905_),
    .A2(_00343_),
    .B1(_00344_),
    .B2(_03906_),
    .Y(_04628_));
 AND2x2_ASAP7_75t_R _11472_ (.A(_04267_),
    .B(_00346_),
    .Y(_04629_));
 AO21x1_ASAP7_75t_R _11473_ (.A1(_03945_),
    .A2(_00345_),
    .B(_04629_),
    .Y(_04630_));
 AO21x1_ASAP7_75t_R _11474_ (.A1(_03074_),
    .A2(_04630_),
    .B(_03623_),
    .Y(_04631_));
 AO21x1_ASAP7_75t_R _11475_ (.A1(_03904_),
    .A2(_04628_),
    .B(_04631_),
    .Y(_04632_));
 AND3x1_ASAP7_75t_R _11476_ (.A(_04098_),
    .B(_04627_),
    .C(_04632_),
    .Y(_04633_));
 OR3x1_ASAP7_75t_R _11477_ (.A(_04043_),
    .B(_04622_),
    .C(_04633_),
    .Y(_04634_));
 AND2x2_ASAP7_75t_R _11478_ (.A(_03155_),
    .B(_00366_),
    .Y(_04635_));
 AO21x1_ASAP7_75t_R _11479_ (.A1(_03056_),
    .A2(_00365_),
    .B(_04635_),
    .Y(_04636_));
 AND3x1_ASAP7_75t_R _11480_ (.A(_03894_),
    .B(_03020_),
    .C(_00364_),
    .Y(_04637_));
 AO21x1_ASAP7_75t_R _11481_ (.A1(_00363_),
    .A2(_04071_),
    .B(_04637_),
    .Y(_04638_));
 AO221x1_ASAP7_75t_R _11482_ (.A1(_03893_),
    .A2(_04636_),
    .B1(_04638_),
    .B2(_03901_),
    .C(_04075_),
    .Y(_04639_));
 AND2x2_ASAP7_75t_R _11483_ (.A(_03088_),
    .B(_00361_),
    .Y(_04640_));
 AO21x1_ASAP7_75t_R _11484_ (.A1(_03665_),
    .A2(_00359_),
    .B(_04640_),
    .Y(_04641_));
 AO21x1_ASAP7_75t_R _11485_ (.A1(_00360_),
    .A2(_04081_),
    .B(_04529_),
    .Y(_04642_));
 AO221x1_ASAP7_75t_R _11486_ (.A1(_00362_),
    .A2(_04077_),
    .B1(_04641_),
    .B2(_03082_),
    .C(_04642_),
    .Y(_04643_));
 AND3x1_ASAP7_75t_R _11487_ (.A(_04098_),
    .B(_04639_),
    .C(_04643_),
    .Y(_04644_));
 AND2x2_ASAP7_75t_R _11488_ (.A(_03058_),
    .B(_00358_),
    .Y(_04645_));
 AO21x1_ASAP7_75t_R _11489_ (.A1(_03056_),
    .A2(_00357_),
    .B(_04645_),
    .Y(_04646_));
 AND3x1_ASAP7_75t_R _11490_ (.A(_03155_),
    .B(_03020_),
    .C(_00356_),
    .Y(_04647_));
 AO21x1_ASAP7_75t_R _11491_ (.A1(_00355_),
    .A2(_04071_),
    .B(_04647_),
    .Y(_04648_));
 AO221x1_ASAP7_75t_R _11492_ (.A1(_04068_),
    .A2(_04646_),
    .B1(_04648_),
    .B2(_03901_),
    .C(_04075_),
    .Y(_04649_));
 AND2x2_ASAP7_75t_R _11493_ (.A(_03088_),
    .B(_00353_),
    .Y(_04650_));
 AO21x1_ASAP7_75t_R _11494_ (.A1(_03665_),
    .A2(_00351_),
    .B(_04650_),
    .Y(_04651_));
 AO21x1_ASAP7_75t_R _11495_ (.A1(_00352_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_04652_));
 AO221x1_ASAP7_75t_R _11496_ (.A1(_00354_),
    .A2(_04077_),
    .B1(_04651_),
    .B2(_03082_),
    .C(_04652_),
    .Y(_04653_));
 AND3x1_ASAP7_75t_R _11497_ (.A(_04085_),
    .B(_04649_),
    .C(_04653_),
    .Y(_04654_));
 OR3x1_ASAP7_75t_R _11498_ (.A(_04100_),
    .B(_04644_),
    .C(_04654_),
    .Y(_04655_));
 AO21x2_ASAP7_75t_R _11499_ (.A1(_04634_),
    .A2(_04655_),
    .B(_03781_),
    .Y(_04656_));
 BUFx6f_ASAP7_75t_R _11500_ (.A(_04397_),
    .Y(_04657_));
 OA21x2_ASAP7_75t_R _11501_ (.A1(_04657_),
    .A2(_03777_),
    .B(_03712_),
    .Y(_04658_));
 OR3x1_ASAP7_75t_R _11502_ (.A(_04422_),
    .B(_03718_),
    .C(_04658_),
    .Y(_04659_));
 OA21x2_ASAP7_75t_R _11503_ (.A1(_03780_),
    .A2(_04656_),
    .B(_04659_),
    .Y(_04660_));
 XNOR2x1_ASAP7_75t_R _11504_ (.B(_04660_),
    .Y(_09606_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _11505_ (.A(_09606_),
    .Y(_09608_));
 OAI22x1_ASAP7_75t_R _11506_ (.A1(_00348_),
    .A2(_04550_),
    .B1(_03410_),
    .B2(_00347_),
    .Y(_04661_));
 OA211x2_ASAP7_75t_R _11507_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03328_),
    .C(_00344_),
    .Y(_04662_));
 AOI21x1_ASAP7_75t_R _11508_ (.A1(_00343_),
    .A2(_03740_),
    .B(_04662_),
    .Y(_04663_));
 INVx1_ASAP7_75t_R _11509_ (.A(_00345_),
    .Y(_04664_));
 INVx1_ASAP7_75t_R _11510_ (.A(_00346_),
    .Y(_04665_));
 OA211x2_ASAP7_75t_R _11511_ (.A1(_03225_),
    .A2(_03310_),
    .B(_03304_),
    .C(_04665_),
    .Y(_04666_));
 AO221x1_ASAP7_75t_R _11512_ (.A1(_03208_),
    .A2(_03988_),
    .B1(_03436_),
    .B2(_04664_),
    .C(_04666_),
    .Y(_04667_));
 OA211x2_ASAP7_75t_R _11513_ (.A1(_03502_),
    .A2(_04663_),
    .B(_04667_),
    .C(_03393_),
    .Y(_04668_));
 OR3x1_ASAP7_75t_R _11514_ (.A(_04492_),
    .B(_04561_),
    .C(_00350_),
    .Y(_04669_));
 OAI21x1_ASAP7_75t_R _11515_ (.A1(_00349_),
    .A2(_04560_),
    .B(_04669_),
    .Y(_04670_));
 AND3x1_ASAP7_75t_R _11516_ (.A(_03502_),
    .B(_04444_),
    .C(_04670_),
    .Y(_04671_));
 OR3x1_ASAP7_75t_R _11517_ (.A(_04552_),
    .B(_04668_),
    .C(_04671_),
    .Y(_04672_));
 AO21x2_ASAP7_75t_R _11518_ (.A1(_04549_),
    .A2(_04661_),
    .B(_04672_),
    .Y(_04673_));
 NAND2x1_ASAP7_75t_R _11519_ (.A(_00335_),
    .B(_03415_),
    .Y(_04674_));
 NAND2x1_ASAP7_75t_R _11520_ (.A(_00336_),
    .B(_03401_),
    .Y(_04675_));
 BUFx12f_ASAP7_75t_R _11521_ (.A(_03418_),
    .Y(_04676_));
 OAI22x1_ASAP7_75t_R _11522_ (.A1(_00339_),
    .A2(_03330_),
    .B1(_04676_),
    .B2(_00340_),
    .Y(_04677_));
 AO32x1_ASAP7_75t_R _11523_ (.A1(_04469_),
    .A2(_04674_),
    .A3(_04675_),
    .B1(_03483_),
    .B2(_04677_),
    .Y(_04678_));
 INVx1_ASAP7_75t_R _11524_ (.A(_00338_),
    .Y(_04679_));
 OA211x2_ASAP7_75t_R _11525_ (.A1(_03225_),
    .A2(_03365_),
    .B(_03837_),
    .C(_04679_),
    .Y(_04680_));
 NOR2x1_ASAP7_75t_R _11526_ (.A(_00337_),
    .B(_03305_),
    .Y(_04681_));
 OA211x2_ASAP7_75t_R _11527_ (.A1(_04680_),
    .A2(_04681_),
    .B(_04574_),
    .C(_04460_),
    .Y(_04682_));
 AND2x2_ASAP7_75t_R _11528_ (.A(_00341_),
    .B(_03436_),
    .Y(_04683_));
 AOI221x1_ASAP7_75t_R _11529_ (.A1(_03325_),
    .A2(_04441_),
    .B1(_03385_),
    .B2(_00342_),
    .C(_04683_),
    .Y(_04684_));
 OA21x2_ASAP7_75t_R _11530_ (.A1(_04682_),
    .A2(_04684_),
    .B(_04432_),
    .Y(_04685_));
 OA21x2_ASAP7_75t_R _11531_ (.A1(_03461_),
    .A2(_04685_),
    .B(_03246_),
    .Y(_04686_));
 OA21x2_ASAP7_75t_R _11532_ (.A1(_04678_),
    .A2(_04686_),
    .B(_03499_),
    .Y(_04687_));
 NAND2x1_ASAP7_75t_R _11533_ (.A(_00351_),
    .B(_03415_),
    .Y(_04688_));
 NAND2x1_ASAP7_75t_R _11534_ (.A(_00352_),
    .B(_03401_),
    .Y(_04689_));
 OAI22x1_ASAP7_75t_R _11535_ (.A1(_00355_),
    .A2(_03330_),
    .B1(_04676_),
    .B2(_00356_),
    .Y(_04690_));
 AO32x1_ASAP7_75t_R _11536_ (.A1(_04469_),
    .A2(_04688_),
    .A3(_04689_),
    .B1(_03540_),
    .B2(_04690_),
    .Y(_04691_));
 BUFx6f_ASAP7_75t_R _11537_ (.A(_03031_),
    .Y(_04692_));
 AND3x1_ASAP7_75t_R _11538_ (.A(_04692_),
    .B(_04586_),
    .C(_00358_),
    .Y(_04693_));
 AOI221x1_ASAP7_75t_R _11539_ (.A1(_03251_),
    .A2(_04441_),
    .B1(_03396_),
    .B2(_00357_),
    .C(_04693_),
    .Y(_04694_));
 INVx1_ASAP7_75t_R _11540_ (.A(_00354_),
    .Y(_04695_));
 OA211x2_ASAP7_75t_R _11541_ (.A1(_03225_),
    .A2(_03310_),
    .B(_03837_),
    .C(_04695_),
    .Y(_04696_));
 NOR2x1_ASAP7_75t_R _11542_ (.A(_00353_),
    .B(_03384_),
    .Y(_04697_));
 OA211x2_ASAP7_75t_R _11543_ (.A1(_04696_),
    .A2(_04697_),
    .B(_04574_),
    .C(_04460_),
    .Y(_04698_));
 OA21x2_ASAP7_75t_R _11544_ (.A1(_04694_),
    .A2(_04698_),
    .B(_04432_),
    .Y(_04699_));
 OA21x2_ASAP7_75t_R _11545_ (.A1(_03461_),
    .A2(_04699_),
    .B(_03246_),
    .Y(_04700_));
 OAI22x1_ASAP7_75t_R _11546_ (.A1(_00364_),
    .A2(_03378_),
    .B1(_03401_),
    .B2(_00363_),
    .Y(_04701_));
 AND3x1_ASAP7_75t_R _11547_ (.A(_03539_),
    .B(_03483_),
    .C(_04701_),
    .Y(_04702_));
 INVx1_ASAP7_75t_R _11548_ (.A(_00362_),
    .Y(_04703_));
 OA211x2_ASAP7_75t_R _11549_ (.A1(_03225_),
    .A2(_03310_),
    .B(_03837_),
    .C(_04703_),
    .Y(_04704_));
 NOR2x1_ASAP7_75t_R _11550_ (.A(_00361_),
    .B(_03384_),
    .Y(_04705_));
 OA211x2_ASAP7_75t_R _11551_ (.A1(_04704_),
    .A2(_04705_),
    .B(_04574_),
    .C(_04460_),
    .Y(_04706_));
 AND2x2_ASAP7_75t_R _11552_ (.A(_00365_),
    .B(_03334_),
    .Y(_04707_));
 AOI221x1_ASAP7_75t_R _11553_ (.A1(_03325_),
    .A2(_04441_),
    .B1(_03385_),
    .B2(_00366_),
    .C(_04707_),
    .Y(_04708_));
 OA21x2_ASAP7_75t_R _11554_ (.A1(_04706_),
    .A2(_04708_),
    .B(_04432_),
    .Y(_04709_));
 OA211x2_ASAP7_75t_R _11555_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03384_),
    .C(_00360_),
    .Y(_04710_));
 AOI21x1_ASAP7_75t_R _11556_ (.A1(_00359_),
    .A2(_04005_),
    .B(_04710_),
    .Y(_04711_));
 AO21x1_ASAP7_75t_R _11557_ (.A1(_03484_),
    .A2(_04711_),
    .B(_03299_),
    .Y(_04712_));
 OA21x2_ASAP7_75t_R _11558_ (.A1(_04709_),
    .A2(_04712_),
    .B(_03495_),
    .Y(_04713_));
 OA22x2_ASAP7_75t_R _11559_ (.A1(_04691_),
    .A2(_04700_),
    .B1(_04702_),
    .B2(_04713_),
    .Y(_04714_));
 AO21x1_ASAP7_75t_R _11560_ (.A1(_04673_),
    .A2(_04687_),
    .B(_04714_),
    .Y(_04715_));
 BUFx6f_ASAP7_75t_R _11561_ (.A(_04715_),
    .Y(_09605_));
 INVx1_ASAP7_75t_R _11562_ (.A(_09605_),
    .Y(_09607_));
 AND2x2_ASAP7_75t_R _11563_ (.A(_03926_),
    .B(_00371_),
    .Y(_04716_));
 AO21x1_ASAP7_75t_R _11564_ (.A1(_03910_),
    .A2(_00370_),
    .B(_04716_),
    .Y(_04717_));
 AO21x1_ASAP7_75t_R _11565_ (.A1(_03571_),
    .A2(_04717_),
    .B(_04529_),
    .Y(_04718_));
 AO22x1_ASAP7_75t_R _11566_ (.A1(_03111_),
    .A2(_00368_),
    .B1(_00369_),
    .B2(_03626_),
    .Y(_04719_));
 AO22x1_ASAP7_75t_R _11567_ (.A1(_03130_),
    .A2(_00368_),
    .B1(_04719_),
    .B2(_03665_),
    .Y(_04720_));
 AO21x1_ASAP7_75t_R _11568_ (.A1(_03215_),
    .A2(_04718_),
    .B(_04720_),
    .Y(_04721_));
 BUFx6f_ASAP7_75t_R _11569_ (.A(_03593_),
    .Y(_04722_));
 AND2x2_ASAP7_75t_R _11570_ (.A(_04488_),
    .B(_00375_),
    .Y(_04723_));
 AO21x1_ASAP7_75t_R _11571_ (.A1(_03081_),
    .A2(_00374_),
    .B(_04723_),
    .Y(_04724_));
 AND3x1_ASAP7_75t_R _11572_ (.A(_03065_),
    .B(_03044_),
    .C(_00373_),
    .Y(_04725_));
 AO21x1_ASAP7_75t_R _11573_ (.A1(_00372_),
    .A2(_04376_),
    .B(_04725_),
    .Y(_04726_));
 AO221x1_ASAP7_75t_R _11574_ (.A1(_04722_),
    .A2(_04724_),
    .B1(_04726_),
    .B2(_03582_),
    .C(_03583_),
    .Y(_04727_));
 AND3x1_ASAP7_75t_R _11575_ (.A(_04085_),
    .B(_04721_),
    .C(_04727_),
    .Y(_04728_));
 AND2x2_ASAP7_75t_R _11576_ (.A(_04488_),
    .B(_00383_),
    .Y(_04729_));
 AO21x1_ASAP7_75t_R _11577_ (.A1(_03081_),
    .A2(_00382_),
    .B(_04729_),
    .Y(_04730_));
 AND3x1_ASAP7_75t_R _11578_ (.A(_03040_),
    .B(_03044_),
    .C(_00381_),
    .Y(_04731_));
 AO21x1_ASAP7_75t_R _11579_ (.A1(_00380_),
    .A2(_03577_),
    .B(_04731_),
    .Y(_04732_));
 AO221x1_ASAP7_75t_R _11580_ (.A1(_04722_),
    .A2(_04730_),
    .B1(_04732_),
    .B2(_03582_),
    .C(_03583_),
    .Y(_04733_));
 AO22x1_ASAP7_75t_R _11581_ (.A1(_03056_),
    .A2(_00376_),
    .B1(_00377_),
    .B2(_04361_),
    .Y(_04734_));
 AND2x2_ASAP7_75t_R _11582_ (.A(_03926_),
    .B(_00379_),
    .Y(_04735_));
 AO21x1_ASAP7_75t_R _11583_ (.A1(_03932_),
    .A2(_00378_),
    .B(_04735_),
    .Y(_04736_));
 AO21x1_ASAP7_75t_R _11584_ (.A1(_03571_),
    .A2(_04736_),
    .B(_04529_),
    .Y(_04737_));
 AO21x1_ASAP7_75t_R _11585_ (.A1(_04381_),
    .A2(_04734_),
    .B(_04737_),
    .Y(_04738_));
 AND3x1_ASAP7_75t_R _11586_ (.A(_03119_),
    .B(_04733_),
    .C(_04738_),
    .Y(_04739_));
 OR3x1_ASAP7_75t_R _11587_ (.A(_04043_),
    .B(_04728_),
    .C(_04739_),
    .Y(_04740_));
 AND2x2_ASAP7_75t_R _11588_ (.A(_04488_),
    .B(_00399_),
    .Y(_04741_));
 AO21x1_ASAP7_75t_R _11589_ (.A1(_03081_),
    .A2(_00398_),
    .B(_04741_),
    .Y(_04742_));
 AND3x1_ASAP7_75t_R _11590_ (.A(_03065_),
    .B(_03044_),
    .C(_00397_),
    .Y(_04743_));
 AO21x1_ASAP7_75t_R _11591_ (.A1(_00396_),
    .A2(_03577_),
    .B(_04743_),
    .Y(_04744_));
 AO221x1_ASAP7_75t_R _11592_ (.A1(_04722_),
    .A2(_04742_),
    .B1(_04744_),
    .B2(_03582_),
    .C(_03583_),
    .Y(_04745_));
 AND2x2_ASAP7_75t_R _11593_ (.A(_03647_),
    .B(_00394_),
    .Y(_04746_));
 AO21x1_ASAP7_75t_R _11594_ (.A1(_03160_),
    .A2(_00392_),
    .B(_04746_),
    .Y(_04747_));
 BUFx12f_ASAP7_75t_R _11595_ (.A(_03620_),
    .Y(_04748_));
 AO21x1_ASAP7_75t_R _11596_ (.A1(_00393_),
    .A2(_03560_),
    .B(_03077_),
    .Y(_04749_));
 AO221x1_ASAP7_75t_R _11597_ (.A1(_00395_),
    .A2(_03697_),
    .B1(_04747_),
    .B2(_04748_),
    .C(_04749_),
    .Y(_04750_));
 AND3x1_ASAP7_75t_R _11598_ (.A(_03119_),
    .B(_04745_),
    .C(_04750_),
    .Y(_04751_));
 AND2x2_ASAP7_75t_R _11599_ (.A(_04488_),
    .B(_00391_),
    .Y(_04752_));
 AO21x1_ASAP7_75t_R _11600_ (.A1(_03081_),
    .A2(_00390_),
    .B(_04752_),
    .Y(_04753_));
 AND3x1_ASAP7_75t_R _11601_ (.A(_03040_),
    .B(_03044_),
    .C(_00389_),
    .Y(_04754_));
 AO21x1_ASAP7_75t_R _11602_ (.A1(_00388_),
    .A2(_03577_),
    .B(_04754_),
    .Y(_04755_));
 AO221x1_ASAP7_75t_R _11603_ (.A1(_04722_),
    .A2(_04753_),
    .B1(_04755_),
    .B2(_03582_),
    .C(_03583_),
    .Y(_04756_));
 AND2x2_ASAP7_75t_R _11604_ (.A(_03647_),
    .B(_00386_),
    .Y(_04757_));
 AO21x1_ASAP7_75t_R _11605_ (.A1(_03160_),
    .A2(_00384_),
    .B(_04757_),
    .Y(_04758_));
 AO21x1_ASAP7_75t_R _11606_ (.A1(_00385_),
    .A2(_03560_),
    .B(_03077_),
    .Y(_04759_));
 AO221x2_ASAP7_75t_R _11607_ (.A1(_00387_),
    .A2(_03697_),
    .B1(_04758_),
    .B2(_04748_),
    .C(_04759_),
    .Y(_04760_));
 AND3x1_ASAP7_75t_R _11608_ (.A(_03586_),
    .B(_04756_),
    .C(_04760_),
    .Y(_04761_));
 OR3x1_ASAP7_75t_R _11609_ (.A(_04100_),
    .B(_04751_),
    .C(_04761_),
    .Y(_04762_));
 AO21x2_ASAP7_75t_R _11610_ (.A1(_04740_),
    .A2(_04762_),
    .B(_03781_),
    .Y(_04763_));
 BUFx6f_ASAP7_75t_R _11611_ (.A(_04396_),
    .Y(_04764_));
 OA21x2_ASAP7_75t_R _11612_ (.A1(_04764_),
    .A2(_03777_),
    .B(_03712_),
    .Y(_04765_));
 OR3x1_ASAP7_75t_R _11613_ (.A(_04422_),
    .B(_03718_),
    .C(_04765_),
    .Y(_04766_));
 OA21x2_ASAP7_75t_R _11614_ (.A1(_03780_),
    .A2(_04763_),
    .B(_04766_),
    .Y(_04767_));
 XNOR2x2_ASAP7_75t_R _11615_ (.A(_04610_),
    .B(_04767_),
    .Y(_09611_));
 INVx1_ASAP7_75t_R _11616_ (.A(_09611_),
    .Y(_09613_));
 BUFx12_ASAP7_75t_R _11617_ (.A(_04466_),
    .Y(_04768_));
 AND2x2_ASAP7_75t_R _11618_ (.A(_00368_),
    .B(_04445_),
    .Y(_04769_));
 AO221x1_ASAP7_75t_R _11619_ (.A1(_00369_),
    .A2(_04768_),
    .B1(_03411_),
    .B2(_03246_),
    .C(_04769_),
    .Y(_04770_));
 BUFx12_ASAP7_75t_R _11620_ (.A(_03550_),
    .Y(_04771_));
 NOR2x1_ASAP7_75t_R _11621_ (.A(_00370_),
    .B(_04022_),
    .Y(_04772_));
 INVx1_ASAP7_75t_R _11622_ (.A(_00371_),
    .Y(_04773_));
 OA211x2_ASAP7_75t_R _11623_ (.A1(_03364_),
    .A2(_03490_),
    .B(_03328_),
    .C(_04773_),
    .Y(_04774_));
 OA211x2_ASAP7_75t_R _11624_ (.A1(_04772_),
    .A2(_04774_),
    .B(_03325_),
    .C(_04018_),
    .Y(_04775_));
 AND2x2_ASAP7_75t_R _11625_ (.A(_00374_),
    .B(_03466_),
    .Y(_04776_));
 AOI221x1_ASAP7_75t_R _11626_ (.A1(_03209_),
    .A2(_04020_),
    .B1(_04023_),
    .B2(_00375_),
    .C(_04776_),
    .Y(_04777_));
 OAI21x1_ASAP7_75t_R _11627_ (.A1(_04775_),
    .A2(_04777_),
    .B(_04026_),
    .Y(_04778_));
 NOR2x1_ASAP7_75t_R _11628_ (.A(_00372_),
    .B(_04023_),
    .Y(_04779_));
 INVx1_ASAP7_75t_R _11629_ (.A(_00373_),
    .Y(_04780_));
 AND3x1_ASAP7_75t_R _11630_ (.A(_04780_),
    .B(_03735_),
    .C(_03759_),
    .Y(_04781_));
 OAI21x1_ASAP7_75t_R _11631_ (.A1(_04779_),
    .A2(_04781_),
    .B(_03457_),
    .Y(_04782_));
 BUFx12_ASAP7_75t_R _11632_ (.A(_03243_),
    .Y(_04783_));
 BUFx12_ASAP7_75t_R _11633_ (.A(_03233_),
    .Y(_04784_));
 AO32x2_ASAP7_75t_R _11634_ (.A1(_04771_),
    .A2(_04778_),
    .A3(_04782_),
    .B1(_04783_),
    .B2(_04784_),
    .Y(_04785_));
 BUFx6f_ASAP7_75t_R _11635_ (.A(_03855_),
    .Y(_04786_));
 OA22x2_ASAP7_75t_R _11636_ (.A1(_00378_),
    .A2(_03329_),
    .B1(_03414_),
    .B2(_00379_),
    .Y(_04787_));
 AND2x2_ASAP7_75t_R _11637_ (.A(_00382_),
    .B(_03334_),
    .Y(_04788_));
 AO221x1_ASAP7_75t_R _11638_ (.A1(_03261_),
    .A2(_04018_),
    .B1(_03349_),
    .B2(_00383_),
    .C(_04788_),
    .Y(_04789_));
 OA21x2_ASAP7_75t_R _11639_ (.A1(_03441_),
    .A2(_04787_),
    .B(_04789_),
    .Y(_04790_));
 BUFx10_ASAP7_75t_R _11640_ (.A(_03888_),
    .Y(_04791_));
 OA21x2_ASAP7_75t_R _11641_ (.A1(_04786_),
    .A2(_04790_),
    .B(_04791_),
    .Y(_04792_));
 OA22x2_ASAP7_75t_R _11642_ (.A1(_00381_),
    .A2(_04480_),
    .B1(_03541_),
    .B2(_00380_),
    .Y(_04793_));
 AND2x2_ASAP7_75t_R _11643_ (.A(_00377_),
    .B(_03511_),
    .Y(_04794_));
 AO21x1_ASAP7_75t_R _11644_ (.A1(_00376_),
    .A2(_03383_),
    .B(_04794_),
    .Y(_04795_));
 OA22x2_ASAP7_75t_R _11645_ (.A1(_04107_),
    .A2(_04793_),
    .B1(_04795_),
    .B2(_03845_),
    .Y(_04796_));
 AOI22x1_ASAP7_75t_R _11646_ (.A1(_04770_),
    .A2(_04785_),
    .B1(_04792_),
    .B2(_04796_),
    .Y(_04797_));
 INVx1_ASAP7_75t_R _11647_ (.A(_00385_),
    .Y(_04798_));
 NAND2x1_ASAP7_75t_R _11648_ (.A(_00384_),
    .B(_04445_),
    .Y(_04799_));
 OA211x2_ASAP7_75t_R _11649_ (.A1(_04798_),
    .A2(_04451_),
    .B(_03520_),
    .C(_04799_),
    .Y(_04800_));
 AND3x1_ASAP7_75t_R _11650_ (.A(_03044_),
    .B(_04586_),
    .C(_00391_),
    .Y(_04801_));
 AOI221x1_ASAP7_75t_R _11651_ (.A1(_03325_),
    .A2(_04441_),
    .B1(_03396_),
    .B2(_00390_),
    .C(_04801_),
    .Y(_04802_));
 INVx1_ASAP7_75t_R _11652_ (.A(_00387_),
    .Y(_04803_));
 OA211x2_ASAP7_75t_R _11653_ (.A1(_03225_),
    .A2(_03310_),
    .B(_03304_),
    .C(_04803_),
    .Y(_04804_));
 NOR2x1_ASAP7_75t_R _11654_ (.A(_00386_),
    .B(_03522_),
    .Y(_04805_));
 OA211x2_ASAP7_75t_R _11655_ (.A1(_04804_),
    .A2(_04805_),
    .B(_03316_),
    .C(_03321_),
    .Y(_04806_));
 OA21x2_ASAP7_75t_R _11656_ (.A1(_04802_),
    .A2(_04806_),
    .B(_03502_),
    .Y(_04807_));
 OAI22x1_ASAP7_75t_R _11657_ (.A1(_00388_),
    .A2(_03306_),
    .B1(_03486_),
    .B2(_00389_),
    .Y(_04808_));
 AO21x1_ASAP7_75t_R _11658_ (.A1(_03457_),
    .A2(_04808_),
    .B(_03997_),
    .Y(_04809_));
 OA21x2_ASAP7_75t_R _11659_ (.A1(_04807_),
    .A2(_04809_),
    .B(_03246_),
    .Y(_04810_));
 OAI22x1_ASAP7_75t_R _11660_ (.A1(_00397_),
    .A2(_03397_),
    .B1(_03401_),
    .B2(_00396_),
    .Y(_04811_));
 AND3x1_ASAP7_75t_R _11661_ (.A(_03539_),
    .B(_03540_),
    .C(_04811_),
    .Y(_04812_));
 AND3x1_ASAP7_75t_R _11662_ (.A(_03063_),
    .B(_04586_),
    .C(_00399_),
    .Y(_04813_));
 AOI221x1_ASAP7_75t_R _11663_ (.A1(_03261_),
    .A2(_04018_),
    .B1(_03396_),
    .B2(_00398_),
    .C(_04813_),
    .Y(_04814_));
 INVx1_ASAP7_75t_R _11664_ (.A(_00395_),
    .Y(_04815_));
 OA211x2_ASAP7_75t_R _11665_ (.A1(_03225_),
    .A2(_03310_),
    .B(_03304_),
    .C(_04815_),
    .Y(_04816_));
 NOR2x1_ASAP7_75t_R _11666_ (.A(_00394_),
    .B(_03328_),
    .Y(_04817_));
 OA211x2_ASAP7_75t_R _11667_ (.A1(_04816_),
    .A2(_04817_),
    .B(_03208_),
    .C(_03736_),
    .Y(_04818_));
 OA21x2_ASAP7_75t_R _11668_ (.A1(_04814_),
    .A2(_04818_),
    .B(_03502_),
    .Y(_04819_));
 INVx1_ASAP7_75t_R _11669_ (.A(_00393_),
    .Y(_04820_));
 NAND2x1_ASAP7_75t_R _11670_ (.A(_00392_),
    .B(_03356_),
    .Y(_04821_));
 OA211x2_ASAP7_75t_R _11671_ (.A1(_04820_),
    .A2(_03450_),
    .B(_03420_),
    .C(_04821_),
    .Y(_04822_));
 OA31x2_ASAP7_75t_R _11672_ (.A1(_03405_),
    .A2(_04819_),
    .A3(_04822_),
    .B1(_03495_),
    .Y(_04823_));
 OA22x2_ASAP7_75t_R _11673_ (.A1(_04800_),
    .A2(_04810_),
    .B1(_04812_),
    .B2(_04823_),
    .Y(_04824_));
 AO21x1_ASAP7_75t_R _11674_ (.A1(_03499_),
    .A2(_04797_),
    .B(_04824_),
    .Y(_04825_));
 BUFx6f_ASAP7_75t_R _11675_ (.A(_04825_),
    .Y(_09610_));
 INVx1_ASAP7_75t_R _11676_ (.A(_09610_),
    .Y(_09612_));
 AND2x2_ASAP7_75t_R _11677_ (.A(_04488_),
    .B(_00404_),
    .Y(_04826_));
 AO21x1_ASAP7_75t_R _11678_ (.A1(_03081_),
    .A2(_00403_),
    .B(_04826_),
    .Y(_04827_));
 AO21x1_ASAP7_75t_R _11679_ (.A1(_04487_),
    .A2(_04827_),
    .B(_04416_),
    .Y(_04828_));
 AO22x1_ASAP7_75t_R _11680_ (.A1(_03573_),
    .A2(_00401_),
    .B1(_00402_),
    .B2(_03946_),
    .Y(_04829_));
 AO22x1_ASAP7_75t_R _11681_ (.A1(_04493_),
    .A2(_00401_),
    .B1(_04829_),
    .B2(_03132_),
    .Y(_04830_));
 AO21x1_ASAP7_75t_R _11682_ (.A1(_03022_),
    .A2(_04828_),
    .B(_04830_),
    .Y(_04831_));
 AND2x2_ASAP7_75t_R _11683_ (.A(_04499_),
    .B(_00408_),
    .Y(_04832_));
 AO21x1_ASAP7_75t_R _11684_ (.A1(_04498_),
    .A2(_00407_),
    .B(_04832_),
    .Y(_04833_));
 AND3x1_ASAP7_75t_R _11685_ (.A(_04502_),
    .B(_04503_),
    .C(_00406_),
    .Y(_04834_));
 AO21x1_ASAP7_75t_R _11686_ (.A1(_00405_),
    .A2(_04393_),
    .B(_04834_),
    .Y(_04835_));
 AO221x1_ASAP7_75t_R _11687_ (.A1(_04497_),
    .A2(_04833_),
    .B1(_04835_),
    .B2(_03922_),
    .C(_04397_),
    .Y(_04836_));
 AND3x1_ASAP7_75t_R _11688_ (.A(_04404_),
    .B(_04831_),
    .C(_04836_),
    .Y(_04837_));
 AND2x2_ASAP7_75t_R _11689_ (.A(_04499_),
    .B(_00416_),
    .Y(_04838_));
 AO21x1_ASAP7_75t_R _11690_ (.A1(_04498_),
    .A2(_00415_),
    .B(_04838_),
    .Y(_04839_));
 AND3x1_ASAP7_75t_R _11691_ (.A(_04502_),
    .B(_04503_),
    .C(_00414_),
    .Y(_04840_));
 AO21x1_ASAP7_75t_R _11692_ (.A1(_00413_),
    .A2(_03897_),
    .B(_04840_),
    .Y(_04841_));
 AO221x1_ASAP7_75t_R _11693_ (.A1(_04497_),
    .A2(_04839_),
    .B1(_04841_),
    .B2(_03922_),
    .C(_03902_),
    .Y(_04842_));
 AO22x1_ASAP7_75t_R _11694_ (.A1(_03566_),
    .A2(_00409_),
    .B1(_00410_),
    .B2(_04513_),
    .Y(_04843_));
 AND2x2_ASAP7_75t_R _11695_ (.A(_04488_),
    .B(_00412_),
    .Y(_04844_));
 AO21x1_ASAP7_75t_R _11696_ (.A1(_03081_),
    .A2(_00411_),
    .B(_04844_),
    .Y(_04845_));
 AO21x1_ASAP7_75t_R _11697_ (.A1(_04487_),
    .A2(_04845_),
    .B(_04416_),
    .Y(_04846_));
 AO21x1_ASAP7_75t_R _11698_ (.A1(_03029_),
    .A2(_04843_),
    .B(_04846_),
    .Y(_04847_));
 AND3x1_ASAP7_75t_R _11699_ (.A(_04098_),
    .B(_04842_),
    .C(_04847_),
    .Y(_04848_));
 OR3x1_ASAP7_75t_R _11700_ (.A(_04486_),
    .B(_04837_),
    .C(_04848_),
    .Y(_04849_));
 BUFx6f_ASAP7_75t_R _11701_ (.A(_03689_),
    .Y(_04850_));
 BUFx4f_ASAP7_75t_R _11702_ (.A(_03910_),
    .Y(_04851_));
 AND2x2_ASAP7_75t_R _11703_ (.A(_04408_),
    .B(_00432_),
    .Y(_04852_));
 AO21x1_ASAP7_75t_R _11704_ (.A1(_04851_),
    .A2(_00431_),
    .B(_04852_),
    .Y(_04853_));
 AND3x1_ASAP7_75t_R _11705_ (.A(_04408_),
    .B(_03064_),
    .C(_00430_),
    .Y(_04854_));
 AO21x1_ASAP7_75t_R _11706_ (.A1(_00429_),
    .A2(_03290_),
    .B(_04854_),
    .Y(_04855_));
 BUFx6f_ASAP7_75t_R _11707_ (.A(_03604_),
    .Y(_04856_));
 AO221x1_ASAP7_75t_R _11708_ (.A1(_04850_),
    .A2(_04853_),
    .B1(_04855_),
    .B2(_04856_),
    .C(_04411_),
    .Y(_04857_));
 AND2x2_ASAP7_75t_R _11709_ (.A(_03593_),
    .B(_00427_),
    .Y(_04858_));
 AO21x1_ASAP7_75t_R _11710_ (.A1(_03068_),
    .A2(_00425_),
    .B(_04858_),
    .Y(_04859_));
 BUFx6f_ASAP7_75t_R _11711_ (.A(_03905_),
    .Y(_04860_));
 BUFx10_ASAP7_75t_R _11712_ (.A(_03560_),
    .Y(_04861_));
 BUFx10_ASAP7_75t_R _11713_ (.A(_03077_),
    .Y(_04862_));
 AO21x1_ASAP7_75t_R _11714_ (.A1(_00426_),
    .A2(_04861_),
    .B(_04862_),
    .Y(_04863_));
 AO221x1_ASAP7_75t_R _11715_ (.A1(_00428_),
    .A2(_04413_),
    .B1(_04859_),
    .B2(_04860_),
    .C(_04863_),
    .Y(_04864_));
 AO21x1_ASAP7_75t_R _11716_ (.A1(_04857_),
    .A2(_04864_),
    .B(_04404_),
    .Y(_04865_));
 AND2x2_ASAP7_75t_R _11717_ (.A(_04408_),
    .B(_00424_),
    .Y(_04866_));
 AO21x1_ASAP7_75t_R _11718_ (.A1(_04851_),
    .A2(_00423_),
    .B(_04866_),
    .Y(_04867_));
 AND3x1_ASAP7_75t_R _11719_ (.A(_04408_),
    .B(_03064_),
    .C(_00422_),
    .Y(_04868_));
 AO21x1_ASAP7_75t_R _11720_ (.A1(_00421_),
    .A2(_03290_),
    .B(_04868_),
    .Y(_04869_));
 AO221x1_ASAP7_75t_R _11721_ (.A1(_04850_),
    .A2(_04867_),
    .B1(_04869_),
    .B2(_04396_),
    .C(_04411_),
    .Y(_04870_));
 AND2x2_ASAP7_75t_R _11722_ (.A(_03593_),
    .B(_00419_),
    .Y(_04871_));
 AO21x1_ASAP7_75t_R _11723_ (.A1(_03068_),
    .A2(_00417_),
    .B(_04871_),
    .Y(_04872_));
 AO21x1_ASAP7_75t_R _11724_ (.A1(_00418_),
    .A2(_03561_),
    .B(_04862_),
    .Y(_04873_));
 AO221x1_ASAP7_75t_R _11725_ (.A1(_00420_),
    .A2(_04413_),
    .B1(_04872_),
    .B2(_04860_),
    .C(_04873_),
    .Y(_04874_));
 AO21x1_ASAP7_75t_R _11726_ (.A1(_04870_),
    .A2(_04874_),
    .B(_03174_),
    .Y(_04875_));
 AO21x1_ASAP7_75t_R _11727_ (.A1(_04865_),
    .A2(_04875_),
    .B(_04100_),
    .Y(_04876_));
 AO21x2_ASAP7_75t_R _11728_ (.A1(_04849_),
    .A2(_04876_),
    .B(_03781_),
    .Y(_04877_));
 OA21x2_ASAP7_75t_R _11729_ (.A1(_03291_),
    .A2(_03777_),
    .B(_03711_),
    .Y(_04878_));
 OR3x1_ASAP7_75t_R _11730_ (.A(_04422_),
    .B(_03718_),
    .C(_04878_),
    .Y(_04879_));
 OA21x2_ASAP7_75t_R _11731_ (.A1(_03780_),
    .A2(_04877_),
    .B(_04879_),
    .Y(_04880_));
 XNOR2x1_ASAP7_75t_R _11732_ (.B(_04880_),
    .Y(_09616_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _11733_ (.A(_09616_),
    .Y(_09618_));
 BUFx6f_ASAP7_75t_R _11734_ (.A(_03520_),
    .Y(_04881_));
 BUFx12_ASAP7_75t_R _11735_ (.A(_03455_),
    .Y(_04882_));
 OR2x2_ASAP7_75t_R _11736_ (.A(_00410_),
    .B(_04451_),
    .Y(_04883_));
 OAI21x1_ASAP7_75t_R _11737_ (.A1(_00409_),
    .A2(_04882_),
    .B(_04883_),
    .Y(_04884_));
 BUFx12_ASAP7_75t_R _11738_ (.A(_03504_),
    .Y(_04885_));
 OA22x2_ASAP7_75t_R _11739_ (.A1(_00411_),
    .A2(_04560_),
    .B1(_03450_),
    .B2(_00412_),
    .Y(_04886_));
 AND2x2_ASAP7_75t_R _11740_ (.A(_00415_),
    .B(_03436_),
    .Y(_04887_));
 AO221x1_ASAP7_75t_R _11741_ (.A1(_03325_),
    .A2(_04441_),
    .B1(_03385_),
    .B2(_00416_),
    .C(_04887_),
    .Y(_04888_));
 OAI21x1_ASAP7_75t_R _11742_ (.A1(_04885_),
    .A2(_04886_),
    .B(_04888_),
    .Y(_04889_));
 OAI22x1_ASAP7_75t_R _11743_ (.A1(_00414_),
    .A2(_03377_),
    .B1(_03455_),
    .B2(_00413_),
    .Y(_04890_));
 BUFx6f_ASAP7_75t_R _11744_ (.A(_03516_),
    .Y(_04891_));
 AO221x1_ASAP7_75t_R _11745_ (.A1(_03341_),
    .A2(_04889_),
    .B1(_04890_),
    .B2(_04891_),
    .C(_04552_),
    .Y(_04892_));
 AO21x1_ASAP7_75t_R _11746_ (.A1(_04881_),
    .A2(_04884_),
    .B(_04892_),
    .Y(_04893_));
 NAND2x1_ASAP7_75t_R _11747_ (.A(_00401_),
    .B(_04472_),
    .Y(_04894_));
 NAND2x1_ASAP7_75t_R _11748_ (.A(_00402_),
    .B(_03455_),
    .Y(_04895_));
 BUFx6f_ASAP7_75t_R _11749_ (.A(_03329_),
    .Y(_04896_));
 OAI22x1_ASAP7_75t_R _11750_ (.A1(_00405_),
    .A2(_04896_),
    .B1(_04472_),
    .B2(_00406_),
    .Y(_04897_));
 AO32x1_ASAP7_75t_R _11751_ (.A1(_03448_),
    .A2(_04894_),
    .A3(_04895_),
    .B1(_04891_),
    .B2(_04897_),
    .Y(_04898_));
 BUFx6f_ASAP7_75t_R _11752_ (.A(_03997_),
    .Y(_04899_));
 NOR2x1_ASAP7_75t_R _11753_ (.A(_00403_),
    .B(_03313_),
    .Y(_04900_));
 INVx1_ASAP7_75t_R _11754_ (.A(_00404_),
    .Y(_04901_));
 OA211x2_ASAP7_75t_R _11755_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03507_),
    .C(_04901_),
    .Y(_04902_));
 OA211x2_ASAP7_75t_R _11756_ (.A1(_04900_),
    .A2(_04902_),
    .B(_03325_),
    .C(_04018_),
    .Y(_04903_));
 AND2x2_ASAP7_75t_R _11757_ (.A(_00407_),
    .B(_03975_),
    .Y(_04904_));
 AOI221x1_ASAP7_75t_R _11758_ (.A1(_03209_),
    .A2(_04020_),
    .B1(_04560_),
    .B2(_00408_),
    .C(_04904_),
    .Y(_04905_));
 OA21x2_ASAP7_75t_R _11759_ (.A1(_04903_),
    .A2(_04905_),
    .B(_04026_),
    .Y(_04906_));
 OA21x2_ASAP7_75t_R _11760_ (.A1(_04899_),
    .A2(_04906_),
    .B(_03412_),
    .Y(_04907_));
 OA21x2_ASAP7_75t_R _11761_ (.A1(_04898_),
    .A2(_04907_),
    .B(_03499_),
    .Y(_04908_));
 OAI22x1_ASAP7_75t_R _11762_ (.A1(_00430_),
    .A2(_03377_),
    .B1(_03455_),
    .B2(_00429_),
    .Y(_04909_));
 AND2x2_ASAP7_75t_R _11763_ (.A(_04891_),
    .B(_04909_),
    .Y(_04910_));
 OR3x1_ASAP7_75t_R _11764_ (.A(_03096_),
    .B(_03749_),
    .C(_00428_),
    .Y(_04911_));
 OA22x2_ASAP7_75t_R _11765_ (.A1(_00427_),
    .A2(_03329_),
    .B1(_03748_),
    .B2(_04911_),
    .Y(_04912_));
 AND3x1_ASAP7_75t_R _11766_ (.A(_03044_),
    .B(_04586_),
    .C(_00432_),
    .Y(_04913_));
 AO221x1_ASAP7_75t_R _11767_ (.A1(_03261_),
    .A2(_04575_),
    .B1(_03847_),
    .B2(_00431_),
    .C(_04913_),
    .Y(_04914_));
 OAI21x1_ASAP7_75t_R _11768_ (.A1(_03472_),
    .A2(_04912_),
    .B(_04914_),
    .Y(_04915_));
 OR2x2_ASAP7_75t_R _11769_ (.A(_00425_),
    .B(_03400_),
    .Y(_04916_));
 OAI21x1_ASAP7_75t_R _11770_ (.A1(_00426_),
    .A2(_04676_),
    .B(_04916_),
    .Y(_04917_));
 AO221x1_ASAP7_75t_R _11771_ (.A1(_03341_),
    .A2(_04915_),
    .B1(_04917_),
    .B2(_04469_),
    .C(_04552_),
    .Y(_04918_));
 OA22x2_ASAP7_75t_R _11772_ (.A1(_00419_),
    .A2(_03994_),
    .B1(_03765_),
    .B2(_00420_),
    .Y(_04919_));
 AND2x2_ASAP7_75t_R _11773_ (.A(_00423_),
    .B(_03395_),
    .Y(_04920_));
 AO221x1_ASAP7_75t_R _11774_ (.A1(_04574_),
    .A2(_04575_),
    .B1(_03428_),
    .B2(_00424_),
    .C(_04920_),
    .Y(_04921_));
 OAI21x1_ASAP7_75t_R _11775_ (.A1(_03441_),
    .A2(_04919_),
    .B(_04921_),
    .Y(_04922_));
 OR2x2_ASAP7_75t_R _11776_ (.A(_00417_),
    .B(_03467_),
    .Y(_04923_));
 OAI21x1_ASAP7_75t_R _11777_ (.A1(_00418_),
    .A2(_03383_),
    .B(_04923_),
    .Y(_04924_));
 OAI22x1_ASAP7_75t_R _11778_ (.A1(_00421_),
    .A2(_03306_),
    .B1(_03486_),
    .B2(_00422_),
    .Y(_04925_));
 AO21x1_ASAP7_75t_R _11779_ (.A1(_03457_),
    .A2(_04925_),
    .B(_03997_),
    .Y(_04926_));
 AO221x1_ASAP7_75t_R _11780_ (.A1(_04026_),
    .A2(_04922_),
    .B1(_04924_),
    .B2(_04469_),
    .C(_04926_),
    .Y(_04927_));
 OA211x2_ASAP7_75t_R _11781_ (.A1(_04910_),
    .A2(_04918_),
    .B(_04927_),
    .C(_03495_),
    .Y(_04928_));
 AO21x1_ASAP7_75t_R _11782_ (.A1(_04893_),
    .A2(_04908_),
    .B(_04928_),
    .Y(_04929_));
 BUFx6f_ASAP7_75t_R _11783_ (.A(_04929_),
    .Y(_09615_));
 INVx1_ASAP7_75t_R _11784_ (.A(_09615_),
    .Y(_09617_));
 AND2x2_ASAP7_75t_R _11785_ (.A(_03894_),
    .B(_00457_),
    .Y(_04930_));
 AO21x1_ASAP7_75t_R _11786_ (.A1(_03685_),
    .A2(_00456_),
    .B(_04930_),
    .Y(_04931_));
 AND3x1_ASAP7_75t_R _11787_ (.A(_03898_),
    .B(_03473_),
    .C(_00455_),
    .Y(_04932_));
 AO21x1_ASAP7_75t_R _11788_ (.A1(_00454_),
    .A2(_03897_),
    .B(_04932_),
    .Y(_04933_));
 AO221x1_ASAP7_75t_R _11789_ (.A1(_03893_),
    .A2(_04931_),
    .B1(_04933_),
    .B2(_03901_),
    .C(_03902_),
    .Y(_04934_));
 AO22x1_ASAP7_75t_R _11790_ (.A1(_03905_),
    .A2(_00450_),
    .B1(_00451_),
    .B2(_03906_),
    .Y(_04935_));
 AND2x2_ASAP7_75t_R _11791_ (.A(_03692_),
    .B(_00453_),
    .Y(_04936_));
 AO21x1_ASAP7_75t_R _11792_ (.A1(_03910_),
    .A2(_00452_),
    .B(_04936_),
    .Y(_04937_));
 AO221x1_ASAP7_75t_R _11793_ (.A1(_03097_),
    .A2(_00450_),
    .B1(_03909_),
    .B2(_04937_),
    .C(_03914_),
    .Y(_04938_));
 AO21x1_ASAP7_75t_R _11794_ (.A1(_03904_),
    .A2(_04935_),
    .B(_04938_),
    .Y(_04939_));
 AND3x1_ASAP7_75t_R _11795_ (.A(_03143_),
    .B(_04934_),
    .C(_04939_),
    .Y(_04940_));
 AND2x2_ASAP7_75t_R _11796_ (.A(_03894_),
    .B(_00441_),
    .Y(_04941_));
 AO21x1_ASAP7_75t_R _11797_ (.A1(_03685_),
    .A2(_00440_),
    .B(_04941_),
    .Y(_04942_));
 AND3x1_ASAP7_75t_R _11798_ (.A(_04499_),
    .B(_03020_),
    .C(_00439_),
    .Y(_04943_));
 AO21x1_ASAP7_75t_R _11799_ (.A1(_00438_),
    .A2(_04071_),
    .B(_04943_),
    .Y(_04944_));
 AO221x1_ASAP7_75t_R _11800_ (.A1(_03893_),
    .A2(_04942_),
    .B1(_04944_),
    .B2(_03901_),
    .C(_04075_),
    .Y(_04945_));
 AO22x1_ASAP7_75t_R _11801_ (.A1(_03905_),
    .A2(_00434_),
    .B1(_00435_),
    .B2(_03906_),
    .Y(_04946_));
 AND2x2_ASAP7_75t_R _11802_ (.A(_03692_),
    .B(_00437_),
    .Y(_04947_));
 AO21x1_ASAP7_75t_R _11803_ (.A1(_03565_),
    .A2(_00436_),
    .B(_04947_),
    .Y(_04948_));
 AO221x1_ASAP7_75t_R _11804_ (.A1(_03097_),
    .A2(_00434_),
    .B1(_03909_),
    .B2(_04948_),
    .C(_03914_),
    .Y(_04949_));
 AO21x1_ASAP7_75t_R _11805_ (.A1(_03904_),
    .A2(_04946_),
    .B(_04949_),
    .Y(_04950_));
 AND3x1_ASAP7_75t_R _11806_ (.A(_03703_),
    .B(_04945_),
    .C(_04950_),
    .Y(_04951_));
 OR3x1_ASAP7_75t_R _11807_ (.A(_03127_),
    .B(_04940_),
    .C(_04951_),
    .Y(_04952_));
 AO22x1_ASAP7_75t_R _11808_ (.A1(_04851_),
    .A2(_00458_),
    .B1(_00459_),
    .B2(_04513_),
    .Y(_04953_));
 AND2x2_ASAP7_75t_R _11809_ (.A(_03091_),
    .B(_00461_),
    .Y(_04954_));
 AO21x1_ASAP7_75t_R _11810_ (.A1(_03573_),
    .A2(_00460_),
    .B(_04954_),
    .Y(_04955_));
 AO221x1_ASAP7_75t_R _11811_ (.A1(_03130_),
    .A2(_00458_),
    .B1(_03925_),
    .B2(_04955_),
    .C(_03914_),
    .Y(_04956_));
 AO21x1_ASAP7_75t_R _11812_ (.A1(_03029_),
    .A2(_04953_),
    .B(_04956_),
    .Y(_04957_));
 AND2x2_ASAP7_75t_R _11813_ (.A(_04502_),
    .B(_00465_),
    .Y(_04958_));
 AO21x1_ASAP7_75t_R _11814_ (.A1(_03112_),
    .A2(_00464_),
    .B(_04958_),
    .Y(_04959_));
 AND3x1_ASAP7_75t_R _11815_ (.A(_03048_),
    .B(_03034_),
    .C(_00463_),
    .Y(_04960_));
 AO21x1_ASAP7_75t_R _11816_ (.A1(_00462_),
    .A2(_04393_),
    .B(_04960_),
    .Y(_04961_));
 AO221x1_ASAP7_75t_R _11817_ (.A1(_04389_),
    .A2(_04959_),
    .B1(_04961_),
    .B2(_04396_),
    .C(_04397_),
    .Y(_04962_));
 AND3x1_ASAP7_75t_R _11818_ (.A(_03143_),
    .B(_04957_),
    .C(_04962_),
    .Y(_04963_));
 AO22x1_ASAP7_75t_R _11819_ (.A1(_04851_),
    .A2(_00442_),
    .B1(_00443_),
    .B2(_04513_),
    .Y(_04964_));
 AND2x2_ASAP7_75t_R _11820_ (.A(_03091_),
    .B(_00445_),
    .Y(_04965_));
 AO21x1_ASAP7_75t_R _11821_ (.A1(_03573_),
    .A2(_00444_),
    .B(_04965_),
    .Y(_04966_));
 AO221x1_ASAP7_75t_R _11822_ (.A1(_03130_),
    .A2(_00442_),
    .B1(_03925_),
    .B2(_04966_),
    .C(_03914_),
    .Y(_04967_));
 AO21x1_ASAP7_75t_R _11823_ (.A1(_03029_),
    .A2(_04964_),
    .B(_04967_),
    .Y(_04968_));
 AND2x2_ASAP7_75t_R _11824_ (.A(_03898_),
    .B(_00449_),
    .Y(_04969_));
 AO21x1_ASAP7_75t_R _11825_ (.A1(_03112_),
    .A2(_00448_),
    .B(_04969_),
    .Y(_04970_));
 AND3x1_ASAP7_75t_R _11826_ (.A(_03048_),
    .B(_03034_),
    .C(_00447_),
    .Y(_04971_));
 AO21x1_ASAP7_75t_R _11827_ (.A1(_00446_),
    .A2(_04393_),
    .B(_04971_),
    .Y(_04972_));
 AO221x1_ASAP7_75t_R _11828_ (.A1(_04497_),
    .A2(_04970_),
    .B1(_04972_),
    .B2(_04396_),
    .C(_04397_),
    .Y(_04973_));
 AND3x1_ASAP7_75t_R _11829_ (.A(_03703_),
    .B(_04968_),
    .C(_04973_),
    .Y(_04974_));
 OR3x1_ASAP7_75t_R _11830_ (.A(_04545_),
    .B(_04963_),
    .C(_04974_),
    .Y(_04975_));
 OA21x2_ASAP7_75t_R _11831_ (.A1(_03175_),
    .A2(_04952_),
    .B(_04975_),
    .Y(_04976_));
 OAI21x1_ASAP7_75t_R _11832_ (.A1(_03708_),
    .A2(_03642_),
    .B(_03709_),
    .Y(_04977_));
 AND4x1_ASAP7_75t_R _11833_ (.A(_03063_),
    .B(net27),
    .C(_03194_),
    .D(net26),
    .Y(_04978_));
 AND3x4_ASAP7_75t_R _11834_ (.A(_03240_),
    .B(_03267_),
    .C(_04978_),
    .Y(_04979_));
 AO32x1_ASAP7_75t_R _11835_ (.A1(_04784_),
    .A2(_04783_),
    .A3(_04899_),
    .B1(_03539_),
    .B2(_04979_),
    .Y(_04980_));
 INVx2_ASAP7_75t_R _11836_ (.A(_03717_),
    .Y(_04981_));
 OA21x2_ASAP7_75t_R _11837_ (.A1(_04977_),
    .A2(_04980_),
    .B(_04981_),
    .Y(_04982_));
 AO21x1_ASAP7_75t_R _11838_ (.A1(_03192_),
    .A2(_03264_),
    .B(_03241_),
    .Y(_04983_));
 AO21x2_ASAP7_75t_R _11839_ (.A1(_03249_),
    .A2(_04983_),
    .B(_03254_),
    .Y(_04984_));
 INVx2_ASAP7_75t_R _11840_ (.A(_04984_),
    .Y(_04985_));
 OA21x2_ASAP7_75t_R _11841_ (.A1(_03247_),
    .A2(_03861_),
    .B(_03711_),
    .Y(_04986_));
 OR2x2_ASAP7_75t_R _11842_ (.A(_03718_),
    .B(_04985_),
    .Y(_04987_));
 NOR2x1_ASAP7_75t_R _11843_ (.A(_04986_),
    .B(_04987_),
    .Y(_04988_));
 AO21x1_ASAP7_75t_R _11844_ (.A1(_04982_),
    .A2(_04985_),
    .B(_04988_),
    .Y(_09754_));
 NOR2x1_ASAP7_75t_R _11845_ (.A(_04159_),
    .B(_09754_),
    .Y(_04989_));
 AO21x1_ASAP7_75t_R _11846_ (.A1(_04159_),
    .A2(_04976_),
    .B(_04989_),
    .Y(_04990_));
 XNOR2x1_ASAP7_75t_R _11847_ (.B(_04990_),
    .Y(_09621_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _11848_ (.A(_09621_),
    .Y(_09623_));
 OAI22x1_ASAP7_75t_R _11849_ (.A1(_00447_),
    .A2(_04550_),
    .B1(_03410_),
    .B2(_00446_),
    .Y(_04991_));
 OA22x2_ASAP7_75t_R _11850_ (.A1(_00444_),
    .A2(_03735_),
    .B1(_03740_),
    .B2(_00445_),
    .Y(_04992_));
 AND2x2_ASAP7_75t_R _11851_ (.A(_00448_),
    .B(_03334_),
    .Y(_04993_));
 AO221x1_ASAP7_75t_R _11852_ (.A1(_03261_),
    .A2(_04018_),
    .B1(_03994_),
    .B2(_00449_),
    .C(_04993_),
    .Y(_04994_));
 OAI21x1_ASAP7_75t_R _11853_ (.A1(_03472_),
    .A2(_04992_),
    .B(_04994_),
    .Y(_04995_));
 OR2x2_ASAP7_75t_R _11854_ (.A(_00443_),
    .B(_03765_),
    .Y(_04996_));
 OAI21x1_ASAP7_75t_R _11855_ (.A1(_00442_),
    .A2(_03479_),
    .B(_04996_),
    .Y(_04997_));
 AO221x1_ASAP7_75t_R _11856_ (.A1(_03341_),
    .A2(_04995_),
    .B1(_04997_),
    .B2(_03448_),
    .C(_04552_),
    .Y(_04998_));
 AO21x1_ASAP7_75t_R _11857_ (.A1(_04549_),
    .A2(_04991_),
    .B(_04998_),
    .Y(_04999_));
 NAND2x1_ASAP7_75t_R _11858_ (.A(_00434_),
    .B(_04451_),
    .Y(_05000_));
 NAND2x1_ASAP7_75t_R _11859_ (.A(_00435_),
    .B(_03479_),
    .Y(_05001_));
 OAI22x1_ASAP7_75t_R _11860_ (.A1(_00438_),
    .A2(_03330_),
    .B1(_03415_),
    .B2(_00439_),
    .Y(_05002_));
 AO32x1_ASAP7_75t_R _11861_ (.A1(_03448_),
    .A2(_05000_),
    .A3(_05001_),
    .B1(_03483_),
    .B2(_05002_),
    .Y(_05003_));
 NOR2x1_ASAP7_75t_R _11862_ (.A(_00436_),
    .B(_03305_),
    .Y(_05004_));
 INVx1_ASAP7_75t_R _11863_ (.A(_00437_),
    .Y(_05005_));
 OA211x2_ASAP7_75t_R _11864_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03837_),
    .C(_05005_),
    .Y(_05006_));
 OA211x2_ASAP7_75t_R _11865_ (.A1(_05004_),
    .A2(_05006_),
    .B(_04574_),
    .C(_04575_),
    .Y(_05007_));
 AND2x2_ASAP7_75t_R _11866_ (.A(_00440_),
    .B(_03436_),
    .Y(_05008_));
 AOI221x1_ASAP7_75t_R _11867_ (.A1(_03251_),
    .A2(_03388_),
    .B1(_03735_),
    .B2(_00441_),
    .C(_05008_),
    .Y(_05009_));
 OA21x2_ASAP7_75t_R _11868_ (.A1(_05007_),
    .A2(_05009_),
    .B(_04432_),
    .Y(_05010_));
 OA21x2_ASAP7_75t_R _11869_ (.A1(_03461_),
    .A2(_05010_),
    .B(_03246_),
    .Y(_05011_));
 OA21x2_ASAP7_75t_R _11870_ (.A1(_05003_),
    .A2(_05011_),
    .B(_03499_),
    .Y(_05012_));
 INVx1_ASAP7_75t_R _11871_ (.A(_00451_),
    .Y(_05013_));
 NAND2x1_ASAP7_75t_R _11872_ (.A(_00450_),
    .B(_03383_),
    .Y(_05014_));
 OA211x2_ASAP7_75t_R _11873_ (.A1(_05013_),
    .A2(_03451_),
    .B(_04469_),
    .C(_05014_),
    .Y(_05015_));
 OA22x2_ASAP7_75t_R _11874_ (.A1(_00452_),
    .A2(_03329_),
    .B1(_03414_),
    .B2(_00453_),
    .Y(_05016_));
 AND3x1_ASAP7_75t_R _11875_ (.A(_03063_),
    .B(_04586_),
    .C(_00457_),
    .Y(_05017_));
 AO221x1_ASAP7_75t_R _11876_ (.A1(_03261_),
    .A2(_04575_),
    .B1(_03847_),
    .B2(_00456_),
    .C(_05017_),
    .Y(_05018_));
 OAI21x1_ASAP7_75t_R _11877_ (.A1(_03441_),
    .A2(_05016_),
    .B(_05018_),
    .Y(_05019_));
 OAI22x1_ASAP7_75t_R _11878_ (.A1(_00454_),
    .A2(_03350_),
    .B1(_03357_),
    .B2(_00455_),
    .Y(_05020_));
 AO221x1_ASAP7_75t_R _11879_ (.A1(_04026_),
    .A2(_05019_),
    .B1(_05020_),
    .B2(_03540_),
    .C(_03461_),
    .Y(_05021_));
 INVx1_ASAP7_75t_R _11880_ (.A(_00459_),
    .Y(_05022_));
 NAND2x1_ASAP7_75t_R _11881_ (.A(_00458_),
    .B(_03383_),
    .Y(_05023_));
 OA211x2_ASAP7_75t_R _11882_ (.A1(_05022_),
    .A2(_03451_),
    .B(_04469_),
    .C(_05023_),
    .Y(_05024_));
 OA22x2_ASAP7_75t_R _11883_ (.A1(_00460_),
    .A2(_03994_),
    .B1(_03765_),
    .B2(_00461_),
    .Y(_05025_));
 AND3x1_ASAP7_75t_R _11884_ (.A(_03063_),
    .B(_04586_),
    .C(_00465_),
    .Y(_05026_));
 AO221x1_ASAP7_75t_R _11885_ (.A1(_03261_),
    .A2(_04575_),
    .B1(_03847_),
    .B2(_00464_),
    .C(_05026_),
    .Y(_05027_));
 OAI21x1_ASAP7_75t_R _11886_ (.A1(_03441_),
    .A2(_05025_),
    .B(_05027_),
    .Y(_05028_));
 OAI22x1_ASAP7_75t_R _11887_ (.A1(_00463_),
    .A2(_03397_),
    .B1(_03401_),
    .B2(_00462_),
    .Y(_05029_));
 AO221x1_ASAP7_75t_R _11888_ (.A1(_04026_),
    .A2(_05028_),
    .B1(_05029_),
    .B2(_03540_),
    .C(_04552_),
    .Y(_05030_));
 OA22x2_ASAP7_75t_R _11889_ (.A1(_05015_),
    .A2(_05021_),
    .B1(_05024_),
    .B2(_05030_),
    .Y(_05031_));
 BUFx6f_ASAP7_75t_R _11890_ (.A(_03495_),
    .Y(_05032_));
 AO22x2_ASAP7_75t_R _11891_ (.A1(_04999_),
    .A2(_05012_),
    .B1(_05031_),
    .B2(_05032_),
    .Y(_05033_));
 BUFx6f_ASAP7_75t_R _11892_ (.A(_05033_),
    .Y(_09620_));
 INVx1_ASAP7_75t_R _11893_ (.A(_09620_),
    .Y(_09622_));
 BUFx6f_ASAP7_75t_R _11894_ (.A(_03586_),
    .Y(_05034_));
 AND2x2_ASAP7_75t_R _11895_ (.A(_04390_),
    .B(_00470_),
    .Y(_05035_));
 AO21x1_ASAP7_75t_R _11896_ (.A1(_04851_),
    .A2(_00469_),
    .B(_05035_),
    .Y(_05036_));
 AO21x1_ASAP7_75t_R _11897_ (.A1(_04850_),
    .A2(_05036_),
    .B(_03078_),
    .Y(_05037_));
 AO22x1_ASAP7_75t_R _11898_ (.A1(_04498_),
    .A2(_00467_),
    .B1(_00468_),
    .B2(_04361_),
    .Y(_05038_));
 AO22x1_ASAP7_75t_R _11899_ (.A1(_03098_),
    .A2(_00467_),
    .B1(_05038_),
    .B2(_04381_),
    .Y(_05039_));
 AO21x1_ASAP7_75t_R _11900_ (.A1(_03216_),
    .A2(_05037_),
    .B(_05039_),
    .Y(_05040_));
 BUFx6f_ASAP7_75t_R _11901_ (.A(_03074_),
    .Y(_05041_));
 AND2x2_ASAP7_75t_R _11902_ (.A(_03092_),
    .B(_00474_),
    .Y(_05042_));
 AO21x1_ASAP7_75t_R _11903_ (.A1(_04095_),
    .A2(_00473_),
    .B(_05042_),
    .Y(_05043_));
 BUFx6f_ASAP7_75t_R _11904_ (.A(_04267_),
    .Y(_05044_));
 AND3x1_ASAP7_75t_R _11905_ (.A(_05044_),
    .B(_03045_),
    .C(_00472_),
    .Y(_05045_));
 AO21x1_ASAP7_75t_R _11906_ (.A1(_00471_),
    .A2(_03290_),
    .B(_05045_),
    .Y(_05046_));
 AO221x1_ASAP7_75t_R _11907_ (.A1(_05041_),
    .A2(_05043_),
    .B1(_05046_),
    .B2(_04856_),
    .C(_04411_),
    .Y(_05047_));
 AND3x1_ASAP7_75t_R _11908_ (.A(_05034_),
    .B(_05040_),
    .C(_05047_),
    .Y(_05048_));
 AND2x2_ASAP7_75t_R _11909_ (.A(_03092_),
    .B(_00482_),
    .Y(_05049_));
 AO21x1_ASAP7_75t_R _11910_ (.A1(_04080_),
    .A2(_00481_),
    .B(_05049_),
    .Y(_05050_));
 AND3x1_ASAP7_75t_R _11911_ (.A(_05044_),
    .B(_03045_),
    .C(_00480_),
    .Y(_05051_));
 AO21x1_ASAP7_75t_R _11912_ (.A1(_00479_),
    .A2(_03290_),
    .B(_05051_),
    .Y(_05052_));
 AO221x1_ASAP7_75t_R _11913_ (.A1(_05041_),
    .A2(_05050_),
    .B1(_05052_),
    .B2(_04856_),
    .C(_04411_),
    .Y(_05053_));
 AO22x1_ASAP7_75t_R _11914_ (.A1(_03139_),
    .A2(_00475_),
    .B1(_00476_),
    .B2(_04513_),
    .Y(_05054_));
 AND2x2_ASAP7_75t_R _11915_ (.A(_04390_),
    .B(_00478_),
    .Y(_05055_));
 AO21x1_ASAP7_75t_R _11916_ (.A1(_03566_),
    .A2(_00477_),
    .B(_05055_),
    .Y(_05056_));
 AO21x1_ASAP7_75t_R _11917_ (.A1(_04389_),
    .A2(_05056_),
    .B(_03078_),
    .Y(_05057_));
 AO21x1_ASAP7_75t_R _11918_ (.A1(_03137_),
    .A2(_05054_),
    .B(_05057_),
    .Y(_05058_));
 AND3x1_ASAP7_75t_R _11919_ (.A(_03174_),
    .B(_05053_),
    .C(_05058_),
    .Y(_05059_));
 NOR3x1_ASAP7_75t_R _11920_ (.A(_04486_),
    .B(_05048_),
    .C(_05059_),
    .Y(_05060_));
 BUFx6f_ASAP7_75t_R _11921_ (.A(_03697_),
    .Y(_05061_));
 AND2x2_ASAP7_75t_R _11922_ (.A(_03107_),
    .B(_00485_),
    .Y(_05062_));
 AO21x1_ASAP7_75t_R _11923_ (.A1(_03904_),
    .A2(_00483_),
    .B(_05062_),
    .Y(_05063_));
 BUFx6f_ASAP7_75t_R _11924_ (.A(_03082_),
    .Y(_05064_));
 AO22x1_ASAP7_75t_R _11925_ (.A1(_00486_),
    .A2(_05061_),
    .B1(_05063_),
    .B2(_05064_),
    .Y(_05065_));
 BUFx6f_ASAP7_75t_R _11926_ (.A(_03561_),
    .Y(_05066_));
 BUFx6f_ASAP7_75t_R _11927_ (.A(_04862_),
    .Y(_05067_));
 AO21x1_ASAP7_75t_R _11928_ (.A1(_00484_),
    .A2(_05066_),
    .B(_05067_),
    .Y(_05068_));
 BUFx6f_ASAP7_75t_R _11929_ (.A(_03893_),
    .Y(_05069_));
 BUFx6f_ASAP7_75t_R _11930_ (.A(_04087_),
    .Y(_05070_));
 AND2x2_ASAP7_75t_R _11931_ (.A(_05070_),
    .B(_00490_),
    .Y(_05071_));
 AO21x1_ASAP7_75t_R _11932_ (.A1(_03139_),
    .A2(_00489_),
    .B(_05071_),
    .Y(_05072_));
 BUFx10_ASAP7_75t_R _11933_ (.A(_03577_),
    .Y(_05073_));
 AND3x1_ASAP7_75t_R _11934_ (.A(_03041_),
    .B(_03200_),
    .C(_00488_),
    .Y(_05074_));
 AO21x1_ASAP7_75t_R _11935_ (.A1(_00487_),
    .A2(_05073_),
    .B(_05074_),
    .Y(_05075_));
 BUFx6f_ASAP7_75t_R _11936_ (.A(_04074_),
    .Y(_05076_));
 BUFx6f_ASAP7_75t_R _11937_ (.A(_04379_),
    .Y(_05077_));
 AO221x1_ASAP7_75t_R _11938_ (.A1(_05069_),
    .A2(_05072_),
    .B1(_05075_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_05078_));
 OA21x2_ASAP7_75t_R _11939_ (.A1(_05065_),
    .A2(_05068_),
    .B(_05078_),
    .Y(_05079_));
 AND2x2_ASAP7_75t_R _11940_ (.A(_03571_),
    .B(_00493_),
    .Y(_05080_));
 AO21x1_ASAP7_75t_R _11941_ (.A1(_04381_),
    .A2(_00491_),
    .B(_05080_),
    .Y(_05081_));
 AO22x1_ASAP7_75t_R _11942_ (.A1(_00494_),
    .A2(_05061_),
    .B1(_05081_),
    .B2(_05064_),
    .Y(_05082_));
 AO21x1_ASAP7_75t_R _11943_ (.A1(_00492_),
    .A2(_05066_),
    .B(_05067_),
    .Y(_05083_));
 AND2x2_ASAP7_75t_R _11944_ (.A(_03092_),
    .B(_00498_),
    .Y(_05084_));
 AO21x1_ASAP7_75t_R _11945_ (.A1(_04080_),
    .A2(_00497_),
    .B(_05084_),
    .Y(_05085_));
 AND3x1_ASAP7_75t_R _11946_ (.A(_05044_),
    .B(_03045_),
    .C(_00496_),
    .Y(_05086_));
 AO21x1_ASAP7_75t_R _11947_ (.A1(_00495_),
    .A2(_03290_),
    .B(_05086_),
    .Y(_05087_));
 AO221x1_ASAP7_75t_R _11948_ (.A1(_05041_),
    .A2(_05085_),
    .B1(_05087_),
    .B2(_04856_),
    .C(_04411_),
    .Y(_05088_));
 OA211x2_ASAP7_75t_R _11949_ (.A1(_05082_),
    .A2(_05083_),
    .B(_03174_),
    .C(_05088_),
    .Y(_05089_));
 AOI211x1_ASAP7_75t_R _11950_ (.A1(_04545_),
    .A2(_05079_),
    .B(_05089_),
    .C(_04423_),
    .Y(_05090_));
 OAI21x1_ASAP7_75t_R _11951_ (.A1(_05060_),
    .A2(_05090_),
    .B(_03705_),
    .Y(_05091_));
 BUFx4f_ASAP7_75t_R _11952_ (.A(_04984_),
    .Y(_05092_));
 BUFx12f_ASAP7_75t_R _11953_ (.A(_03472_),
    .Y(_05093_));
 AO32x1_ASAP7_75t_R _11954_ (.A1(_04784_),
    .A2(_04783_),
    .A3(_05093_),
    .B1(_04899_),
    .B2(_04979_),
    .Y(_05094_));
 OA21x2_ASAP7_75t_R _11955_ (.A1(_04977_),
    .A2(_05094_),
    .B(_04981_),
    .Y(_05095_));
 AND2x2_ASAP7_75t_R _11956_ (.A(_04985_),
    .B(_05095_),
    .Y(_05096_));
 AO21x1_ASAP7_75t_R _11957_ (.A1(_04982_),
    .A2(_05092_),
    .B(_05096_),
    .Y(_09752_));
 NOR2x1_ASAP7_75t_R _11958_ (.A(_04159_),
    .B(_09752_),
    .Y(_05097_));
 AO21x1_ASAP7_75t_R _11959_ (.A1(_04159_),
    .A2(_05091_),
    .B(_05097_),
    .Y(_05098_));
 XNOR2x1_ASAP7_75t_R _11960_ (.B(_05098_),
    .Y(_09626_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _11961_ (.A(_09626_),
    .Y(_09628_));
 INVx1_ASAP7_75t_R _11962_ (.A(_00476_),
    .Y(_05099_));
 NAND2x1_ASAP7_75t_R _11963_ (.A(_00475_),
    .B(_04153_),
    .Y(_05100_));
 OA211x2_ASAP7_75t_R _11964_ (.A1(_05099_),
    .A2(_03486_),
    .B(_05100_),
    .C(_03393_),
    .Y(_05101_));
 OR3x1_ASAP7_75t_R _11965_ (.A(_03277_),
    .B(_03550_),
    .C(_03381_),
    .Y(_05102_));
 OAI22x1_ASAP7_75t_R _11966_ (.A1(_00480_),
    .A2(_03847_),
    .B1(_03400_),
    .B2(_00479_),
    .Y(_05103_));
 AND2x2_ASAP7_75t_R _11967_ (.A(_03747_),
    .B(_05103_),
    .Y(_05104_));
 OR4x1_ASAP7_75t_R _11968_ (.A(_03344_),
    .B(_05101_),
    .C(_05102_),
    .D(_05104_),
    .Y(_05105_));
 BUFx12_ASAP7_75t_R _11969_ (.A(_04022_),
    .Y(_05106_));
 AND3x1_ASAP7_75t_R _11970_ (.A(_00477_),
    .B(_03261_),
    .C(_04018_),
    .Y(_05107_));
 AOI211x1_ASAP7_75t_R _11971_ (.A1(_00481_),
    .A2(_04444_),
    .B(_05106_),
    .C(_05107_),
    .Y(_05108_));
 OAI22x1_ASAP7_75t_R _11972_ (.A1(_00482_),
    .A2(_03732_),
    .B1(_03733_),
    .B2(_00478_),
    .Y(_05109_));
 OR4x2_ASAP7_75t_R _11973_ (.A(_04786_),
    .B(_03405_),
    .C(_05108_),
    .D(_05109_),
    .Y(_05110_));
 AND3x1_ASAP7_75t_R _11974_ (.A(_03499_),
    .B(_05105_),
    .C(_05110_),
    .Y(_05111_));
 AND3x1_ASAP7_75t_R _11975_ (.A(_00469_),
    .B(_03251_),
    .C(_03388_),
    .Y(_05112_));
 AO21x1_ASAP7_75t_R _11976_ (.A1(_00473_),
    .A2(_03472_),
    .B(_05112_),
    .Y(_05113_));
 OA222x2_ASAP7_75t_R _11977_ (.A1(_00474_),
    .A2(_03732_),
    .B1(_05113_),
    .B2(_04440_),
    .C1(_03733_),
    .C2(_00470_),
    .Y(_05114_));
 OA22x2_ASAP7_75t_R _11978_ (.A1(_00471_),
    .A2(_04560_),
    .B1(_03450_),
    .B2(_00472_),
    .Y(_05115_));
 OA21x2_ASAP7_75t_R _11979_ (.A1(_03979_),
    .A2(_05115_),
    .B(_04771_),
    .Y(_05116_));
 AND2x2_ASAP7_75t_R _11980_ (.A(_00468_),
    .B(_04466_),
    .Y(_05117_));
 AO21x1_ASAP7_75t_R _11981_ (.A1(_00467_),
    .A2(_04472_),
    .B(_05117_),
    .Y(_05118_));
 OA22x2_ASAP7_75t_R _11982_ (.A1(_03344_),
    .A2(_05116_),
    .B1(_05118_),
    .B2(_04450_),
    .Y(_05119_));
 OAI21x1_ASAP7_75t_R _11983_ (.A1(_04214_),
    .A2(_05114_),
    .B(_05119_),
    .Y(_05120_));
 OA21x2_ASAP7_75t_R _11984_ (.A1(_00493_),
    .A2(_03384_),
    .B(_03736_),
    .Y(_05121_));
 OA21x2_ASAP7_75t_R _11985_ (.A1(_00494_),
    .A2(_03414_),
    .B(_05121_),
    .Y(_05122_));
 OR2x2_ASAP7_75t_R _11986_ (.A(_03988_),
    .B(_05122_),
    .Y(_05123_));
 BUFx12_ASAP7_75t_R _11987_ (.A(_04586_),
    .Y(_05124_));
 AND3x1_ASAP7_75t_R _11988_ (.A(_03200_),
    .B(_05124_),
    .C(_00498_),
    .Y(_05125_));
 AO21x1_ASAP7_75t_R _11989_ (.A1(_00497_),
    .A2(_03377_),
    .B(_05125_),
    .Y(_05126_));
 BUFx12f_ASAP7_75t_R _11990_ (.A(_04444_),
    .Y(_05127_));
 AOI22x1_ASAP7_75t_R _11991_ (.A1(_03210_),
    .A2(_05123_),
    .B1(_05126_),
    .B2(_05127_),
    .Y(_05128_));
 OR2x2_ASAP7_75t_R _11992_ (.A(_00491_),
    .B(_03467_),
    .Y(_05129_));
 OAI21x1_ASAP7_75t_R _11993_ (.A1(_00492_),
    .A2(_03383_),
    .B(_05129_),
    .Y(_05130_));
 OAI22x1_ASAP7_75t_R _11994_ (.A1(_00496_),
    .A2(_03397_),
    .B1(_03401_),
    .B2(_00495_),
    .Y(_05131_));
 AO221x1_ASAP7_75t_R _11995_ (.A1(_04469_),
    .A2(_05130_),
    .B1(_05131_),
    .B2(_03362_),
    .C(_04552_),
    .Y(_05132_));
 AND3x1_ASAP7_75t_R _11996_ (.A(_04503_),
    .B(_03475_),
    .C(_00490_),
    .Y(_05133_));
 AO21x1_ASAP7_75t_R _11997_ (.A1(_00489_),
    .A2(_03437_),
    .B(_05133_),
    .Y(_05134_));
 AO21x1_ASAP7_75t_R _11998_ (.A1(_03472_),
    .A2(_05134_),
    .B(_04786_),
    .Y(_05135_));
 OA21x2_ASAP7_75t_R _11999_ (.A1(_00485_),
    .A2(_03329_),
    .B(_03550_),
    .Y(_05136_));
 OA211x2_ASAP7_75t_R _12000_ (.A1(_00486_),
    .A2(_04676_),
    .B(_05136_),
    .C(_04447_),
    .Y(_05137_));
 AOI211x1_ASAP7_75t_R _12001_ (.A1(_04771_),
    .A2(_05135_),
    .B(_05137_),
    .C(_03862_),
    .Y(_05138_));
 OAI22x1_ASAP7_75t_R _12002_ (.A1(_00487_),
    .A2(_03385_),
    .B1(_03414_),
    .B2(_00488_),
    .Y(_05139_));
 AND2x2_ASAP7_75t_R _12003_ (.A(_03361_),
    .B(_05139_),
    .Y(_05140_));
 INVx1_ASAP7_75t_R _12004_ (.A(_00484_),
    .Y(_05141_));
 NAND2x1_ASAP7_75t_R _12005_ (.A(_00483_),
    .B(_03418_),
    .Y(_05142_));
 OA211x2_ASAP7_75t_R _12006_ (.A1(_05141_),
    .A2(_04005_),
    .B(_03420_),
    .C(_05142_),
    .Y(_05143_));
 OA211x2_ASAP7_75t_R _12007_ (.A1(_05140_),
    .A2(_05143_),
    .B(_03521_),
    .C(_03539_),
    .Y(_05144_));
 OA22x2_ASAP7_75t_R _12008_ (.A1(_05128_),
    .A2(_05132_),
    .B1(_05138_),
    .B2(_05144_),
    .Y(_05145_));
 AO21x2_ASAP7_75t_R _12009_ (.A1(_05111_),
    .A2(_05120_),
    .B(_05145_),
    .Y(_05146_));
 BUFx6f_ASAP7_75t_R _12010_ (.A(_05146_),
    .Y(_09625_));
 INVx1_ASAP7_75t_R _12011_ (.A(_09625_),
    .Y(_09627_));
 AO22x1_ASAP7_75t_R _12012_ (.A1(_03945_),
    .A2(_00500_),
    .B1(_00501_),
    .B2(_03946_),
    .Y(_05147_));
 AND2x2_ASAP7_75t_R _12013_ (.A(_03047_),
    .B(_00503_),
    .Y(_05148_));
 AO21x1_ASAP7_75t_R _12014_ (.A1(_03630_),
    .A2(_00502_),
    .B(_05148_),
    .Y(_05149_));
 AO21x1_ASAP7_75t_R _12015_ (.A1(_03087_),
    .A2(_05149_),
    .B(_03077_),
    .Y(_05150_));
 AND2x2_ASAP7_75t_R _12016_ (.A(_03097_),
    .B(_00500_),
    .Y(_05151_));
 AO221x1_ASAP7_75t_R _12017_ (.A1(_03068_),
    .A2(_05147_),
    .B1(_05150_),
    .B2(_03215_),
    .C(_05151_),
    .Y(_05152_));
 BUFx10_ASAP7_75t_R _12018_ (.A(_03055_),
    .Y(_05153_));
 AND2x2_ASAP7_75t_R _12019_ (.A(_03040_),
    .B(_00507_),
    .Y(_05154_));
 AO21x1_ASAP7_75t_R _12020_ (.A1(_05153_),
    .A2(_00506_),
    .B(_05154_),
    .Y(_05155_));
 AND3x1_ASAP7_75t_R _12021_ (.A(_04087_),
    .B(_04692_),
    .C(_00505_),
    .Y(_05156_));
 AO21x1_ASAP7_75t_R _12022_ (.A1(_00504_),
    .A2(_04376_),
    .B(_05156_),
    .Y(_05157_));
 AO221x2_ASAP7_75t_R _12023_ (.A1(_04487_),
    .A2(_05155_),
    .B1(_05157_),
    .B2(_04074_),
    .C(_04379_),
    .Y(_05158_));
 AND3x1_ASAP7_75t_R _12024_ (.A(_04085_),
    .B(_05152_),
    .C(_05158_),
    .Y(_05159_));
 AND2x2_ASAP7_75t_R _12025_ (.A(_03040_),
    .B(_00515_),
    .Y(_05160_));
 AO21x1_ASAP7_75t_R _12026_ (.A1(_05153_),
    .A2(_00514_),
    .B(_05160_),
    .Y(_05161_));
 AND3x1_ASAP7_75t_R _12027_ (.A(_04087_),
    .B(_04692_),
    .C(_00513_),
    .Y(_05162_));
 AO21x1_ASAP7_75t_R _12028_ (.A1(_00512_),
    .A2(_04376_),
    .B(_05162_),
    .Y(_05163_));
 AO221x1_ASAP7_75t_R _12029_ (.A1(_04487_),
    .A2(_05161_),
    .B1(_05163_),
    .B2(_03582_),
    .C(_04379_),
    .Y(_05164_));
 AO22x1_ASAP7_75t_R _12030_ (.A1(_03685_),
    .A2(_00508_),
    .B1(_00509_),
    .B2(_04361_),
    .Y(_05165_));
 AND2x2_ASAP7_75t_R _12031_ (.A(_03091_),
    .B(_00511_),
    .Y(_05166_));
 AO21x1_ASAP7_75t_R _12032_ (.A1(_03573_),
    .A2(_00510_),
    .B(_05166_),
    .Y(_05167_));
 AO21x1_ASAP7_75t_R _12033_ (.A1(_03107_),
    .A2(_05167_),
    .B(_03623_),
    .Y(_05168_));
 AO21x1_ASAP7_75t_R _12034_ (.A1(_04381_),
    .A2(_05165_),
    .B(_05168_),
    .Y(_05169_));
 AND3x1_ASAP7_75t_R _12035_ (.A(_03119_),
    .B(_05164_),
    .C(_05169_),
    .Y(_05170_));
 OR3x1_ASAP7_75t_R _12036_ (.A(_04043_),
    .B(_05159_),
    .C(_05170_),
    .Y(_05171_));
 AND2x2_ASAP7_75t_R _12037_ (.A(_03040_),
    .B(_00531_),
    .Y(_05172_));
 AO21x1_ASAP7_75t_R _12038_ (.A1(_05153_),
    .A2(_00530_),
    .B(_05172_),
    .Y(_05173_));
 AND3x1_ASAP7_75t_R _12039_ (.A(_04087_),
    .B(_04692_),
    .C(_00529_),
    .Y(_05174_));
 AO21x1_ASAP7_75t_R _12040_ (.A1(_00528_),
    .A2(_04376_),
    .B(_05174_),
    .Y(_05175_));
 AO221x1_ASAP7_75t_R _12041_ (.A1(_04487_),
    .A2(_05173_),
    .B1(_05175_),
    .B2(_04074_),
    .C(_04379_),
    .Y(_05176_));
 AND2x2_ASAP7_75t_R _12042_ (.A(_03647_),
    .B(_00526_),
    .Y(_05177_));
 AO21x1_ASAP7_75t_R _12043_ (.A1(_03160_),
    .A2(_00524_),
    .B(_05177_),
    .Y(_05178_));
 AO21x1_ASAP7_75t_R _12044_ (.A1(_00525_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_05179_));
 AO221x1_ASAP7_75t_R _12045_ (.A1(_00527_),
    .A2(_03697_),
    .B1(_05178_),
    .B2(_04080_),
    .C(_05179_),
    .Y(_05180_));
 AND3x1_ASAP7_75t_R _12046_ (.A(_03119_),
    .B(_05176_),
    .C(_05180_),
    .Y(_05181_));
 AND2x2_ASAP7_75t_R _12047_ (.A(_03040_),
    .B(_00523_),
    .Y(_05182_));
 AO21x1_ASAP7_75t_R _12048_ (.A1(_05153_),
    .A2(_00522_),
    .B(_05182_),
    .Y(_05183_));
 AND3x1_ASAP7_75t_R _12049_ (.A(_03065_),
    .B(_04692_),
    .C(_00521_),
    .Y(_05184_));
 AO21x1_ASAP7_75t_R _12050_ (.A1(_00520_),
    .A2(_04376_),
    .B(_05184_),
    .Y(_05185_));
 AO221x1_ASAP7_75t_R _12051_ (.A1(_04722_),
    .A2(_05183_),
    .B1(_05185_),
    .B2(_03582_),
    .C(_04379_),
    .Y(_05186_));
 AND2x2_ASAP7_75t_R _12052_ (.A(_03647_),
    .B(_00518_),
    .Y(_05187_));
 AO21x1_ASAP7_75t_R _12053_ (.A1(_03160_),
    .A2(_00516_),
    .B(_05187_),
    .Y(_05188_));
 AO21x1_ASAP7_75t_R _12054_ (.A1(_00517_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_05189_));
 AO221x1_ASAP7_75t_R _12055_ (.A1(_00519_),
    .A2(_03697_),
    .B1(_05188_),
    .B2(_04080_),
    .C(_05189_),
    .Y(_05190_));
 AND3x1_ASAP7_75t_R _12056_ (.A(_04085_),
    .B(_05186_),
    .C(_05190_),
    .Y(_05191_));
 OR3x2_ASAP7_75t_R _12057_ (.A(_04100_),
    .B(_05181_),
    .C(_05191_),
    .Y(_05192_));
 AND2x2_ASAP7_75t_R _12058_ (.A(_05171_),
    .B(_05192_),
    .Y(_05193_));
 OR2x4_ASAP7_75t_R _12059_ (.A(_04163_),
    .B(_05193_),
    .Y(_05194_));
 BUFx10_ASAP7_75t_R _12060_ (.A(_04026_),
    .Y(_05195_));
 AOI22x1_ASAP7_75t_R _12061_ (.A1(_03345_),
    .A2(_05195_),
    .B1(_05093_),
    .B2(_04979_),
    .Y(_05196_));
 AO21x1_ASAP7_75t_R _12062_ (.A1(_03710_),
    .A2(_05196_),
    .B(_03718_),
    .Y(_05197_));
 NOR2x1_ASAP7_75t_R _12063_ (.A(_05092_),
    .B(_05197_),
    .Y(_05198_));
 AO21x1_ASAP7_75t_R _12064_ (.A1(_05092_),
    .A2(_05095_),
    .B(_05198_),
    .Y(_09750_));
 NOR2x1_ASAP7_75t_R _12065_ (.A(_04159_),
    .B(_09750_),
    .Y(_05199_));
 AO21x1_ASAP7_75t_R _12066_ (.A1(_04159_),
    .A2(_05194_),
    .B(_05199_),
    .Y(_05200_));
 XNOR2x1_ASAP7_75t_R _12067_ (.B(_05200_),
    .Y(_09631_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _12068_ (.A(_09631_),
    .Y(_09633_));
 AND2x2_ASAP7_75t_R _12069_ (.A(_00516_),
    .B(_04445_),
    .Y(_05201_));
 AO221x2_ASAP7_75t_R _12070_ (.A1(_00517_),
    .A2(_04768_),
    .B1(_03411_),
    .B2(_03246_),
    .C(_05201_),
    .Y(_05202_));
 AND3x1_ASAP7_75t_R _12071_ (.A(_03064_),
    .B(_05124_),
    .C(_00523_),
    .Y(_05203_));
 AOI221x1_ASAP7_75t_R _12072_ (.A1(_03317_),
    .A2(_03322_),
    .B1(_04480_),
    .B2(_00522_),
    .C(_05203_),
    .Y(_05204_));
 INVx1_ASAP7_75t_R _12073_ (.A(_00519_),
    .Y(_05205_));
 OA211x2_ASAP7_75t_R _12074_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03305_),
    .C(_05205_),
    .Y(_05206_));
 NOR2x1_ASAP7_75t_R _12075_ (.A(_00518_),
    .B(_03329_),
    .Y(_05207_));
 OA211x2_ASAP7_75t_R _12076_ (.A1(_05206_),
    .A2(_05207_),
    .B(_03209_),
    .C(_04020_),
    .Y(_05208_));
 OAI21x1_ASAP7_75t_R _12077_ (.A1(_05204_),
    .A2(_05208_),
    .B(_03341_),
    .Y(_05209_));
 OA22x2_ASAP7_75t_R _12078_ (.A1(_00520_),
    .A2(_03735_),
    .B1(_03740_),
    .B2(_00521_),
    .Y(_05210_));
 OA21x2_ASAP7_75t_R _12079_ (.A1(_03979_),
    .A2(_05210_),
    .B(_04771_),
    .Y(_05211_));
 AO21x1_ASAP7_75t_R _12080_ (.A1(_05209_),
    .A2(_05211_),
    .B(_03344_),
    .Y(_05212_));
 OAI22x1_ASAP7_75t_R _12081_ (.A1(_00529_),
    .A2(_03377_),
    .B1(_04768_),
    .B2(_00528_),
    .Y(_05213_));
 NAND2x2_ASAP7_75t_R _12082_ (.A(_04891_),
    .B(_05213_),
    .Y(_05214_));
 INVx1_ASAP7_75t_R _12083_ (.A(_00525_),
    .Y(_05215_));
 NAND2x1_ASAP7_75t_R _12084_ (.A(_00524_),
    .B(_03722_),
    .Y(_05216_));
 OA211x2_ASAP7_75t_R _12085_ (.A1(_05215_),
    .A2(_04676_),
    .B(_03484_),
    .C(_05216_),
    .Y(_05217_));
 AND3x1_ASAP7_75t_R _12086_ (.A(_03034_),
    .B(_03475_),
    .C(_00531_),
    .Y(_05218_));
 AOI21x1_ASAP7_75t_R _12087_ (.A1(_00530_),
    .A2(_03976_),
    .B(_05218_),
    .Y(_05219_));
 OA21x2_ASAP7_75t_R _12088_ (.A1(_00526_),
    .A2(_04022_),
    .B(_04575_),
    .Y(_05220_));
 OAI21x1_ASAP7_75t_R _12089_ (.A1(_00527_),
    .A2(_03722_),
    .B(_05220_),
    .Y(_05221_));
 OA211x2_ASAP7_75t_R _12090_ (.A1(_04447_),
    .A2(_05219_),
    .B(_05221_),
    .C(_03382_),
    .Y(_05222_));
 NOR3x2_ASAP7_75t_R _12091_ (.B(_05217_),
    .C(_05222_),
    .Y(_05223_),
    .A(_03406_));
 AO221x2_ASAP7_75t_R _12092_ (.A1(_05202_),
    .A2(_05212_),
    .B1(_05214_),
    .B2(_05223_),
    .C(_04003_),
    .Y(_05224_));
 INVx1_ASAP7_75t_R _12093_ (.A(_00500_),
    .Y(_01230_));
 NAND2x1_ASAP7_75t_R _12094_ (.A(_00501_),
    .B(_03541_),
    .Y(_05225_));
 OA21x2_ASAP7_75t_R _12095_ (.A1(_01230_),
    .A2(_03479_),
    .B(_05225_),
    .Y(_05226_));
 BUFx12_ASAP7_75t_R _12096_ (.A(_03306_),
    .Y(_05227_));
 OAI22x1_ASAP7_75t_R _12097_ (.A1(_00504_),
    .A2(_05227_),
    .B1(_03451_),
    .B2(_00505_),
    .Y(_05228_));
 BUFx6f_ASAP7_75t_R _12098_ (.A(_03149_),
    .Y(_05229_));
 OAI22x1_ASAP7_75t_R _12099_ (.A1(_00502_),
    .A2(_04023_),
    .B1(_03722_),
    .B2(_00503_),
    .Y(_05230_));
 AND2x2_ASAP7_75t_R _12100_ (.A(_00506_),
    .B(_03975_),
    .Y(_05231_));
 AOI221x1_ASAP7_75t_R _12101_ (.A1(_03209_),
    .A2(_04020_),
    .B1(_04560_),
    .B2(_00507_),
    .C(_05231_),
    .Y(_05232_));
 AO221x1_ASAP7_75t_R _12102_ (.A1(_05229_),
    .A2(net9),
    .B1(_04447_),
    .B2(_05230_),
    .C(_05232_),
    .Y(_05233_));
 AO222x2_ASAP7_75t_R _12103_ (.A1(_03448_),
    .A2(_05226_),
    .B1(_05228_),
    .B2(_04891_),
    .C1(_04349_),
    .C2(_05233_),
    .Y(_05234_));
 OA21x2_ASAP7_75t_R _12104_ (.A1(_00510_),
    .A2(_03994_),
    .B(_04441_),
    .Y(_05235_));
 OAI21x1_ASAP7_75t_R _12105_ (.A1(_00511_),
    .A2(_04473_),
    .B(_05235_),
    .Y(_05236_));
 AO21x1_ASAP7_75t_R _12106_ (.A1(_03382_),
    .A2(_05236_),
    .B(_03278_),
    .Y(_05237_));
 AND3x1_ASAP7_75t_R _12107_ (.A(_03064_),
    .B(_05124_),
    .C(_00515_),
    .Y(_05238_));
 AO21x1_ASAP7_75t_R _12108_ (.A1(_00514_),
    .A2(_04480_),
    .B(_05238_),
    .Y(_05239_));
 NAND2x1_ASAP7_75t_R _12109_ (.A(_04885_),
    .B(_05239_),
    .Y(_05240_));
 BUFx10_ASAP7_75t_R _12110_ (.A(_03722_),
    .Y(_05241_));
 OR2x2_ASAP7_75t_R _12111_ (.A(_00508_),
    .B(_04466_),
    .Y(_05242_));
 OAI21x1_ASAP7_75t_R _12112_ (.A1(_00509_),
    .A2(_05241_),
    .B(_05242_),
    .Y(_05243_));
 OAI22x1_ASAP7_75t_R _12113_ (.A1(_00513_),
    .A2(_03976_),
    .B1(_04466_),
    .B2(_00512_),
    .Y(_05244_));
 AO221x1_ASAP7_75t_R _12114_ (.A1(_04784_),
    .A2(_04783_),
    .B1(_03457_),
    .B2(_05244_),
    .C(_03299_),
    .Y(_05245_));
 AO221x2_ASAP7_75t_R _12115_ (.A1(_05237_),
    .A2(_05240_),
    .B1(_05243_),
    .B2(_04881_),
    .C(_05245_),
    .Y(_05246_));
 NAND3x2_ASAP7_75t_R _12116_ (.B(_05234_),
    .C(_05246_),
    .Y(_05247_),
    .A(_04484_));
 NAND2x2_ASAP7_75t_R _12117_ (.A(_05224_),
    .B(_05247_),
    .Y(_09630_));
 INVx1_ASAP7_75t_R _12118_ (.A(_09630_),
    .Y(_09632_));
 BUFx10_ASAP7_75t_R _12119_ (.A(_03350_),
    .Y(_05248_));
 AO221x1_ASAP7_75t_R _12120_ (.A1(_04979_),
    .A2(_05195_),
    .B1(_05248_),
    .B2(_03345_),
    .C(_04977_),
    .Y(_05249_));
 NAND2x1_ASAP7_75t_R _12121_ (.A(_05092_),
    .B(_05197_),
    .Y(_05250_));
 OA21x2_ASAP7_75t_R _12122_ (.A1(_05092_),
    .A2(_05249_),
    .B(_05250_),
    .Y(_09748_));
 AND2x2_ASAP7_75t_R _12123_ (.A(_03578_),
    .B(_00556_),
    .Y(_05251_));
 AO21x1_ASAP7_75t_R _12124_ (.A1(_03573_),
    .A2(_00555_),
    .B(_05251_),
    .Y(_05252_));
 OR3x4_ASAP7_75t_R _12125_ (.A(_03052_),
    .B(net14),
    .C(_04492_),
    .Y(_05253_));
 AO21x1_ASAP7_75t_R _12126_ (.A1(_03107_),
    .A2(_05252_),
    .B(_05253_),
    .Y(_05254_));
 AND3x1_ASAP7_75t_R _12127_ (.A(_03048_),
    .B(_04503_),
    .C(_00554_),
    .Y(_05255_));
 OA21x2_ASAP7_75t_R _12128_ (.A1(_03625_),
    .A2(_03104_),
    .B(_00553_),
    .Y(_05256_));
 OA21x2_ASAP7_75t_R _12129_ (.A1(_05255_),
    .A2(_05256_),
    .B(_03604_),
    .Y(_05257_));
 AND2x2_ASAP7_75t_R _12130_ (.A(_03578_),
    .B(_00564_),
    .Y(_05258_));
 AO21x1_ASAP7_75t_R _12131_ (.A1(_03620_),
    .A2(_00563_),
    .B(_05258_),
    .Y(_05259_));
 OR3x4_ASAP7_75t_R _12132_ (.A(_03052_),
    .B(_03959_),
    .C(_04492_),
    .Y(_05260_));
 AO21x1_ASAP7_75t_R _12133_ (.A1(_03107_),
    .A2(_05259_),
    .B(_05260_),
    .Y(_05261_));
 AND3x1_ASAP7_75t_R _12134_ (.A(_04502_),
    .B(_04503_),
    .C(_00562_),
    .Y(_05262_));
 OA21x2_ASAP7_75t_R _12135_ (.A1(_03625_),
    .A2(_03104_),
    .B(_00561_),
    .Y(_05263_));
 OA21x2_ASAP7_75t_R _12136_ (.A1(_05262_),
    .A2(_05263_),
    .B(_03604_),
    .Y(_05264_));
 OA22x2_ASAP7_75t_R _12137_ (.A1(_05254_),
    .A2(_05257_),
    .B1(_05261_),
    .B2(_05264_),
    .Y(_05265_));
 BUFx6f_ASAP7_75t_R _12138_ (.A(_03040_),
    .Y(_05266_));
 AND2x2_ASAP7_75t_R _12139_ (.A(_03072_),
    .B(_00551_),
    .Y(_05267_));
 AO21x1_ASAP7_75t_R _12140_ (.A1(_03588_),
    .A2(_00549_),
    .B(_05267_),
    .Y(_05268_));
 NOR2x2_ASAP7_75t_R _12141_ (.A(_03085_),
    .B(_03103_),
    .Y(_05269_));
 AO221x1_ASAP7_75t_R _12142_ (.A1(_03086_),
    .A2(_00552_),
    .B1(_05269_),
    .B2(_00550_),
    .C(_03080_),
    .Y(_05270_));
 OA211x2_ASAP7_75t_R _12143_ (.A1(_05266_),
    .A2(_05268_),
    .B(_05270_),
    .C(_03585_),
    .Y(_05271_));
 BUFx6f_ASAP7_75t_R _12144_ (.A(_03040_),
    .Y(_05272_));
 AND2x2_ASAP7_75t_R _12145_ (.A(_03072_),
    .B(_00559_),
    .Y(_05273_));
 AO21x1_ASAP7_75t_R _12146_ (.A1(_03588_),
    .A2(_00557_),
    .B(_05273_),
    .Y(_05274_));
 AO221x1_ASAP7_75t_R _12147_ (.A1(_03086_),
    .A2(_00560_),
    .B1(_05269_),
    .B2(_00558_),
    .C(_03061_),
    .Y(_05275_));
 OA211x2_ASAP7_75t_R _12148_ (.A1(_05272_),
    .A2(_05274_),
    .B(_05275_),
    .C(_03118_),
    .Y(_05276_));
 OR3x1_ASAP7_75t_R _12149_ (.A(_03078_),
    .B(_05271_),
    .C(_05276_),
    .Y(_05277_));
 AOI21x1_ASAP7_75t_R _12150_ (.A1(_05265_),
    .A2(_05277_),
    .B(_03703_),
    .Y(_05278_));
 AO22x1_ASAP7_75t_R _12151_ (.A1(_05153_),
    .A2(_00533_),
    .B1(_00534_),
    .B2(_04361_),
    .Y(_05279_));
 AND2x2_ASAP7_75t_R _12152_ (.A(_03678_),
    .B(_00536_),
    .Y(_05280_));
 AO21x1_ASAP7_75t_R _12153_ (.A1(_03625_),
    .A2(_00535_),
    .B(_05280_),
    .Y(_05281_));
 AO21x1_ASAP7_75t_R _12154_ (.A1(_03689_),
    .A2(_05281_),
    .B(_04082_),
    .Y(_05282_));
 AND2x2_ASAP7_75t_R _12155_ (.A(_03097_),
    .B(_00533_),
    .Y(_05283_));
 AOI221x1_ASAP7_75t_R _12156_ (.A1(_03161_),
    .A2(_05279_),
    .B1(_05282_),
    .B2(_03215_),
    .C(_05283_),
    .Y(_05284_));
 AND2x2_ASAP7_75t_R _12157_ (.A(_03692_),
    .B(_00540_),
    .Y(_05285_));
 AO21x1_ASAP7_75t_R _12158_ (.A1(_03910_),
    .A2(_00539_),
    .B(_05285_),
    .Y(_05286_));
 AO21x1_ASAP7_75t_R _12159_ (.A1(_03689_),
    .A2(_05286_),
    .B(_03695_),
    .Y(_05287_));
 AND3x1_ASAP7_75t_R _12160_ (.A(_04499_),
    .B(_03020_),
    .C(_00538_),
    .Y(_05288_));
 OA21x2_ASAP7_75t_R _12161_ (.A1(_03111_),
    .A2(_03104_),
    .B(_00537_),
    .Y(_05289_));
 OA21x2_ASAP7_75t_R _12162_ (.A1(_05288_),
    .A2(_05289_),
    .B(_03604_),
    .Y(_05290_));
 OAI21x1_ASAP7_75t_R _12163_ (.A1(_05287_),
    .A2(_05290_),
    .B(_03586_),
    .Y(_05291_));
 NAND2x2_ASAP7_75t_R _12164_ (.A(_03080_),
    .B(_00541_),
    .Y(_05292_));
 INVx2_ASAP7_75t_R _12165_ (.A(_00542_),
    .Y(_05293_));
 OR3x1_ASAP7_75t_R _12166_ (.A(_03564_),
    .B(_03103_),
    .C(_05293_),
    .Y(_05294_));
 INVx3_ASAP7_75t_R _12167_ (.A(_00543_),
    .Y(_05295_));
 NAND2x1_ASAP7_75t_R _12168_ (.A(_03667_),
    .B(_00544_),
    .Y(_05296_));
 OA211x2_ASAP7_75t_R _12169_ (.A1(_03047_),
    .A2(_05295_),
    .B(_05296_),
    .C(_03085_),
    .Y(_05297_));
 AO31x2_ASAP7_75t_R _12170_ (.A1(_03027_),
    .A2(_05292_),
    .A3(_05294_),
    .B(_05297_),
    .Y(_05298_));
 AND2x2_ASAP7_75t_R _12171_ (.A(_03057_),
    .B(_00548_),
    .Y(_05299_));
 AO21x1_ASAP7_75t_R _12172_ (.A1(_03055_),
    .A2(_00547_),
    .B(_05299_),
    .Y(_05300_));
 AOI21x1_ASAP7_75t_R _12173_ (.A1(_03087_),
    .A2(_05300_),
    .B(_03617_),
    .Y(_05301_));
 AND3x1_ASAP7_75t_R _12174_ (.A(_04267_),
    .B(_03044_),
    .C(_00546_),
    .Y(_05302_));
 OA21x2_ASAP7_75t_R _12175_ (.A1(_03055_),
    .A2(_03096_),
    .B(_00545_),
    .Y(_05303_));
 OAI21x1_ASAP7_75t_R _12176_ (.A1(_05302_),
    .A2(_05303_),
    .B(_03635_),
    .Y(_05304_));
 AO221x1_ASAP7_75t_R _12177_ (.A1(_03052_),
    .A2(_05298_),
    .B1(_05301_),
    .B2(_05304_),
    .C(_03585_),
    .Y(_05305_));
 OA211x2_ASAP7_75t_R _12178_ (.A1(_05284_),
    .A2(_05291_),
    .B(_05305_),
    .C(_03154_),
    .Y(_05306_));
 OA21x2_ASAP7_75t_R _12179_ (.A1(_05278_),
    .A2(_05306_),
    .B(_03705_),
    .Y(_05307_));
 AND2x2_ASAP7_75t_R _12180_ (.A(_04422_),
    .B(_05307_),
    .Y(_05308_));
 AOI21x1_ASAP7_75t_R _12181_ (.A1(_03645_),
    .A2(_09748_),
    .B(_05308_),
    .Y(_05309_));
 XNOR2x1_ASAP7_75t_R _12182_ (.B(_05309_),
    .Y(_09636_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _12183_ (.A(_09636_),
    .Y(_09638_));
 OA22x2_ASAP7_75t_R _12184_ (.A1(_00551_),
    .A2(_03350_),
    .B1(_03357_),
    .B2(_00552_),
    .Y(_05310_));
 AND3x1_ASAP7_75t_R _12185_ (.A(_03149_),
    .B(_03475_),
    .C(_00556_),
    .Y(_05311_));
 AO221x1_ASAP7_75t_R _12186_ (.A1(_03317_),
    .A2(_04020_),
    .B1(_03976_),
    .B2(_00555_),
    .C(_05311_),
    .Y(_05312_));
 OA211x2_ASAP7_75t_R _12187_ (.A1(_05127_),
    .A2(_05310_),
    .B(_05312_),
    .C(_04771_),
    .Y(_05313_));
 BUFx6f_ASAP7_75t_R _12188_ (.A(_03359_),
    .Y(_05314_));
 OA22x2_ASAP7_75t_R _12189_ (.A1(_00553_),
    .A2(_03350_),
    .B1(_03357_),
    .B2(_00554_),
    .Y(_05315_));
 OA211x2_ASAP7_75t_R _12190_ (.A1(_03226_),
    .A2(_03311_),
    .B(_03994_),
    .C(_00550_),
    .Y(_05316_));
 AO21x1_ASAP7_75t_R _12191_ (.A1(_00549_),
    .A2(_03415_),
    .B(_05316_),
    .Y(_05317_));
 BUFx12_ASAP7_75t_R _12192_ (.A(_03393_),
    .Y(_05318_));
 AO221x1_ASAP7_75t_R _12193_ (.A1(_05314_),
    .A2(_05315_),
    .B1(_05317_),
    .B2(_05318_),
    .C(_03341_),
    .Y(_05319_));
 OA21x2_ASAP7_75t_R _12194_ (.A1(_04458_),
    .A2(_05313_),
    .B(_05319_),
    .Y(_05320_));
 OA22x2_ASAP7_75t_R _12195_ (.A1(_00562_),
    .A2(_03377_),
    .B1(_04768_),
    .B2(_00561_),
    .Y(_05321_));
 OA211x2_ASAP7_75t_R _12196_ (.A1(_03226_),
    .A2(_03311_),
    .B(_03349_),
    .C(_00558_),
    .Y(_05322_));
 AO21x1_ASAP7_75t_R _12197_ (.A1(_00557_),
    .A2(_03383_),
    .B(_05322_),
    .Y(_05323_));
 OA21x2_ASAP7_75t_R _12198_ (.A1(_03411_),
    .A2(_05323_),
    .B(_04899_),
    .Y(_05324_));
 OR3x1_ASAP7_75t_R _12199_ (.A(_03096_),
    .B(_04561_),
    .C(_00560_),
    .Y(_05325_));
 AO21x1_ASAP7_75t_R _12200_ (.A1(_03351_),
    .A2(_03352_),
    .B(_05325_),
    .Y(_05326_));
 OA21x2_ASAP7_75t_R _12201_ (.A1(_00559_),
    .A2(_03329_),
    .B(_03388_),
    .Y(_05327_));
 AO21x1_ASAP7_75t_R _12202_ (.A1(_05326_),
    .A2(_05327_),
    .B(_03988_),
    .Y(_05328_));
 AND3x1_ASAP7_75t_R _12203_ (.A(_03045_),
    .B(_05124_),
    .C(_00564_),
    .Y(_05329_));
 AO21x1_ASAP7_75t_R _12204_ (.A1(_00563_),
    .A2(_03397_),
    .B(_05329_),
    .Y(_05330_));
 AO22x1_ASAP7_75t_R _12205_ (.A1(_03210_),
    .A2(_05328_),
    .B1(_05330_),
    .B2(_04885_),
    .Y(_05331_));
 OA211x2_ASAP7_75t_R _12206_ (.A1(_04107_),
    .A2(_05321_),
    .B(_05324_),
    .C(_05331_),
    .Y(_05332_));
 NOR3x2_ASAP7_75t_R _12207_ (.B(_05320_),
    .C(_05332_),
    .Y(_05333_),
    .A(_04003_));
 OA22x2_ASAP7_75t_R _12208_ (.A1(_00540_),
    .A2(_03732_),
    .B1(_03733_),
    .B2(_00536_),
    .Y(_05334_));
 BUFx10_ASAP7_75t_R _12209_ (.A(_03475_),
    .Y(_05335_));
 AND3x1_ASAP7_75t_R _12210_ (.A(_00535_),
    .B(_03326_),
    .C(_03322_),
    .Y(_05336_));
 AO221x1_ASAP7_75t_R _12211_ (.A1(_03022_),
    .A2(_05335_),
    .B1(_00539_),
    .B2(_05127_),
    .C(_05336_),
    .Y(_05337_));
 AO21x2_ASAP7_75t_R _12212_ (.A1(_05334_),
    .A2(_05337_),
    .B(_04214_),
    .Y(_05338_));
 INVx1_ASAP7_75t_R _12213_ (.A(_00533_),
    .Y(_01229_));
 NAND2x1_ASAP7_75t_R _12214_ (.A(_00534_),
    .B(_04768_),
    .Y(_05339_));
 OA21x2_ASAP7_75t_R _12215_ (.A1(_01229_),
    .A2(_03410_),
    .B(_05339_),
    .Y(_05340_));
 BUFx12_ASAP7_75t_R _12216_ (.A(_04472_),
    .Y(_05341_));
 OAI22x1_ASAP7_75t_R _12217_ (.A1(_00537_),
    .A2(_05248_),
    .B1(_05341_),
    .B2(_00538_),
    .Y(_05342_));
 AOI221x1_ASAP7_75t_R _12218_ (.A1(_04881_),
    .A2(_05340_),
    .B1(_05342_),
    .B2(_04549_),
    .C(_04791_),
    .Y(_05343_));
 OA22x2_ASAP7_75t_R _12219_ (.A1(_00546_),
    .A2(_04550_),
    .B1(_03410_),
    .B2(_00545_),
    .Y(_05344_));
 INVx1_ASAP7_75t_R _12220_ (.A(_00541_),
    .Y(_05345_));
 OA211x2_ASAP7_75t_R _12221_ (.A1(_03226_),
    .A2(_03311_),
    .B(_03735_),
    .C(_05293_),
    .Y(_05346_));
 AO21x1_ASAP7_75t_R _12222_ (.A1(_05345_),
    .A2(_04472_),
    .B(_05346_),
    .Y(_05347_));
 AOI221x1_ASAP7_75t_R _12223_ (.A1(_04784_),
    .A2(_04783_),
    .B1(_03484_),
    .B2(_05347_),
    .C(_03300_),
    .Y(_05348_));
 INVx1_ASAP7_75t_R _12224_ (.A(_00544_),
    .Y(_05349_));
 OA211x2_ASAP7_75t_R _12225_ (.A1(_03226_),
    .A2(_03311_),
    .B(_03385_),
    .C(_05349_),
    .Y(_05350_));
 AO21x1_ASAP7_75t_R _12226_ (.A1(_05295_),
    .A2(_03437_),
    .B(_05314_),
    .Y(_05351_));
 OA21x2_ASAP7_75t_R _12227_ (.A1(_05350_),
    .A2(_05351_),
    .B(_03382_),
    .Y(_05352_));
 AND3x1_ASAP7_75t_R _12228_ (.A(_03021_),
    .B(_05335_),
    .C(_00548_),
    .Y(_05353_));
 AOI21x1_ASAP7_75t_R _12229_ (.A1(_00547_),
    .A2(_03377_),
    .B(_05353_),
    .Y(_05354_));
 OAI22x1_ASAP7_75t_R _12230_ (.A1(_03278_),
    .A2(_05352_),
    .B1(_05354_),
    .B2(_05318_),
    .Y(_05355_));
 OA211x2_ASAP7_75t_R _12231_ (.A1(_04107_),
    .A2(_05344_),
    .B(_05348_),
    .C(_05355_),
    .Y(_05356_));
 AOI211x1_ASAP7_75t_R _12232_ (.A1(_05338_),
    .A2(_05343_),
    .B(_05356_),
    .C(_03426_),
    .Y(_05357_));
 NOR2x2_ASAP7_75t_R _12233_ (.A(_05333_),
    .B(_05357_),
    .Y(_09637_));
 BUFx6f_ASAP7_75t_R _12234_ (.A(net6),
    .Y(_05358_));
 AND3x1_ASAP7_75t_R _12235_ (.A(net89),
    .B(_05358_),
    .C(_04985_),
    .Y(_05359_));
 AO21x1_ASAP7_75t_R _12236_ (.A1(_05248_),
    .A2(_04984_),
    .B(_05359_),
    .Y(_05360_));
 OR2x2_ASAP7_75t_R _12237_ (.A(_05248_),
    .B(_04984_),
    .Y(_05361_));
 OA211x2_ASAP7_75t_R _12238_ (.A1(_05195_),
    .A2(_04985_),
    .B(_05361_),
    .C(_04979_),
    .Y(_05362_));
 AO21x1_ASAP7_75t_R _12239_ (.A1(_03345_),
    .A2(_05360_),
    .B(_05362_),
    .Y(_05363_));
 OA21x2_ASAP7_75t_R _12240_ (.A1(_04977_),
    .A2(_05363_),
    .B(_04981_),
    .Y(_09746_));
 BUFx6f_ASAP7_75t_R _12241_ (.A(_04487_),
    .Y(_05364_));
 BUFx6f_ASAP7_75t_R _12242_ (.A(_05364_),
    .Y(_05365_));
 BUFx6f_ASAP7_75t_R _12243_ (.A(_05070_),
    .Y(_05366_));
 AND2x2_ASAP7_75t_R _12244_ (.A(_05366_),
    .B(_00569_),
    .Y(_05367_));
 AO21x1_ASAP7_75t_R _12245_ (.A1(_05064_),
    .A2(_00568_),
    .B(_05367_),
    .Y(_05368_));
 AO21x1_ASAP7_75t_R _12246_ (.A1(_05365_),
    .A2(_05368_),
    .B(_05067_),
    .Y(_05369_));
 BUFx6f_ASAP7_75t_R _12247_ (.A(_04361_),
    .Y(_05370_));
 AO22x1_ASAP7_75t_R _12248_ (.A1(_05064_),
    .A2(_00566_),
    .B1(_00567_),
    .B2(_05370_),
    .Y(_05371_));
 BUFx6f_ASAP7_75t_R _12249_ (.A(_04381_),
    .Y(_05372_));
 AO22x1_ASAP7_75t_R _12250_ (.A1(_03099_),
    .A2(_00566_),
    .B1(_05371_),
    .B2(_05372_),
    .Y(_05373_));
 AO21x1_ASAP7_75t_R _12251_ (.A1(_03023_),
    .A2(_05369_),
    .B(_05373_),
    .Y(_05374_));
 BUFx6f_ASAP7_75t_R _12252_ (.A(_04401_),
    .Y(_05375_));
 BUFx6f_ASAP7_75t_R _12253_ (.A(_03071_),
    .Y(_05376_));
 AND2x2_ASAP7_75t_R _12254_ (.A(_05376_),
    .B(_00573_),
    .Y(_05377_));
 AO21x1_ASAP7_75t_R _12255_ (.A1(_05375_),
    .A2(_00572_),
    .B(_05377_),
    .Y(_05378_));
 AND3x1_ASAP7_75t_R _12256_ (.A(_05376_),
    .B(_03022_),
    .C(_00571_),
    .Y(_05379_));
 AO21x1_ASAP7_75t_R _12257_ (.A1(_00570_),
    .A2(_03291_),
    .B(_05379_),
    .Y(_05380_));
 AO221x1_ASAP7_75t_R _12258_ (.A1(_05365_),
    .A2(_05378_),
    .B1(_05380_),
    .B2(_04764_),
    .C(_04657_),
    .Y(_05381_));
 AND3x1_ASAP7_75t_R _12259_ (.A(_04545_),
    .B(_05374_),
    .C(_05381_),
    .Y(_05382_));
 AND2x2_ASAP7_75t_R _12260_ (.A(_05376_),
    .B(_00581_),
    .Y(_05383_));
 AO21x1_ASAP7_75t_R _12261_ (.A1(_05375_),
    .A2(_00580_),
    .B(_05383_),
    .Y(_05384_));
 AND3x1_ASAP7_75t_R _12262_ (.A(_05376_),
    .B(_03022_),
    .C(_00579_),
    .Y(_05385_));
 AO21x1_ASAP7_75t_R _12263_ (.A1(_00578_),
    .A2(_03291_),
    .B(_05385_),
    .Y(_05386_));
 AO221x1_ASAP7_75t_R _12264_ (.A1(_05365_),
    .A2(_05384_),
    .B1(_05386_),
    .B2(_04764_),
    .C(_04657_),
    .Y(_05387_));
 AO22x1_ASAP7_75t_R _12265_ (.A1(_05375_),
    .A2(_00574_),
    .B1(_00575_),
    .B2(_05370_),
    .Y(_05388_));
 AND2x2_ASAP7_75t_R _12266_ (.A(_05366_),
    .B(_00577_),
    .Y(_05389_));
 AO21x1_ASAP7_75t_R _12267_ (.A1(_05064_),
    .A2(_00576_),
    .B(_05389_),
    .Y(_05390_));
 AO21x1_ASAP7_75t_R _12268_ (.A1(_05365_),
    .A2(_05390_),
    .B(_05067_),
    .Y(_05391_));
 AO21x1_ASAP7_75t_R _12269_ (.A1(_05372_),
    .A2(_05388_),
    .B(_05391_),
    .Y(_05392_));
 AND3x1_ASAP7_75t_R _12270_ (.A(_03175_),
    .B(_05387_),
    .C(_05392_),
    .Y(_05393_));
 OR3x1_ASAP7_75t_R _12271_ (.A(_04486_),
    .B(_05382_),
    .C(_05393_),
    .Y(_05394_));
 AND2x2_ASAP7_75t_R _12272_ (.A(_05376_),
    .B(_00597_),
    .Y(_05395_));
 AO21x1_ASAP7_75t_R _12273_ (.A1(_05375_),
    .A2(_00596_),
    .B(_05395_),
    .Y(_05396_));
 AND3x1_ASAP7_75t_R _12274_ (.A(_05376_),
    .B(_03022_),
    .C(_00595_),
    .Y(_05397_));
 AO21x1_ASAP7_75t_R _12275_ (.A1(_00594_),
    .A2(_03291_),
    .B(_05397_),
    .Y(_05398_));
 AO221x1_ASAP7_75t_R _12276_ (.A1(_05365_),
    .A2(_05396_),
    .B1(_05398_),
    .B2(_04764_),
    .C(_04657_),
    .Y(_05399_));
 AND2x2_ASAP7_75t_R _12277_ (.A(_05364_),
    .B(_00592_),
    .Y(_05400_));
 AO21x1_ASAP7_75t_R _12278_ (.A1(_05372_),
    .A2(_00590_),
    .B(_05400_),
    .Y(_05401_));
 AO21x1_ASAP7_75t_R _12279_ (.A1(_00591_),
    .A2(_05066_),
    .B(_05067_),
    .Y(_05402_));
 AO221x1_ASAP7_75t_R _12280_ (.A1(_00593_),
    .A2(_05061_),
    .B1(_05401_),
    .B2(_05375_),
    .C(_05402_),
    .Y(_05403_));
 AND3x1_ASAP7_75t_R _12281_ (.A(_03175_),
    .B(_05399_),
    .C(_05403_),
    .Y(_05404_));
 AND2x2_ASAP7_75t_R _12282_ (.A(_05376_),
    .B(_00589_),
    .Y(_05405_));
 AO21x1_ASAP7_75t_R _12283_ (.A1(_05375_),
    .A2(_00588_),
    .B(_05405_),
    .Y(_05406_));
 AND3x1_ASAP7_75t_R _12284_ (.A(_05376_),
    .B(_03022_),
    .C(_00587_),
    .Y(_05407_));
 AO21x1_ASAP7_75t_R _12285_ (.A1(_00586_),
    .A2(_03291_),
    .B(_05407_),
    .Y(_05408_));
 AO221x1_ASAP7_75t_R _12286_ (.A1(_05365_),
    .A2(_05406_),
    .B1(_05408_),
    .B2(_04764_),
    .C(_04657_),
    .Y(_05409_));
 BUFx6f_ASAP7_75t_R _12287_ (.A(_03107_),
    .Y(_05410_));
 AND2x2_ASAP7_75t_R _12288_ (.A(_05410_),
    .B(_00584_),
    .Y(_05411_));
 AO21x1_ASAP7_75t_R _12289_ (.A1(_05372_),
    .A2(_00582_),
    .B(_05411_),
    .Y(_05412_));
 AO21x1_ASAP7_75t_R _12290_ (.A1(_00583_),
    .A2(_05066_),
    .B(_05067_),
    .Y(_05413_));
 AO221x1_ASAP7_75t_R _12291_ (.A1(_00585_),
    .A2(_05061_),
    .B1(_05412_),
    .B2(_05375_),
    .C(_05413_),
    .Y(_05414_));
 AND3x1_ASAP7_75t_R _12292_ (.A(_04545_),
    .B(_05409_),
    .C(_05414_),
    .Y(_05415_));
 OR3x1_ASAP7_75t_R _12293_ (.A(_04423_),
    .B(_05404_),
    .C(_05415_),
    .Y(_05416_));
 AOI21x1_ASAP7_75t_R _12294_ (.A1(_05394_),
    .A2(_05416_),
    .B(_04163_),
    .Y(_05417_));
 AND2x2_ASAP7_75t_R _12295_ (.A(_04422_),
    .B(_05417_),
    .Y(_05418_));
 AOI21x1_ASAP7_75t_R _12296_ (.A1(_03645_),
    .A2(_09746_),
    .B(_05418_),
    .Y(_05419_));
 XNOR2x1_ASAP7_75t_R _12297_ (.B(_05419_),
    .Y(_09641_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _12298_ (.A(_09641_),
    .Y(_09643_));
 OAI22x1_ASAP7_75t_R _12299_ (.A1(_00592_),
    .A2(_03429_),
    .B1(_03529_),
    .B2(_00593_),
    .Y(_05420_));
 NAND2x1_ASAP7_75t_R _12300_ (.A(_03444_),
    .B(_05420_),
    .Y(_05421_));
 AND2x2_ASAP7_75t_R _12301_ (.A(_00590_),
    .B(_04153_),
    .Y(_05422_));
 AO221x1_ASAP7_75t_R _12302_ (.A1(_03245_),
    .A2(_03340_),
    .B1(_04132_),
    .B2(_00591_),
    .C(_05422_),
    .Y(_05423_));
 AND3x1_ASAP7_75t_R _12303_ (.A(_03317_),
    .B(_03997_),
    .C(_03322_),
    .Y(_05424_));
 OA22x2_ASAP7_75t_R _12304_ (.A1(_00586_),
    .A2(_03349_),
    .B1(_03418_),
    .B2(_00587_),
    .Y(_05425_));
 OA22x2_ASAP7_75t_R _12305_ (.A1(_00588_),
    .A2(_03348_),
    .B1(_03355_),
    .B2(_00589_),
    .Y(_05426_));
 OA211x2_ASAP7_75t_R _12306_ (.A1(_03273_),
    .A2(_03287_),
    .B(_03501_),
    .C(_05426_),
    .Y(_05427_));
 AO21x1_ASAP7_75t_R _12307_ (.A1(_04214_),
    .A2(_05425_),
    .B(_05427_),
    .Y(_05428_));
 AND2x2_ASAP7_75t_R _12308_ (.A(_03550_),
    .B(_04444_),
    .Y(_05429_));
 AO32x1_ASAP7_75t_R _12309_ (.A1(_05421_),
    .A2(_05423_),
    .A3(_05424_),
    .B1(_05428_),
    .B2(_05429_),
    .Y(_05430_));
 OA22x2_ASAP7_75t_R _12310_ (.A1(_00584_),
    .A2(_03306_),
    .B1(_03486_),
    .B2(_00585_),
    .Y(_05431_));
 AND3x1_ASAP7_75t_R _12311_ (.A(_03299_),
    .B(_03394_),
    .C(_05431_),
    .Y(_05432_));
 AND2x2_ASAP7_75t_R _12312_ (.A(_00583_),
    .B(_03467_),
    .Y(_05433_));
 AO21x1_ASAP7_75t_R _12313_ (.A1(_00582_),
    .A2(_03529_),
    .B(_05433_),
    .Y(_05434_));
 AO21x1_ASAP7_75t_R _12314_ (.A1(_03421_),
    .A2(_05434_),
    .B(_03862_),
    .Y(_05435_));
 AO21x1_ASAP7_75t_R _12315_ (.A1(_03444_),
    .A2(_05432_),
    .B(_05435_),
    .Y(_05436_));
 OR2x2_ASAP7_75t_R _12316_ (.A(_00597_),
    .B(_03431_),
    .Y(_05437_));
 OA211x2_ASAP7_75t_R _12317_ (.A1(_00596_),
    .A2(_05106_),
    .B(_03443_),
    .C(_05437_),
    .Y(_05438_));
 OA222x2_ASAP7_75t_R _12318_ (.A1(_03344_),
    .A2(_03855_),
    .B1(_03976_),
    .B2(_00595_),
    .C1(_00594_),
    .C2(_03409_),
    .Y(_05439_));
 OA21x2_ASAP7_75t_R _12319_ (.A1(_03273_),
    .A2(_03287_),
    .B(_03747_),
    .Y(_05440_));
 OA211x2_ASAP7_75t_R _12320_ (.A1(_05438_),
    .A2(_05439_),
    .B(_05440_),
    .C(_03888_),
    .Y(_05441_));
 AOI211x1_ASAP7_75t_R _12321_ (.A1(_03247_),
    .A2(_05430_),
    .B(_05436_),
    .C(_05441_),
    .Y(_05442_));
 AO21x2_ASAP7_75t_R _12322_ (.A1(_03233_),
    .A2(_03243_),
    .B(_03393_),
    .Y(_05443_));
 BUFx4f_ASAP7_75t_R _12323_ (.A(_05443_),
    .Y(_05444_));
 OA22x2_ASAP7_75t_R _12324_ (.A1(_00576_),
    .A2(_03735_),
    .B1(_03740_),
    .B2(_00577_),
    .Y(_05445_));
 OA22x2_ASAP7_75t_R _12325_ (.A1(_00580_),
    .A2(_03522_),
    .B1(_03485_),
    .B2(_00581_),
    .Y(_05446_));
 OA211x2_ASAP7_75t_R _12326_ (.A1(_03273_),
    .A2(_03287_),
    .B(_03440_),
    .C(_05446_),
    .Y(_05447_));
 AO21x1_ASAP7_75t_R _12327_ (.A1(_05444_),
    .A2(_05445_),
    .B(_05447_),
    .Y(_05448_));
 AND2x2_ASAP7_75t_R _12328_ (.A(_00575_),
    .B(_03400_),
    .Y(_05449_));
 AOI21x1_ASAP7_75t_R _12329_ (.A1(_00574_),
    .A2(_04473_),
    .B(_05449_),
    .Y(_05450_));
 OAI22x1_ASAP7_75t_R _12330_ (.A1(_00579_),
    .A2(_03847_),
    .B1(_03408_),
    .B2(_00578_),
    .Y(_05451_));
 OA211x2_ASAP7_75t_R _12331_ (.A1(_03273_),
    .A2(_03287_),
    .B(_03504_),
    .C(_05451_),
    .Y(_05452_));
 AOI211x1_ASAP7_75t_R _12332_ (.A1(_05444_),
    .A2(_05450_),
    .B(_05452_),
    .C(_03444_),
    .Y(_05453_));
 AO21x1_ASAP7_75t_R _12333_ (.A1(_03444_),
    .A2(_05448_),
    .B(_05453_),
    .Y(_05454_));
 OA22x2_ASAP7_75t_R _12334_ (.A1(_00568_),
    .A2(_03385_),
    .B1(_03740_),
    .B2(_00569_),
    .Y(_05455_));
 OA22x2_ASAP7_75t_R _12335_ (.A1(_00572_),
    .A2(_03328_),
    .B1(_03413_),
    .B2(_00573_),
    .Y(_05456_));
 OA211x2_ASAP7_75t_R _12336_ (.A1(_03273_),
    .A2(_03287_),
    .B(_03440_),
    .C(_05456_),
    .Y(_05457_));
 AO21x1_ASAP7_75t_R _12337_ (.A1(_05443_),
    .A2(_05455_),
    .B(_05457_),
    .Y(_05458_));
 AND2x2_ASAP7_75t_R _12338_ (.A(_00567_),
    .B(_03453_),
    .Y(_05459_));
 AO21x1_ASAP7_75t_R _12339_ (.A1(_00566_),
    .A2(_03418_),
    .B(_05459_),
    .Y(_05460_));
 OA22x2_ASAP7_75t_R _12340_ (.A1(_00570_),
    .A2(_03837_),
    .B1(_03430_),
    .B2(_00571_),
    .Y(_05461_));
 OA211x2_ASAP7_75t_R _12341_ (.A1(_03272_),
    .A2(_03287_),
    .B(_03440_),
    .C(_05461_),
    .Y(_05462_));
 AO221x1_ASAP7_75t_R _12342_ (.A1(_03245_),
    .A2(_03502_),
    .B1(_05443_),
    .B2(_05460_),
    .C(_05462_),
    .Y(_05463_));
 OA211x2_ASAP7_75t_R _12343_ (.A1(_04214_),
    .A2(_05458_),
    .B(_05463_),
    .C(_04552_),
    .Y(_05464_));
 AOI211x1_ASAP7_75t_R _12344_ (.A1(_04791_),
    .A2(_05454_),
    .B(_05464_),
    .C(_03426_),
    .Y(_05465_));
 OR2x2_ASAP7_75t_R _12345_ (.A(_05442_),
    .B(_05465_),
    .Y(_05466_));
 BUFx2_ASAP7_75t_R _12346_ (.A(_05466_),
    .Y(_09640_));
 INVx2_ASAP7_75t_R _12347_ (.A(_09640_),
    .Y(_09642_));
 AO21x2_ASAP7_75t_R _12348_ (.A1(_03240_),
    .A2(_04978_),
    .B(_03278_),
    .Y(_05467_));
 AND2x4_ASAP7_75t_R _12349_ (.A(_03023_),
    .B(_03212_),
    .Y(_05468_));
 AND3x1_ASAP7_75t_R _12350_ (.A(_03025_),
    .B(_05358_),
    .C(_04984_),
    .Y(_05469_));
 AO21x1_ASAP7_75t_R _12351_ (.A1(_04985_),
    .A2(_05468_),
    .B(_05469_),
    .Y(_05470_));
 AO32x1_ASAP7_75t_R _12352_ (.A1(_03267_),
    .A2(_05467_),
    .A3(_05360_),
    .B1(_05470_),
    .B2(_03345_),
    .Y(_05471_));
 OA21x2_ASAP7_75t_R _12353_ (.A1(_04977_),
    .A2(_05471_),
    .B(_04981_),
    .Y(_09744_));
 AND2x2_ASAP7_75t_R _12354_ (.A(_05070_),
    .B(_00603_),
    .Y(_05472_));
 AO21x1_ASAP7_75t_R _12355_ (.A1(_04528_),
    .A2(_00602_),
    .B(_05472_),
    .Y(_05473_));
 BUFx6f_ASAP7_75t_R _12356_ (.A(_03623_),
    .Y(_05474_));
 AO21x1_ASAP7_75t_R _12357_ (.A1(_05364_),
    .A2(_05473_),
    .B(_05474_),
    .Y(_05475_));
 AO22x1_ASAP7_75t_R _12358_ (.A1(_04748_),
    .A2(_00600_),
    .B1(_00601_),
    .B2(_04513_),
    .Y(_05476_));
 AO22x1_ASAP7_75t_R _12359_ (.A1(_03131_),
    .A2(_00600_),
    .B1(_05476_),
    .B2(_03029_),
    .Y(_05477_));
 AO21x1_ASAP7_75t_R _12360_ (.A1(_03023_),
    .A2(_05475_),
    .B(_05477_),
    .Y(_05478_));
 AND2x2_ASAP7_75t_R _12361_ (.A(_03041_),
    .B(_00607_),
    .Y(_05479_));
 AO21x1_ASAP7_75t_R _12362_ (.A1(_04401_),
    .A2(_00606_),
    .B(_05479_),
    .Y(_05480_));
 AND3x1_ASAP7_75t_R _12363_ (.A(_03071_),
    .B(_03021_),
    .C(_00605_),
    .Y(_05481_));
 AO21x1_ASAP7_75t_R _12364_ (.A1(_00604_),
    .A2(_05073_),
    .B(_05481_),
    .Y(_05482_));
 AO221x1_ASAP7_75t_R _12365_ (.A1(_05069_),
    .A2(_05480_),
    .B1(_05482_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_05483_));
 AND3x1_ASAP7_75t_R _12366_ (.A(_04545_),
    .B(_05478_),
    .C(_05483_),
    .Y(_05484_));
 AND2x2_ASAP7_75t_R _12367_ (.A(_03041_),
    .B(_00615_),
    .Y(_05485_));
 AO21x1_ASAP7_75t_R _12368_ (.A1(_04401_),
    .A2(_00614_),
    .B(_05485_),
    .Y(_05486_));
 AND3x1_ASAP7_75t_R _12369_ (.A(_03071_),
    .B(_03021_),
    .C(_00613_),
    .Y(_05487_));
 AO21x1_ASAP7_75t_R _12370_ (.A1(_00612_),
    .A2(_05073_),
    .B(_05487_),
    .Y(_05488_));
 AO221x1_ASAP7_75t_R _12371_ (.A1(_05069_),
    .A2(_05486_),
    .B1(_05488_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_05489_));
 AO22x1_ASAP7_75t_R _12372_ (.A1(_04860_),
    .A2(_00608_),
    .B1(_00609_),
    .B2(_05370_),
    .Y(_05490_));
 AND2x2_ASAP7_75t_R _12373_ (.A(_05070_),
    .B(_00611_),
    .Y(_05491_));
 AO21x1_ASAP7_75t_R _12374_ (.A1(_04528_),
    .A2(_00610_),
    .B(_05491_),
    .Y(_05492_));
 AO21x1_ASAP7_75t_R _12375_ (.A1(_05364_),
    .A2(_05492_),
    .B(_05474_),
    .Y(_05493_));
 AO21x1_ASAP7_75t_R _12376_ (.A1(_05372_),
    .A2(_05490_),
    .B(_05493_),
    .Y(_05494_));
 AND3x1_ASAP7_75t_R _12377_ (.A(_03175_),
    .B(_05489_),
    .C(_05494_),
    .Y(_05495_));
 OR3x1_ASAP7_75t_R _12378_ (.A(_04486_),
    .B(_05484_),
    .C(_05495_),
    .Y(_05496_));
 AND2x2_ASAP7_75t_R _12379_ (.A(_03071_),
    .B(_00631_),
    .Y(_05497_));
 AO21x1_ASAP7_75t_R _12380_ (.A1(_04860_),
    .A2(_00630_),
    .B(_05497_),
    .Y(_05498_));
 AND3x1_ASAP7_75t_R _12381_ (.A(_03071_),
    .B(_05229_),
    .C(_00629_),
    .Y(_05499_));
 AO21x1_ASAP7_75t_R _12382_ (.A1(_00628_),
    .A2(_05073_),
    .B(_05499_),
    .Y(_05500_));
 AO221x1_ASAP7_75t_R _12383_ (.A1(_05069_),
    .A2(_05498_),
    .B1(_05500_),
    .B2(_05076_),
    .C(_04657_),
    .Y(_05501_));
 AND2x2_ASAP7_75t_R _12384_ (.A(_03074_),
    .B(_00626_),
    .Y(_05502_));
 AO21x1_ASAP7_75t_R _12385_ (.A1(_03029_),
    .A2(_00624_),
    .B(_05502_),
    .Y(_05503_));
 AO21x1_ASAP7_75t_R _12386_ (.A1(_00625_),
    .A2(_05066_),
    .B(_05474_),
    .Y(_05504_));
 AO221x1_ASAP7_75t_R _12387_ (.A1(_00627_),
    .A2(_05061_),
    .B1(_05503_),
    .B2(_05064_),
    .C(_05504_),
    .Y(_05505_));
 AND3x1_ASAP7_75t_R _12388_ (.A(_03175_),
    .B(_05501_),
    .C(_05505_),
    .Y(_05506_));
 AND2x2_ASAP7_75t_R _12389_ (.A(_03071_),
    .B(_00623_),
    .Y(_05507_));
 AO21x1_ASAP7_75t_R _12390_ (.A1(_04860_),
    .A2(_00622_),
    .B(_05507_),
    .Y(_05508_));
 AND3x1_ASAP7_75t_R _12391_ (.A(_03071_),
    .B(_05229_),
    .C(_00621_),
    .Y(_05509_));
 AO21x1_ASAP7_75t_R _12392_ (.A1(_00620_),
    .A2(_05073_),
    .B(_05509_),
    .Y(_05510_));
 AO221x1_ASAP7_75t_R _12393_ (.A1(_05069_),
    .A2(_05508_),
    .B1(_05510_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_05511_));
 AND2x2_ASAP7_75t_R _12394_ (.A(_03074_),
    .B(_00618_),
    .Y(_05512_));
 AO21x1_ASAP7_75t_R _12395_ (.A1(_03904_),
    .A2(_00616_),
    .B(_05512_),
    .Y(_05513_));
 AO21x1_ASAP7_75t_R _12396_ (.A1(_00617_),
    .A2(_05066_),
    .B(_05474_),
    .Y(_05514_));
 AO221x1_ASAP7_75t_R _12397_ (.A1(_00619_),
    .A2(_05061_),
    .B1(_05513_),
    .B2(_05064_),
    .C(_05514_),
    .Y(_05515_));
 AND3x1_ASAP7_75t_R _12398_ (.A(_04545_),
    .B(_05511_),
    .C(_05515_),
    .Y(_05516_));
 OR3x1_ASAP7_75t_R _12399_ (.A(_04423_),
    .B(_05506_),
    .C(_05516_),
    .Y(_05517_));
 AOI21x1_ASAP7_75t_R _12400_ (.A1(_05496_),
    .A2(_05517_),
    .B(_04163_),
    .Y(_05518_));
 AND2x2_ASAP7_75t_R _12401_ (.A(_04422_),
    .B(_05518_),
    .Y(_05519_));
 AOI21x1_ASAP7_75t_R _12402_ (.A1(_03645_),
    .A2(_09744_),
    .B(_05519_),
    .Y(_05520_));
 XNOR2x1_ASAP7_75t_R _12403_ (.B(_05520_),
    .Y(_09646_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _12404_ (.A(_09646_),
    .Y(_09648_));
 OA211x2_ASAP7_75t_R _12405_ (.A1(_03284_),
    .A2(_03288_),
    .B(_03472_),
    .C(_00628_),
    .Y(_05521_));
 AO221x1_ASAP7_75t_R _12406_ (.A1(_05248_),
    .A2(_03759_),
    .B1(_05444_),
    .B2(_00624_),
    .C(_05521_),
    .Y(_05522_));
 NOR2x1_ASAP7_75t_R _12407_ (.A(_00625_),
    .B(_05341_),
    .Y(_05523_));
 NOR2x1_ASAP7_75t_R _12408_ (.A(_00629_),
    .B(_03378_),
    .Y(_05524_));
 OA211x2_ASAP7_75t_R _12409_ (.A1(_03284_),
    .A2(_03288_),
    .B(_04885_),
    .C(_05524_),
    .Y(_05525_));
 AOI21x1_ASAP7_75t_R _12410_ (.A1(_05444_),
    .A2(_05523_),
    .B(_05525_),
    .Y(_05526_));
 AND4x1_ASAP7_75t_R _12411_ (.A(_04786_),
    .B(_04791_),
    .C(_05522_),
    .D(_05526_),
    .Y(_05527_));
 OA22x2_ASAP7_75t_R _12412_ (.A1(_00620_),
    .A2(_04896_),
    .B1(_04472_),
    .B2(_00621_),
    .Y(_05528_));
 AND3x1_ASAP7_75t_R _12413_ (.A(_05440_),
    .B(_03835_),
    .C(_05528_),
    .Y(_05529_));
 OA22x2_ASAP7_75t_R _12414_ (.A1(_00626_),
    .A2(_04560_),
    .B1(_04005_),
    .B2(_00627_),
    .Y(_05530_));
 OA222x2_ASAP7_75t_R _12415_ (.A1(_00630_),
    .A2(_03306_),
    .B1(_03486_),
    .B2(_00631_),
    .C1(_03277_),
    .C2(_03468_),
    .Y(_05531_));
 AO21x1_ASAP7_75t_R _12416_ (.A1(_03394_),
    .A2(_05530_),
    .B(_05531_),
    .Y(_05532_));
 OA22x2_ASAP7_75t_R _12417_ (.A1(_00618_),
    .A2(_03329_),
    .B1(_03765_),
    .B2(_00619_),
    .Y(_05533_));
 OA222x2_ASAP7_75t_R _12418_ (.A1(_00622_),
    .A2(_03428_),
    .B1(_03356_),
    .B2(_00623_),
    .C1(_03277_),
    .C2(_03468_),
    .Y(_05534_));
 AO221x1_ASAP7_75t_R _12419_ (.A1(_05229_),
    .A2(net9),
    .B1(_04447_),
    .B2(_05533_),
    .C(_05534_),
    .Y(_05535_));
 OA211x2_ASAP7_75t_R _12420_ (.A1(_03300_),
    .A2(_05532_),
    .B(_05535_),
    .C(_03444_),
    .Y(_05536_));
 AND2x2_ASAP7_75t_R _12421_ (.A(_00617_),
    .B(_03409_),
    .Y(_05537_));
 AO21x1_ASAP7_75t_R _12422_ (.A1(_00616_),
    .A2(_03451_),
    .B(_05537_),
    .Y(_05538_));
 AND3x1_ASAP7_75t_R _12423_ (.A(_03300_),
    .B(_03484_),
    .C(_05538_),
    .Y(_05539_));
 OR4x1_ASAP7_75t_R _12424_ (.A(_04003_),
    .B(_05529_),
    .C(_05536_),
    .D(_05539_),
    .Y(_05540_));
 OA22x2_ASAP7_75t_R _12425_ (.A1(_00606_),
    .A2(_05227_),
    .B1(_05241_),
    .B2(_00607_),
    .Y(_05541_));
 OR3x1_ASAP7_75t_R _12426_ (.A(_04899_),
    .B(_05444_),
    .C(_05541_),
    .Y(_05542_));
 OA22x2_ASAP7_75t_R _12427_ (.A1(_00610_),
    .A2(_03350_),
    .B1(_03383_),
    .B2(_00611_),
    .Y(_05543_));
 OA222x2_ASAP7_75t_R _12428_ (.A1(_00614_),
    .A2(_05106_),
    .B1(_04445_),
    .B2(_00615_),
    .C1(_03470_),
    .C2(_05314_),
    .Y(_05544_));
 AO21x1_ASAP7_75t_R _12429_ (.A1(_05318_),
    .A2(_05543_),
    .B(_05544_),
    .Y(_05545_));
 OA22x2_ASAP7_75t_R _12430_ (.A1(_00602_),
    .A2(_03350_),
    .B1(_04473_),
    .B2(_00603_),
    .Y(_05546_));
 OR3x2_ASAP7_75t_R _12431_ (.A(_03461_),
    .B(_05127_),
    .C(_05546_),
    .Y(_05547_));
 OA21x2_ASAP7_75t_R _12432_ (.A1(_03300_),
    .A2(_05545_),
    .B(_05547_),
    .Y(_05548_));
 AND3x1_ASAP7_75t_R _12433_ (.A(_03444_),
    .B(_05542_),
    .C(_05548_),
    .Y(_05549_));
 OA22x2_ASAP7_75t_R _12434_ (.A1(_00604_),
    .A2(_05227_),
    .B1(_04472_),
    .B2(_00605_),
    .Y(_05550_));
 AND3x1_ASAP7_75t_R _12435_ (.A(_05440_),
    .B(_03835_),
    .C(_05550_),
    .Y(_05551_));
 OA211x2_ASAP7_75t_R _12436_ (.A1(_03226_),
    .A2(_03311_),
    .B(_04022_),
    .C(_00609_),
    .Y(_05552_));
 AO21x1_ASAP7_75t_R _12437_ (.A1(_00608_),
    .A2(_04445_),
    .B(_05552_),
    .Y(_05553_));
 OA222x2_ASAP7_75t_R _12438_ (.A1(_03470_),
    .A2(_03468_),
    .B1(_03335_),
    .B2(_00613_),
    .C1(_00612_),
    .C2(_04132_),
    .Y(_05554_));
 AO21x1_ASAP7_75t_R _12439_ (.A1(_03394_),
    .A2(_05553_),
    .B(_05554_),
    .Y(_05555_));
 AND3x1_ASAP7_75t_R _12440_ (.A(_04786_),
    .B(_04791_),
    .C(_05555_),
    .Y(_05556_));
 BUFx10_ASAP7_75t_R _12441_ (.A(_04473_),
    .Y(_05557_));
 OA21x2_ASAP7_75t_R _12442_ (.A1(_00601_),
    .A2(_05557_),
    .B(_03421_),
    .Y(_05558_));
 OR4x1_ASAP7_75t_R _12443_ (.A(_05032_),
    .B(_05551_),
    .C(_05556_),
    .D(_05558_),
    .Y(_05559_));
 OAI22x1_ASAP7_75t_R _12444_ (.A1(_05527_),
    .A2(_05540_),
    .B1(_05549_),
    .B2(_05559_),
    .Y(_05560_));
 INVx2_ASAP7_75t_R _12445_ (.A(_05560_),
    .Y(_09647_));
 AOI21x1_ASAP7_75t_R _12446_ (.A1(_04979_),
    .A2(_05470_),
    .B(_04977_),
    .Y(_05561_));
 OR2x2_ASAP7_75t_R _12447_ (.A(_03218_),
    .B(_05092_),
    .Y(_05562_));
 NAND2x1_ASAP7_75t_R _12448_ (.A(_05092_),
    .B(_05468_),
    .Y(_05563_));
 AO21x1_ASAP7_75t_R _12449_ (.A1(_05562_),
    .A2(_05563_),
    .B(_03777_),
    .Y(_05564_));
 AOI21x1_ASAP7_75t_R _12450_ (.A1(_05561_),
    .A2(_05564_),
    .B(_03779_),
    .Y(_09742_));
 AND2x2_ASAP7_75t_R _12451_ (.A(_04267_),
    .B(_00636_),
    .Y(_05565_));
 AO21x1_ASAP7_75t_R _12452_ (.A1(_03062_),
    .A2(_00635_),
    .B(_05565_),
    .Y(_05566_));
 AO21x1_ASAP7_75t_R _12453_ (.A1(_04722_),
    .A2(_05566_),
    .B(_04416_),
    .Y(_05567_));
 AO22x1_ASAP7_75t_R _12454_ (.A1(_03910_),
    .A2(_00633_),
    .B1(_00634_),
    .B2(_03591_),
    .Y(_05568_));
 AO22x1_ASAP7_75t_R _12455_ (.A1(_04493_),
    .A2(_00633_),
    .B1(_05568_),
    .B2(_03028_),
    .Y(_05569_));
 AO21x1_ASAP7_75t_R _12456_ (.A1(_03201_),
    .A2(_05567_),
    .B(_05569_),
    .Y(_05570_));
 AND2x2_ASAP7_75t_R _12457_ (.A(_03894_),
    .B(_00640_),
    .Y(_05571_));
 AO21x1_ASAP7_75t_R _12458_ (.A1(_03685_),
    .A2(_00639_),
    .B(_05571_),
    .Y(_05572_));
 AND3x1_ASAP7_75t_R _12459_ (.A(_03898_),
    .B(_03473_),
    .C(_00638_),
    .Y(_05573_));
 AO21x1_ASAP7_75t_R _12460_ (.A1(_00637_),
    .A2(_03897_),
    .B(_05573_),
    .Y(_05574_));
 AO221x1_ASAP7_75t_R _12461_ (.A1(_03893_),
    .A2(_05572_),
    .B1(_05574_),
    .B2(_03901_),
    .C(_03902_),
    .Y(_05575_));
 AND3x4_ASAP7_75t_R _12462_ (.A(_04404_),
    .B(_05570_),
    .C(_05575_),
    .Y(_05576_));
 AND2x2_ASAP7_75t_R _12463_ (.A(_03894_),
    .B(_00648_),
    .Y(_05577_));
 AO21x1_ASAP7_75t_R _12464_ (.A1(_03685_),
    .A2(_00647_),
    .B(_05577_),
    .Y(_05578_));
 AND3x1_ASAP7_75t_R _12465_ (.A(_03898_),
    .B(_03473_),
    .C(_00646_),
    .Y(_05579_));
 AO21x1_ASAP7_75t_R _12466_ (.A1(_00645_),
    .A2(_03897_),
    .B(_05579_),
    .Y(_05580_));
 AO221x1_ASAP7_75t_R _12467_ (.A1(_03893_),
    .A2(_05578_),
    .B1(_05580_),
    .B2(_03901_),
    .C(_03902_),
    .Y(_05581_));
 AO22x1_ASAP7_75t_R _12468_ (.A1(_03905_),
    .A2(_00641_),
    .B1(_00642_),
    .B2(_03906_),
    .Y(_05582_));
 AND2x2_ASAP7_75t_R _12469_ (.A(_04267_),
    .B(_00644_),
    .Y(_05583_));
 AO21x1_ASAP7_75t_R _12470_ (.A1(_03062_),
    .A2(_00643_),
    .B(_05583_),
    .Y(_05584_));
 AO21x1_ASAP7_75t_R _12471_ (.A1(_04722_),
    .A2(_05584_),
    .B(_04416_),
    .Y(_05585_));
 AO21x1_ASAP7_75t_R _12472_ (.A1(_03904_),
    .A2(_05582_),
    .B(_05585_),
    .Y(_05586_));
 AND3x4_ASAP7_75t_R _12473_ (.A(_04098_),
    .B(_05581_),
    .C(_05586_),
    .Y(_05587_));
 OR3x1_ASAP7_75t_R _12474_ (.A(_04043_),
    .B(_05576_),
    .C(_05587_),
    .Y(_05588_));
 AND2x2_ASAP7_75t_R _12475_ (.A(_03898_),
    .B(_00664_),
    .Y(_05589_));
 AO21x1_ASAP7_75t_R _12476_ (.A1(_03112_),
    .A2(_00663_),
    .B(_05589_),
    .Y(_05590_));
 AND3x1_ASAP7_75t_R _12477_ (.A(_03048_),
    .B(_03034_),
    .C(_00662_),
    .Y(_05591_));
 AO21x1_ASAP7_75t_R _12478_ (.A1(_00661_),
    .A2(_04393_),
    .B(_05591_),
    .Y(_05592_));
 AO221x1_ASAP7_75t_R _12479_ (.A1(_04497_),
    .A2(_05590_),
    .B1(_05592_),
    .B2(_03922_),
    .C(_04397_),
    .Y(_05593_));
 AND2x2_ASAP7_75t_R _12480_ (.A(_03073_),
    .B(_00659_),
    .Y(_05594_));
 AO21x1_ASAP7_75t_R _12481_ (.A1(_03589_),
    .A2(_00657_),
    .B(_05594_),
    .Y(_05595_));
 AO21x1_ASAP7_75t_R _12482_ (.A1(_00658_),
    .A2(_03561_),
    .B(_04529_),
    .Y(_05596_));
 AO221x1_ASAP7_75t_R _12483_ (.A1(_00660_),
    .A2(_04077_),
    .B1(_05595_),
    .B2(_03139_),
    .C(_05596_),
    .Y(_05597_));
 AND3x1_ASAP7_75t_R _12484_ (.A(_03174_),
    .B(_05593_),
    .C(_05597_),
    .Y(_05598_));
 AND2x2_ASAP7_75t_R _12485_ (.A(_04499_),
    .B(_00656_),
    .Y(_05599_));
 AO21x1_ASAP7_75t_R _12486_ (.A1(_04498_),
    .A2(_00655_),
    .B(_05599_),
    .Y(_05600_));
 AND3x1_ASAP7_75t_R _12487_ (.A(_04502_),
    .B(_04503_),
    .C(_00654_),
    .Y(_05601_));
 AO21x1_ASAP7_75t_R _12488_ (.A1(_00653_),
    .A2(_03897_),
    .B(_05601_),
    .Y(_05602_));
 AO221x1_ASAP7_75t_R _12489_ (.A1(_04497_),
    .A2(_05600_),
    .B1(_05602_),
    .B2(_03922_),
    .C(_03902_),
    .Y(_05603_));
 AND2x2_ASAP7_75t_R _12490_ (.A(_03073_),
    .B(_00651_),
    .Y(_05604_));
 AO21x1_ASAP7_75t_R _12491_ (.A1(_03665_),
    .A2(_00649_),
    .B(_05604_),
    .Y(_05605_));
 AO21x1_ASAP7_75t_R _12492_ (.A1(_00650_),
    .A2(_03561_),
    .B(_04529_),
    .Y(_05606_));
 AO221x2_ASAP7_75t_R _12493_ (.A1(_00652_),
    .A2(_04077_),
    .B1(_05605_),
    .B2(_04528_),
    .C(_05606_),
    .Y(_05607_));
 AND3x1_ASAP7_75t_R _12494_ (.A(_04404_),
    .B(_05603_),
    .C(_05607_),
    .Y(_05608_));
 OR3x4_ASAP7_75t_R _12495_ (.A(_04100_),
    .B(_05598_),
    .C(_05608_),
    .Y(_05609_));
 AOI21x1_ASAP7_75t_R _12496_ (.A1(_05588_),
    .A2(_05609_),
    .B(_03781_),
    .Y(_05610_));
 AND2x2_ASAP7_75t_R _12497_ (.A(_04422_),
    .B(_05610_),
    .Y(_05611_));
 AOI21x1_ASAP7_75t_R _12498_ (.A1(_03645_),
    .A2(_09742_),
    .B(_05611_),
    .Y(_05612_));
 XNOR2x1_ASAP7_75t_R _12499_ (.B(_05612_),
    .Y(_09651_),
    .A(_04610_));
 INVx1_ASAP7_75t_R _12500_ (.A(_09651_),
    .Y(_09653_));
 INVx1_ASAP7_75t_R _12501_ (.A(_00662_),
    .Y(_05613_));
 INVx1_ASAP7_75t_R _12502_ (.A(_00661_),
    .Y(_05614_));
 AO32x1_ASAP7_75t_R _12503_ (.A1(_03200_),
    .A2(_05335_),
    .A3(_05613_),
    .B1(_03450_),
    .B2(_05614_),
    .Y(_05615_));
 INVx2_ASAP7_75t_R _12504_ (.A(_00658_),
    .Y(_05616_));
 NAND2x1_ASAP7_75t_R _12505_ (.A(_00657_),
    .B(_03765_),
    .Y(_05617_));
 OA211x2_ASAP7_75t_R _12506_ (.A1(_05616_),
    .A2(_04005_),
    .B(_05617_),
    .C(_03393_),
    .Y(_05618_));
 AOI211x1_ASAP7_75t_R _12507_ (.A1(_05440_),
    .A2(_05615_),
    .B(_05618_),
    .C(_03341_),
    .Y(_05619_));
 AND3x1_ASAP7_75t_R _12508_ (.A(_00659_),
    .B(_03208_),
    .C(_03321_),
    .Y(_05620_));
 AO21x1_ASAP7_75t_R _12509_ (.A1(_00663_),
    .A2(_03747_),
    .B(_05620_),
    .Y(_05621_));
 OA22x2_ASAP7_75t_R _12510_ (.A1(_00664_),
    .A2(_03732_),
    .B1(_03733_),
    .B2(_00660_),
    .Y(_05622_));
 OA211x2_ASAP7_75t_R _12511_ (.A1(_03330_),
    .A2(_05621_),
    .B(_05622_),
    .C(_04432_),
    .Y(_05623_));
 OA21x2_ASAP7_75t_R _12512_ (.A1(_05619_),
    .A2(_05623_),
    .B(_04899_),
    .Y(_05624_));
 INVx1_ASAP7_75t_R _12513_ (.A(_00651_),
    .Y(_05625_));
 INVx1_ASAP7_75t_R _12514_ (.A(_00652_),
    .Y(_05626_));
 AOI22x1_ASAP7_75t_R _12515_ (.A1(_05625_),
    .A2(_03466_),
    .B1(_03408_),
    .B2(_05626_),
    .Y(_05627_));
 AND2x2_ASAP7_75t_R _12516_ (.A(_00655_),
    .B(_03435_),
    .Y(_05628_));
 AO221x2_ASAP7_75t_R _12517_ (.A1(_03250_),
    .A2(_03387_),
    .B1(_03384_),
    .B2(_00656_),
    .C(_05628_),
    .Y(_05629_));
 OA21x2_ASAP7_75t_R _12518_ (.A1(_03504_),
    .A2(_05627_),
    .B(_05629_),
    .Y(_05630_));
 INVx1_ASAP7_75t_R _12519_ (.A(_00653_),
    .Y(_05631_));
 INVx1_ASAP7_75t_R _12520_ (.A(_00654_),
    .Y(_05632_));
 AOI22x1_ASAP7_75t_R _12521_ (.A1(_05631_),
    .A2(_03437_),
    .B1(_04466_),
    .B2(_05632_),
    .Y(_05633_));
 AND2x2_ASAP7_75t_R _12522_ (.A(_00650_),
    .B(_03408_),
    .Y(_05634_));
 AO21x1_ASAP7_75t_R _12523_ (.A1(_00649_),
    .A2(_03486_),
    .B(_05634_),
    .Y(_05635_));
 OA222x2_ASAP7_75t_R _12524_ (.A1(_03855_),
    .A2(_05630_),
    .B1(_05633_),
    .B2(_03979_),
    .C1(_03845_),
    .C2(_05635_),
    .Y(_05636_));
 AO21x1_ASAP7_75t_R _12525_ (.A1(_03300_),
    .A2(_05636_),
    .B(_03862_),
    .Y(_05637_));
 OA222x2_ASAP7_75t_R _12526_ (.A1(_03097_),
    .A2(_03965_),
    .B1(_00640_),
    .B2(_03732_),
    .C1(_03733_),
    .C2(_00636_),
    .Y(_05638_));
 AND3x1_ASAP7_75t_R _12527_ (.A(_00635_),
    .B(_03208_),
    .C(_03736_),
    .Y(_05639_));
 AO221x1_ASAP7_75t_R _12528_ (.A1(_03064_),
    .A2(_05124_),
    .B1(_00639_),
    .B2(_03504_),
    .C(_05639_),
    .Y(_05640_));
 AO21x2_ASAP7_75t_R _12529_ (.A1(_05638_),
    .A2(_05640_),
    .B(_03836_),
    .Y(_05641_));
 INVx2_ASAP7_75t_R _12530_ (.A(_00637_),
    .Y(_05642_));
 INVx2_ASAP7_75t_R _12531_ (.A(_00638_),
    .Y(_05643_));
 AO22x1_ASAP7_75t_R _12532_ (.A1(_05642_),
    .A2(_03437_),
    .B1(_04466_),
    .B2(_05643_),
    .Y(_05644_));
 NAND2x1_ASAP7_75t_R _12533_ (.A(_03540_),
    .B(_05644_),
    .Y(_05645_));
 AND2x2_ASAP7_75t_R _12534_ (.A(_00633_),
    .B(_03765_),
    .Y(_05646_));
 AO221x1_ASAP7_75t_R _12535_ (.A1(_00634_),
    .A2(_03409_),
    .B1(_03411_),
    .B2(_03245_),
    .C(_05646_),
    .Y(_05647_));
 AND3x1_ASAP7_75t_R _12536_ (.A(_04009_),
    .B(_04586_),
    .C(_00648_),
    .Y(_05648_));
 AO21x1_ASAP7_75t_R _12537_ (.A1(_00647_),
    .A2(_03335_),
    .B(_05648_),
    .Y(_05649_));
 OR3x1_ASAP7_75t_R _12538_ (.A(_03855_),
    .B(_04447_),
    .C(_05649_),
    .Y(_05650_));
 OA211x2_ASAP7_75t_R _12539_ (.A1(_03487_),
    .A2(_03310_),
    .B(_03312_),
    .C(_00642_),
    .Y(_05651_));
 AO21x1_ASAP7_75t_R _12540_ (.A1(_00641_),
    .A2(_03431_),
    .B(_05651_),
    .Y(_05652_));
 OA222x2_ASAP7_75t_R _12541_ (.A1(_00643_),
    .A2(_03522_),
    .B1(_03413_),
    .B2(_00644_),
    .C1(_03277_),
    .C2(_03381_),
    .Y(_05653_));
 AO21x1_ASAP7_75t_R _12542_ (.A1(_03855_),
    .A2(_05652_),
    .B(_05653_),
    .Y(_05654_));
 INVx1_ASAP7_75t_R _12543_ (.A(_00646_),
    .Y(_05655_));
 INVx1_ASAP7_75t_R _12544_ (.A(_00645_),
    .Y(_05656_));
 AO32x1_ASAP7_75t_R _12545_ (.A1(_04692_),
    .A2(_04586_),
    .A3(_05655_),
    .B1(_03449_),
    .B2(_05656_),
    .Y(_05657_));
 NAND2x1_ASAP7_75t_R _12546_ (.A(_03361_),
    .B(_05657_),
    .Y(_05658_));
 OA211x2_ASAP7_75t_R _12547_ (.A1(_03441_),
    .A2(_05654_),
    .B(_05658_),
    .C(_03888_),
    .Y(_05659_));
 AO32x1_ASAP7_75t_R _12548_ (.A1(_05641_),
    .A2(_05645_),
    .A3(_05647_),
    .B1(_05650_),
    .B2(_05659_),
    .Y(_05660_));
 OA22x2_ASAP7_75t_R _12549_ (.A1(_05624_),
    .A2(_05637_),
    .B1(_05660_),
    .B2(_03426_),
    .Y(_05661_));
 BUFx6f_ASAP7_75t_R _12550_ (.A(_05661_),
    .Y(_09652_));
 OA21x2_ASAP7_75t_R _12551_ (.A1(_03218_),
    .A2(_03715_),
    .B(_05561_),
    .Y(_05662_));
 OA21x2_ASAP7_75t_R _12552_ (.A1(_03218_),
    .A2(_03265_),
    .B(_03710_),
    .Y(_05663_));
 OAI22x1_ASAP7_75t_R _12553_ (.A1(_04987_),
    .A2(_05662_),
    .B1(_05663_),
    .B2(_05092_),
    .Y(_09740_));
 AO22x1_ASAP7_75t_R _12554_ (.A1(_03932_),
    .A2(_00690_),
    .B1(_00691_),
    .B2(_03591_),
    .Y(_05664_));
 AND2x2_ASAP7_75t_R _12555_ (.A(_03090_),
    .B(_00693_),
    .Y(_05665_));
 AO21x1_ASAP7_75t_R _12556_ (.A1(_03572_),
    .A2(_00692_),
    .B(_05665_),
    .Y(_05666_));
 AO221x1_ASAP7_75t_R _12557_ (.A1(_03104_),
    .A2(_00690_),
    .B1(_03909_),
    .B2(_05666_),
    .C(_03936_),
    .Y(_05667_));
 AO21x1_ASAP7_75t_R _12558_ (.A1(_03132_),
    .A2(_05664_),
    .B(_05667_),
    .Y(_05668_));
 AND2x2_ASAP7_75t_R _12559_ (.A(_03675_),
    .B(_00697_),
    .Y(_05669_));
 AO21x1_ASAP7_75t_R _12560_ (.A1(_03625_),
    .A2(_00696_),
    .B(_05669_),
    .Y(_05670_));
 AND3x1_ASAP7_75t_R _12561_ (.A(_03678_),
    .B(_03117_),
    .C(_00695_),
    .Y(_05671_));
 AO21x1_ASAP7_75t_R _12562_ (.A1(_00694_),
    .A2(_03289_),
    .B(_05671_),
    .Y(_05672_));
 AO221x1_ASAP7_75t_R _12563_ (.A1(_03674_),
    .A2(_05670_),
    .B1(_05672_),
    .B2(_03681_),
    .C(_03636_),
    .Y(_05673_));
 AND3x1_ASAP7_75t_R _12564_ (.A(_03142_),
    .B(_05668_),
    .C(_05673_),
    .Y(_05674_));
 INVx3_ASAP7_75t_R _12565_ (.A(_05674_),
    .Y(_05675_));
 AO22x1_ASAP7_75t_R _12566_ (.A1(_03932_),
    .A2(_00674_),
    .B1(_00675_),
    .B2(_03591_),
    .Y(_05676_));
 AND2x2_ASAP7_75t_R _12567_ (.A(_03090_),
    .B(_00677_),
    .Y(_05677_));
 AO21x1_ASAP7_75t_R _12568_ (.A1(_03572_),
    .A2(_00676_),
    .B(_05677_),
    .Y(_05678_));
 AO221x1_ASAP7_75t_R _12569_ (.A1(_03104_),
    .A2(_00674_),
    .B1(_03908_),
    .B2(_05678_),
    .C(_03913_),
    .Y(_05679_));
 AO21x1_ASAP7_75t_R _12570_ (.A1(_03132_),
    .A2(_05676_),
    .B(_05679_),
    .Y(_05680_));
 AND2x2_ASAP7_75t_R _12571_ (.A(_03675_),
    .B(_00681_),
    .Y(_05681_));
 AO21x1_ASAP7_75t_R _12572_ (.A1(_03111_),
    .A2(_00680_),
    .B(_05681_),
    .Y(_05682_));
 AND3x1_ASAP7_75t_R _12573_ (.A(_03678_),
    .B(_03117_),
    .C(_00679_),
    .Y(_05683_));
 AO21x1_ASAP7_75t_R _12574_ (.A1(_00678_),
    .A2(_03123_),
    .B(_05683_),
    .Y(_05684_));
 AO221x1_ASAP7_75t_R _12575_ (.A1(_03087_),
    .A2(_05682_),
    .B1(_05684_),
    .B2(_03635_),
    .C(_03636_),
    .Y(_05685_));
 AND3x1_ASAP7_75t_R _12576_ (.A(_03154_),
    .B(_05680_),
    .C(_05685_),
    .Y(_05686_));
 INVx1_ASAP7_75t_R _12577_ (.A(_05686_),
    .Y(_05687_));
 INVx2_ASAP7_75t_R _12578_ (.A(_00688_),
    .Y(_05688_));
 NAND2x1_ASAP7_75t_R _12579_ (.A(_04267_),
    .B(_00689_),
    .Y(_05689_));
 OA21x2_ASAP7_75t_R _12580_ (.A1(_03155_),
    .A2(_05688_),
    .B(_05689_),
    .Y(_05690_));
 OA21x2_ASAP7_75t_R _12581_ (.A1(_03665_),
    .A2(_05690_),
    .B(_03936_),
    .Y(_05691_));
 INVx1_ASAP7_75t_R _12582_ (.A(_00687_),
    .Y(_05692_));
 OR3x1_ASAP7_75t_R _12583_ (.A(_03111_),
    .B(_04492_),
    .C(_05692_),
    .Y(_05693_));
 INVx3_ASAP7_75t_R _12584_ (.A(_00686_),
    .Y(_05694_));
 AO21x1_ASAP7_75t_R _12585_ (.A1(_03048_),
    .A2(_03034_),
    .B(_05694_),
    .Y(_05695_));
 AO21x1_ASAP7_75t_R _12586_ (.A1(_05693_),
    .A2(_05695_),
    .B(_03925_),
    .Y(_05696_));
 AO22x1_ASAP7_75t_R _12587_ (.A1(_03932_),
    .A2(_00682_),
    .B1(_00683_),
    .B2(_03591_),
    .Y(_05697_));
 AND2x2_ASAP7_75t_R _12588_ (.A(_03090_),
    .B(_00685_),
    .Y(_05698_));
 AO21x1_ASAP7_75t_R _12589_ (.A1(_03572_),
    .A2(_00684_),
    .B(_05698_),
    .Y(_05699_));
 AO221x1_ASAP7_75t_R _12590_ (.A1(_03104_),
    .A2(_00682_),
    .B1(_03908_),
    .B2(_05699_),
    .C(_03936_),
    .Y(_05700_));
 AOI21x1_ASAP7_75t_R _12591_ (.A1(_03132_),
    .A2(_05697_),
    .B(_05700_),
    .Y(_05701_));
 AO21x1_ASAP7_75t_R _12592_ (.A1(_05691_),
    .A2(_05696_),
    .B(_05701_),
    .Y(_05702_));
 AND2x2_ASAP7_75t_R _12593_ (.A(_03675_),
    .B(_00673_),
    .Y(_05703_));
 AO21x1_ASAP7_75t_R _12594_ (.A1(_03625_),
    .A2(_00672_),
    .B(_05703_),
    .Y(_05704_));
 AND3x1_ASAP7_75t_R _12595_ (.A(_03678_),
    .B(_03117_),
    .C(_00671_),
    .Y(_05705_));
 AO21x1_ASAP7_75t_R _12596_ (.A1(_00670_),
    .A2(_03289_),
    .B(_05705_),
    .Y(_05706_));
 AO221x1_ASAP7_75t_R _12597_ (.A1(_03674_),
    .A2(_05704_),
    .B1(_05706_),
    .B2(_03681_),
    .C(_03695_),
    .Y(_05707_));
 AO22x1_ASAP7_75t_R _12598_ (.A1(_03573_),
    .A2(_00666_),
    .B1(_00667_),
    .B2(_03946_),
    .Y(_05708_));
 AND2x2_ASAP7_75t_R _12599_ (.A(_03090_),
    .B(_00669_),
    .Y(_05709_));
 AO21x1_ASAP7_75t_R _12600_ (.A1(_03572_),
    .A2(_00668_),
    .B(_05709_),
    .Y(_05710_));
 AO221x1_ASAP7_75t_R _12601_ (.A1(_03104_),
    .A2(_00666_),
    .B1(_03909_),
    .B2(_05710_),
    .C(_03936_),
    .Y(_05711_));
 AO21x1_ASAP7_75t_R _12602_ (.A1(_03132_),
    .A2(_05708_),
    .B(_05711_),
    .Y(_05712_));
 AOI21x1_ASAP7_75t_R _12603_ (.A1(_05707_),
    .A2(_05712_),
    .B(_03142_),
    .Y(_05713_));
 AO21x1_ASAP7_75t_R _12604_ (.A1(_03142_),
    .A2(_05702_),
    .B(_05713_),
    .Y(_05714_));
 AO32x2_ASAP7_75t_R _12605_ (.A1(_03174_),
    .A2(_05675_),
    .A3(_05687_),
    .B1(_03128_),
    .B2(_05714_),
    .Y(_05715_));
 OR2x2_ASAP7_75t_R _12606_ (.A(_03270_),
    .B(_05715_),
    .Y(_05716_));
 OA21x2_ASAP7_75t_R _12607_ (.A1(_04159_),
    .A2(_09740_),
    .B(_05716_),
    .Y(_05717_));
 XNOR2x1_ASAP7_75t_R _12608_ (.B(_05717_),
    .Y(_09656_),
    .A(_03259_));
 INVx1_ASAP7_75t_R _12609_ (.A(_09656_),
    .Y(_09658_));
 OA222x2_ASAP7_75t_R _12610_ (.A1(_04493_),
    .A2(_03965_),
    .B1(_00673_),
    .B2(_03732_),
    .C1(_03733_),
    .C2(_00669_),
    .Y(_05718_));
 AND3x1_ASAP7_75t_R _12611_ (.A(_00668_),
    .B(_03261_),
    .C(_04575_),
    .Y(_05719_));
 AO221x1_ASAP7_75t_R _12612_ (.A1(_03021_),
    .A2(_05335_),
    .B1(_00672_),
    .B2(_03747_),
    .C(_05719_),
    .Y(_05720_));
 AO21x2_ASAP7_75t_R _12613_ (.A1(_05718_),
    .A2(_05720_),
    .B(_04458_),
    .Y(_05721_));
 INVx1_ASAP7_75t_R _12614_ (.A(_00670_),
    .Y(_05722_));
 INVx1_ASAP7_75t_R _12615_ (.A(_00671_),
    .Y(_05723_));
 AO22x2_ASAP7_75t_R _12616_ (.A1(_05722_),
    .A2(_03397_),
    .B1(_03401_),
    .B2(_05723_),
    .Y(_05724_));
 INVx3_ASAP7_75t_R _12617_ (.A(_00666_),
    .Y(_01225_));
 INVx1_ASAP7_75t_R _12618_ (.A(_00667_),
    .Y(_05725_));
 AND2x2_ASAP7_75t_R _12619_ (.A(_05725_),
    .B(_03454_),
    .Y(_05726_));
 AO21x1_ASAP7_75t_R _12620_ (.A1(_01225_),
    .A2(_04451_),
    .B(_05726_),
    .Y(_05727_));
 AOI22x1_ASAP7_75t_R _12621_ (.A1(_04891_),
    .A2(_05724_),
    .B1(_05727_),
    .B2(_03448_),
    .Y(_05728_));
 AND2x2_ASAP7_75t_R _12622_ (.A(_00674_),
    .B(_03529_),
    .Y(_05729_));
 AO221x2_ASAP7_75t_R _12623_ (.A1(_00675_),
    .A2(_03455_),
    .B1(_03411_),
    .B2(_03246_),
    .C(_05729_),
    .Y(_05730_));
 INVx1_ASAP7_75t_R _12624_ (.A(_00679_),
    .Y(_05731_));
 INVx1_ASAP7_75t_R _12625_ (.A(_00678_),
    .Y(_05732_));
 AO32x1_ASAP7_75t_R _12626_ (.A1(_03064_),
    .A2(_05124_),
    .A3(_05731_),
    .B1(_03418_),
    .B2(_05732_),
    .Y(_05733_));
 NAND2x1_ASAP7_75t_R _12627_ (.A(_03457_),
    .B(_05733_),
    .Y(_05734_));
 AND3x1_ASAP7_75t_R _12628_ (.A(_03019_),
    .B(_03970_),
    .C(_00681_),
    .Y(_05735_));
 AO21x1_ASAP7_75t_R _12629_ (.A1(_00680_),
    .A2(_03436_),
    .B(_05735_),
    .Y(_05736_));
 INVx1_ASAP7_75t_R _12630_ (.A(_00677_),
    .Y(_05737_));
 NAND2x1_ASAP7_75t_R _12631_ (.A(_05737_),
    .B(_03400_),
    .Y(_05738_));
 OA21x2_ASAP7_75t_R _12632_ (.A1(_00676_),
    .A2(_03313_),
    .B(_03321_),
    .Y(_05739_));
 AO221x1_ASAP7_75t_R _12633_ (.A1(_03504_),
    .A2(_05736_),
    .B1(_05738_),
    .B2(_05739_),
    .C(_03988_),
    .Y(_05740_));
 OR2x2_ASAP7_75t_R _12634_ (.A(_03371_),
    .B(_05736_),
    .Y(_05741_));
 AND4x2_ASAP7_75t_R _12635_ (.A(_03888_),
    .B(_05734_),
    .C(_05740_),
    .D(_05741_),
    .Y(_05742_));
 AO221x2_ASAP7_75t_R _12636_ (.A1(_05721_),
    .A2(_05728_),
    .B1(_05730_),
    .B2(_05742_),
    .C(_03426_),
    .Y(_05743_));
 INVx1_ASAP7_75t_R _12637_ (.A(_00682_),
    .Y(_05744_));
 INVx1_ASAP7_75t_R _12638_ (.A(_00683_),
    .Y(_05745_));
 AND2x2_ASAP7_75t_R _12639_ (.A(_05745_),
    .B(_03511_),
    .Y(_05746_));
 AO21x1_ASAP7_75t_R _12640_ (.A1(_05744_),
    .A2(_04676_),
    .B(_05746_),
    .Y(_05747_));
 AO22x1_ASAP7_75t_R _12641_ (.A1(_05694_),
    .A2(_03397_),
    .B1(_03541_),
    .B2(_05692_),
    .Y(_05748_));
 INVx1_ASAP7_75t_R _12642_ (.A(_00684_),
    .Y(_05749_));
 INVx1_ASAP7_75t_R _12643_ (.A(_00685_),
    .Y(_05750_));
 AO22x1_ASAP7_75t_R _12644_ (.A1(_05749_),
    .A2(_03847_),
    .B1(_03400_),
    .B2(_05750_),
    .Y(_05751_));
 AND2x2_ASAP7_75t_R _12645_ (.A(_00688_),
    .B(_03436_),
    .Y(_05752_));
 AOI221x1_ASAP7_75t_R _12646_ (.A1(_03251_),
    .A2(_04441_),
    .B1(_03735_),
    .B2(_00689_),
    .C(_05752_),
    .Y(_05753_));
 AO221x1_ASAP7_75t_R _12647_ (.A1(_03021_),
    .A2(net9),
    .B1(_04447_),
    .B2(_05751_),
    .C(_05753_),
    .Y(_05754_));
 AO222x2_ASAP7_75t_R _12648_ (.A1(_03448_),
    .A2(_05747_),
    .B1(_05748_),
    .B2(_04891_),
    .C1(_04349_),
    .C2(_05754_),
    .Y(_05755_));
 INVx2_ASAP7_75t_R _12649_ (.A(_00691_),
    .Y(_05756_));
 NAND2x1_ASAP7_75t_R _12650_ (.A(_00690_),
    .B(_03414_),
    .Y(_05757_));
 OA211x2_ASAP7_75t_R _12651_ (.A1(_05756_),
    .A2(_03432_),
    .B(_03484_),
    .C(_05757_),
    .Y(_05758_));
 INVx2_ASAP7_75t_R _12652_ (.A(_00693_),
    .Y(_05759_));
 OA211x2_ASAP7_75t_R _12653_ (.A1(_03364_),
    .A2(_03365_),
    .B(_03348_),
    .C(_05759_),
    .Y(_05760_));
 INVx2_ASAP7_75t_R _12654_ (.A(_00692_),
    .Y(_05761_));
 AO21x1_ASAP7_75t_R _12655_ (.A1(_05761_),
    .A2(_03334_),
    .B(_03359_),
    .Y(_05762_));
 OA21x2_ASAP7_75t_R _12656_ (.A1(_05760_),
    .A2(_05762_),
    .B(_03381_),
    .Y(_05763_));
 INVx1_ASAP7_75t_R _12657_ (.A(_00696_),
    .Y(_05764_));
 INVx1_ASAP7_75t_R _12658_ (.A(_00697_),
    .Y(_05765_));
 OR3x1_ASAP7_75t_R _12659_ (.A(_03096_),
    .B(_03749_),
    .C(_05765_),
    .Y(_05766_));
 OA21x2_ASAP7_75t_R _12660_ (.A1(_05764_),
    .A2(_03349_),
    .B(_05766_),
    .Y(_05767_));
 OA22x2_ASAP7_75t_R _12661_ (.A1(_03470_),
    .A2(_05763_),
    .B1(_05767_),
    .B2(_04447_),
    .Y(_05768_));
 INVx2_ASAP7_75t_R _12662_ (.A(_00695_),
    .Y(_05769_));
 INVx2_ASAP7_75t_R _12663_ (.A(_00694_),
    .Y(_05770_));
 AO32x1_ASAP7_75t_R _12664_ (.A1(_03473_),
    .A2(_03475_),
    .A3(_05769_),
    .B1(_03431_),
    .B2(_05770_),
    .Y(_05771_));
 OA211x2_ASAP7_75t_R _12665_ (.A1(_03273_),
    .A2(_03287_),
    .B(_03361_),
    .C(_05771_),
    .Y(_05772_));
 OR4x2_ASAP7_75t_R _12666_ (.A(_04552_),
    .B(_05758_),
    .C(_05768_),
    .D(_05772_),
    .Y(_05773_));
 NAND3x2_ASAP7_75t_R _12667_ (.B(_05755_),
    .C(_05773_),
    .Y(_05774_),
    .A(_05032_));
 NAND2x2_ASAP7_75t_R _12668_ (.A(_05743_),
    .B(_05774_),
    .Y(_09655_));
 INVx1_ASAP7_75t_R _12669_ (.A(_09655_),
    .Y(_09657_));
 NOR2x2_ASAP7_75t_R _12670_ (.A(_03249_),
    .B(_03254_),
    .Y(_05775_));
 BUFx3_ASAP7_75t_R _12671_ (.A(_05775_),
    .Y(_05776_));
 BUFx4f_ASAP7_75t_R _12672_ (.A(_05776_),
    .Y(_05777_));
 AND3x1_ASAP7_75t_R _12673_ (.A(_04981_),
    .B(_04977_),
    .C(_05092_),
    .Y(_05778_));
 AO221x2_ASAP7_75t_R _12674_ (.A1(_05370_),
    .A2(_04979_),
    .B1(_03279_),
    .B2(_05777_),
    .C(_05778_),
    .Y(_09738_));
 AND2x2_ASAP7_75t_R _12675_ (.A(_04408_),
    .B(_00702_),
    .Y(_05779_));
 AO21x1_ASAP7_75t_R _12676_ (.A1(_04851_),
    .A2(_00701_),
    .B(_05779_),
    .Y(_05780_));
 AO21x1_ASAP7_75t_R _12677_ (.A1(_04850_),
    .A2(_05780_),
    .B(_03078_),
    .Y(_05781_));
 AO22x1_ASAP7_75t_R _12678_ (.A1(_03905_),
    .A2(_00699_),
    .B1(_00700_),
    .B2(_03906_),
    .Y(_05782_));
 AO22x1_ASAP7_75t_R _12679_ (.A1(_03131_),
    .A2(_00699_),
    .B1(_05782_),
    .B2(_04381_),
    .Y(_05783_));
 AO21x1_ASAP7_75t_R _12680_ (.A1(_03216_),
    .A2(_05781_),
    .B(_05783_),
    .Y(_05784_));
 AND2x2_ASAP7_75t_R _12681_ (.A(_05272_),
    .B(_00706_),
    .Y(_05785_));
 AO21x1_ASAP7_75t_R _12682_ (.A1(_03082_),
    .A2(_00705_),
    .B(_05785_),
    .Y(_05786_));
 BUFx6f_ASAP7_75t_R _12683_ (.A(_03577_),
    .Y(_05787_));
 AND3x1_ASAP7_75t_R _12684_ (.A(_05266_),
    .B(_03200_),
    .C(_00704_),
    .Y(_05788_));
 AO21x1_ASAP7_75t_R _12685_ (.A1(_00703_),
    .A2(_05787_),
    .B(_05788_),
    .Y(_05789_));
 BUFx6f_ASAP7_75t_R _12686_ (.A(_03582_),
    .Y(_05790_));
 AO221x1_ASAP7_75t_R _12687_ (.A1(_05410_),
    .A2(_05786_),
    .B1(_05789_),
    .B2(_05790_),
    .C(_05077_),
    .Y(_05791_));
 AND3x1_ASAP7_75t_R _12688_ (.A(_05034_),
    .B(_05784_),
    .C(_05791_),
    .Y(_05792_));
 BUFx6f_ASAP7_75t_R _12689_ (.A(_03119_),
    .Y(_05793_));
 AND2x2_ASAP7_75t_R _12690_ (.A(_05044_),
    .B(_00714_),
    .Y(_05794_));
 AO21x1_ASAP7_75t_R _12691_ (.A1(_04095_),
    .A2(_00713_),
    .B(_05794_),
    .Y(_05795_));
 AND3x1_ASAP7_75t_R _12692_ (.A(_05266_),
    .B(_03145_),
    .C(_00712_),
    .Y(_05796_));
 AO21x1_ASAP7_75t_R _12693_ (.A1(_00711_),
    .A2(_05787_),
    .B(_05796_),
    .Y(_05797_));
 BUFx6f_ASAP7_75t_R _12694_ (.A(_03583_),
    .Y(_05798_));
 AO221x1_ASAP7_75t_R _12695_ (.A1(_05410_),
    .A2(_05795_),
    .B1(_05797_),
    .B2(_05790_),
    .C(_05798_),
    .Y(_05799_));
 AO22x1_ASAP7_75t_R _12696_ (.A1(_03139_),
    .A2(_00707_),
    .B1(_00708_),
    .B2(_05370_),
    .Y(_05800_));
 AND2x2_ASAP7_75t_R _12697_ (.A(_04408_),
    .B(_00710_),
    .Y(_05801_));
 AO21x1_ASAP7_75t_R _12698_ (.A1(_04851_),
    .A2(_00709_),
    .B(_05801_),
    .Y(_05802_));
 AO21x1_ASAP7_75t_R _12699_ (.A1(_04850_),
    .A2(_05802_),
    .B(_03078_),
    .Y(_05803_));
 AO21x1_ASAP7_75t_R _12700_ (.A1(_03137_),
    .A2(_05800_),
    .B(_05803_),
    .Y(_05804_));
 AND3x1_ASAP7_75t_R _12701_ (.A(_05793_),
    .B(_05799_),
    .C(_05804_),
    .Y(_05805_));
 OR3x1_ASAP7_75t_R _12702_ (.A(_04486_),
    .B(_05792_),
    .C(_05805_),
    .Y(_05806_));
 AND2x2_ASAP7_75t_R _12703_ (.A(_05272_),
    .B(_00730_),
    .Y(_05807_));
 AO21x1_ASAP7_75t_R _12704_ (.A1(_03082_),
    .A2(_00729_),
    .B(_05807_),
    .Y(_05808_));
 AND3x1_ASAP7_75t_R _12705_ (.A(_05266_),
    .B(_03145_),
    .C(_00728_),
    .Y(_05809_));
 AO21x1_ASAP7_75t_R _12706_ (.A1(_00727_),
    .A2(_05787_),
    .B(_05809_),
    .Y(_05810_));
 AO221x1_ASAP7_75t_R _12707_ (.A1(_05410_),
    .A2(_05808_),
    .B1(_05810_),
    .B2(_05790_),
    .C(_05077_),
    .Y(_05811_));
 AND2x2_ASAP7_75t_R _12708_ (.A(_03674_),
    .B(_00725_),
    .Y(_05812_));
 AO21x1_ASAP7_75t_R _12709_ (.A1(_03161_),
    .A2(_00723_),
    .B(_05812_),
    .Y(_05813_));
 BUFx6f_ASAP7_75t_R _12710_ (.A(_03905_),
    .Y(_05814_));
 AO21x1_ASAP7_75t_R _12711_ (.A1(_00724_),
    .A2(_04861_),
    .B(_04862_),
    .Y(_05815_));
 AO221x1_ASAP7_75t_R _12712_ (.A1(_00726_),
    .A2(_04413_),
    .B1(_05813_),
    .B2(_05814_),
    .C(_05815_),
    .Y(_05816_));
 AND3x1_ASAP7_75t_R _12713_ (.A(_05793_),
    .B(_05811_),
    .C(_05816_),
    .Y(_05817_));
 AND2x2_ASAP7_75t_R _12714_ (.A(_05044_),
    .B(_00722_),
    .Y(_05818_));
 AO21x1_ASAP7_75t_R _12715_ (.A1(_04095_),
    .A2(_00721_),
    .B(_05818_),
    .Y(_05819_));
 AND3x1_ASAP7_75t_R _12716_ (.A(_05266_),
    .B(_03145_),
    .C(_00720_),
    .Y(_05820_));
 AO21x1_ASAP7_75t_R _12717_ (.A1(_00719_),
    .A2(_05787_),
    .B(_05820_),
    .Y(_05821_));
 AO221x1_ASAP7_75t_R _12718_ (.A1(_05410_),
    .A2(_05819_),
    .B1(_05821_),
    .B2(_05790_),
    .C(_05798_),
    .Y(_05822_));
 AND2x2_ASAP7_75t_R _12719_ (.A(_03087_),
    .B(_00717_),
    .Y(_05823_));
 AO21x1_ASAP7_75t_R _12720_ (.A1(_03161_),
    .A2(_00715_),
    .B(_05823_),
    .Y(_05824_));
 AO21x1_ASAP7_75t_R _12721_ (.A1(_00716_),
    .A2(_04861_),
    .B(_04862_),
    .Y(_05825_));
 AO221x1_ASAP7_75t_R _12722_ (.A1(_00718_),
    .A2(_04413_),
    .B1(_05824_),
    .B2(_05814_),
    .C(_05825_),
    .Y(_05826_));
 AND3x1_ASAP7_75t_R _12723_ (.A(_05034_),
    .B(_05822_),
    .C(_05826_),
    .Y(_05827_));
 OR3x1_ASAP7_75t_R _12724_ (.A(_04423_),
    .B(_05817_),
    .C(_05827_),
    .Y(_05828_));
 AO21x2_ASAP7_75t_R _12725_ (.A1(_05806_),
    .A2(_05828_),
    .B(_04163_),
    .Y(_05829_));
 NAND2x1_ASAP7_75t_R _12726_ (.A(_04422_),
    .B(_05829_),
    .Y(_05830_));
 OA21x2_ASAP7_75t_R _12727_ (.A1(_04159_),
    .A2(_09738_),
    .B(_05830_),
    .Y(_05831_));
 XNOR2x1_ASAP7_75t_R _12728_ (.B(_05831_),
    .Y(_09661_),
    .A(_03259_));
 INVx1_ASAP7_75t_R _12729_ (.A(_09661_),
    .Y(_09663_));
 OA22x2_ASAP7_75t_R _12730_ (.A1(_00712_),
    .A2(_03847_),
    .B1(_03400_),
    .B2(_00711_),
    .Y(_05832_));
 OA211x2_ASAP7_75t_R _12731_ (.A1(_03273_),
    .A2(_03287_),
    .B(_04444_),
    .C(_05832_),
    .Y(_05833_));
 AND2x2_ASAP7_75t_R _12732_ (.A(_00708_),
    .B(_03454_),
    .Y(_05834_));
 AND2x2_ASAP7_75t_R _12733_ (.A(_00707_),
    .B(_03740_),
    .Y(_05835_));
 OA21x2_ASAP7_75t_R _12734_ (.A1(_05834_),
    .A2(_05835_),
    .B(_03394_),
    .Y(_05836_));
 OA211x2_ASAP7_75t_R _12735_ (.A1(_05833_),
    .A2(_05836_),
    .B(_04786_),
    .C(_03888_),
    .Y(_05837_));
 OA22x2_ASAP7_75t_R _12736_ (.A1(_00703_),
    .A2(_04896_),
    .B1(_04451_),
    .B2(_00704_),
    .Y(_05838_));
 AND3x1_ASAP7_75t_R _12737_ (.A(_05440_),
    .B(_03835_),
    .C(_05838_),
    .Y(_05839_));
 OA21x2_ASAP7_75t_R _12738_ (.A1(_00700_),
    .A2(_05557_),
    .B(_03421_),
    .Y(_05840_));
 OR4x2_ASAP7_75t_R _12739_ (.A(_05032_),
    .B(_05837_),
    .C(_05839_),
    .D(_05840_),
    .Y(_05841_));
 BUFx6f_ASAP7_75t_R _12740_ (.A(_04018_),
    .Y(_05842_));
 OAI22x1_ASAP7_75t_R _12741_ (.A1(_00701_),
    .A2(_05248_),
    .B1(_05557_),
    .B2(_00702_),
    .Y(_05843_));
 OAI22x1_ASAP7_75t_R _12742_ (.A1(_00705_),
    .A2(_05248_),
    .B1(_05557_),
    .B2(_00706_),
    .Y(_05844_));
 AO32x1_ASAP7_75t_R _12743_ (.A1(_03210_),
    .A2(_05842_),
    .A3(_05843_),
    .B1(_05844_),
    .B2(_05440_),
    .Y(_05845_));
 OA22x2_ASAP7_75t_R _12744_ (.A1(_00709_),
    .A2(_05248_),
    .B1(_05557_),
    .B2(_00710_),
    .Y(_05846_));
 BUFx10_ASAP7_75t_R _12745_ (.A(_03432_),
    .Y(_05847_));
 OA222x2_ASAP7_75t_R _12746_ (.A1(_00713_),
    .A2(_04440_),
    .B1(_05847_),
    .B2(_00714_),
    .C1(_03278_),
    .C2(_05314_),
    .Y(_05848_));
 AOI211x1_ASAP7_75t_R _12747_ (.A1(_05318_),
    .A2(_05846_),
    .B(_05848_),
    .C(_03300_),
    .Y(_05849_));
 AOI211x1_ASAP7_75t_R _12748_ (.A1(_03300_),
    .A2(_05845_),
    .B(_05849_),
    .C(_04214_),
    .Y(_05850_));
 AND2x2_ASAP7_75t_R _12749_ (.A(_00723_),
    .B(_03451_),
    .Y(_05851_));
 AOI21x1_ASAP7_75t_R _12750_ (.A1(_00724_),
    .A2(_04882_),
    .B(_05851_),
    .Y(_05852_));
 OAI22x1_ASAP7_75t_R _12751_ (.A1(_00728_),
    .A2(_03377_),
    .B1(_03455_),
    .B2(_00727_),
    .Y(_05853_));
 OA211x2_ASAP7_75t_R _12752_ (.A1(_03284_),
    .A2(_03288_),
    .B(_05127_),
    .C(_05853_),
    .Y(_05854_));
 AO21x1_ASAP7_75t_R _12753_ (.A1(_05444_),
    .A2(_05852_),
    .B(_05854_),
    .Y(_05855_));
 AND2x2_ASAP7_75t_R _12754_ (.A(_00715_),
    .B(_03451_),
    .Y(_05856_));
 AOI21x1_ASAP7_75t_R _12755_ (.A1(_00716_),
    .A2(_04882_),
    .B(_05856_),
    .Y(_05857_));
 OAI22x1_ASAP7_75t_R _12756_ (.A1(_00719_),
    .A2(_04896_),
    .B1(_04451_),
    .B2(_00720_),
    .Y(_05858_));
 OA211x2_ASAP7_75t_R _12757_ (.A1(_03284_),
    .A2(_03288_),
    .B(_05127_),
    .C(_05858_),
    .Y(_05859_));
 AO21x1_ASAP7_75t_R _12758_ (.A1(_05444_),
    .A2(_05857_),
    .B(_05859_),
    .Y(_05860_));
 OAI22x1_ASAP7_75t_R _12759_ (.A1(_05102_),
    .A2(_05855_),
    .B1(_05860_),
    .B2(_04348_),
    .Y(_05861_));
 OA22x2_ASAP7_75t_R _12760_ (.A1(_00717_),
    .A2(_05227_),
    .B1(_03451_),
    .B2(_00718_),
    .Y(_05862_));
 OA22x2_ASAP7_75t_R _12761_ (.A1(_00721_),
    .A2(_03306_),
    .B1(_03450_),
    .B2(_00722_),
    .Y(_05863_));
 OA211x2_ASAP7_75t_R _12762_ (.A1(_03284_),
    .A2(_03288_),
    .B(_03472_),
    .C(_05863_),
    .Y(_05864_));
 AO221x1_ASAP7_75t_R _12763_ (.A1(_03412_),
    .A2(_04899_),
    .B1(_05444_),
    .B2(_05862_),
    .C(_05864_),
    .Y(_05865_));
 OR2x2_ASAP7_75t_R _12764_ (.A(_00726_),
    .B(_03414_),
    .Y(_05866_));
 OA211x2_ASAP7_75t_R _12765_ (.A1(_00725_),
    .A2(_04896_),
    .B(_05866_),
    .C(_03394_),
    .Y(_05867_));
 OA222x2_ASAP7_75t_R _12766_ (.A1(_00729_),
    .A2(_04896_),
    .B1(_04451_),
    .B2(_00730_),
    .C1(_03278_),
    .C2(_05314_),
    .Y(_05868_));
 OR3x1_ASAP7_75t_R _12767_ (.A(_03406_),
    .B(_05867_),
    .C(_05868_),
    .Y(_05869_));
 AO31x2_ASAP7_75t_R _12768_ (.A1(_03444_),
    .A2(_05865_),
    .A3(_05869_),
    .B(_04003_),
    .Y(_05870_));
 OAI22x1_ASAP7_75t_R _12769_ (.A1(_05841_),
    .A2(_05850_),
    .B1(_05861_),
    .B2(_05870_),
    .Y(_05871_));
 BUFx6f_ASAP7_75t_R _12770_ (.A(_05871_),
    .Y(_09660_));
 INVx1_ASAP7_75t_R _12771_ (.A(_09660_),
    .Y(_09662_));
 AND2x2_ASAP7_75t_R _12772_ (.A(_04390_),
    .B(_00735_),
    .Y(_05872_));
 AO21x1_ASAP7_75t_R _12773_ (.A1(_04851_),
    .A2(_00734_),
    .B(_05872_),
    .Y(_05873_));
 AO21x1_ASAP7_75t_R _12774_ (.A1(_04850_),
    .A2(_05873_),
    .B(_03078_),
    .Y(_05874_));
 AO22x1_ASAP7_75t_R _12775_ (.A1(_03112_),
    .A2(_00732_),
    .B1(_00733_),
    .B2(_03906_),
    .Y(_05875_));
 AO22x1_ASAP7_75t_R _12776_ (.A1(_03131_),
    .A2(_00732_),
    .B1(_05875_),
    .B2(_04381_),
    .Y(_05876_));
 AO21x1_ASAP7_75t_R _12777_ (.A1(_03216_),
    .A2(_05874_),
    .B(_05876_),
    .Y(_05877_));
 AND2x2_ASAP7_75t_R _12778_ (.A(_05044_),
    .B(_00739_),
    .Y(_05878_));
 AO21x1_ASAP7_75t_R _12779_ (.A1(_04095_),
    .A2(_00738_),
    .B(_05878_),
    .Y(_05879_));
 AND3x1_ASAP7_75t_R _12780_ (.A(_05272_),
    .B(_03145_),
    .C(_00737_),
    .Y(_05880_));
 AO21x1_ASAP7_75t_R _12781_ (.A1(_00736_),
    .A2(_05787_),
    .B(_05880_),
    .Y(_05881_));
 AO221x1_ASAP7_75t_R _12782_ (.A1(_05410_),
    .A2(_05879_),
    .B1(_05881_),
    .B2(_05790_),
    .C(_05798_),
    .Y(_05882_));
 AND3x1_ASAP7_75t_R _12783_ (.A(_05034_),
    .B(_05877_),
    .C(_05882_),
    .Y(_05883_));
 AND2x2_ASAP7_75t_R _12784_ (.A(_03092_),
    .B(_00747_),
    .Y(_05884_));
 AO21x1_ASAP7_75t_R _12785_ (.A1(_04095_),
    .A2(_00746_),
    .B(_05884_),
    .Y(_05885_));
 AND3x1_ASAP7_75t_R _12786_ (.A(_05272_),
    .B(_03145_),
    .C(_00745_),
    .Y(_05886_));
 AO21x1_ASAP7_75t_R _12787_ (.A1(_00744_),
    .A2(_05787_),
    .B(_05886_),
    .Y(_05887_));
 AO221x1_ASAP7_75t_R _12788_ (.A1(_05041_),
    .A2(_05885_),
    .B1(_05887_),
    .B2(_04856_),
    .C(_05798_),
    .Y(_05888_));
 AO22x1_ASAP7_75t_R _12789_ (.A1(_03139_),
    .A2(_00740_),
    .B1(_00741_),
    .B2(_04513_),
    .Y(_05889_));
 AND2x2_ASAP7_75t_R _12790_ (.A(_04390_),
    .B(_00743_),
    .Y(_05890_));
 AO21x1_ASAP7_75t_R _12791_ (.A1(_04851_),
    .A2(_00742_),
    .B(_05890_),
    .Y(_05891_));
 AO21x1_ASAP7_75t_R _12792_ (.A1(_04850_),
    .A2(_05891_),
    .B(_03078_),
    .Y(_05892_));
 AO21x1_ASAP7_75t_R _12793_ (.A1(_03137_),
    .A2(_05889_),
    .B(_05892_),
    .Y(_05893_));
 AND3x1_ASAP7_75t_R _12794_ (.A(_05793_),
    .B(_05888_),
    .C(_05893_),
    .Y(_05894_));
 OR3x1_ASAP7_75t_R _12795_ (.A(_04486_),
    .B(_05883_),
    .C(_05894_),
    .Y(_05895_));
 AND2x2_ASAP7_75t_R _12796_ (.A(_05044_),
    .B(_00763_),
    .Y(_05896_));
 AO21x1_ASAP7_75t_R _12797_ (.A1(_04095_),
    .A2(_00762_),
    .B(_05896_),
    .Y(_05897_));
 AND3x1_ASAP7_75t_R _12798_ (.A(_05272_),
    .B(_03145_),
    .C(_00761_),
    .Y(_05898_));
 AO21x1_ASAP7_75t_R _12799_ (.A1(_00760_),
    .A2(_05787_),
    .B(_05898_),
    .Y(_05899_));
 AO221x1_ASAP7_75t_R _12800_ (.A1(_05410_),
    .A2(_05897_),
    .B1(_05899_),
    .B2(_05790_),
    .C(_05798_),
    .Y(_05900_));
 AND2x2_ASAP7_75t_R _12801_ (.A(_03087_),
    .B(_00758_),
    .Y(_05901_));
 AO21x1_ASAP7_75t_R _12802_ (.A1(_03161_),
    .A2(_00756_),
    .B(_05901_),
    .Y(_05902_));
 AO21x1_ASAP7_75t_R _12803_ (.A1(_00757_),
    .A2(_04861_),
    .B(_04862_),
    .Y(_05903_));
 AO221x1_ASAP7_75t_R _12804_ (.A1(_00759_),
    .A2(_04413_),
    .B1(_05902_),
    .B2(_05814_),
    .C(_05903_),
    .Y(_05904_));
 AND3x1_ASAP7_75t_R _12805_ (.A(_05793_),
    .B(_05900_),
    .C(_05904_),
    .Y(_05905_));
 AND2x2_ASAP7_75t_R _12806_ (.A(_03092_),
    .B(_00755_),
    .Y(_05906_));
 AO21x1_ASAP7_75t_R _12807_ (.A1(_04095_),
    .A2(_00754_),
    .B(_05906_),
    .Y(_05907_));
 AND3x1_ASAP7_75t_R _12808_ (.A(_05272_),
    .B(_03145_),
    .C(_00753_),
    .Y(_05908_));
 AO21x1_ASAP7_75t_R _12809_ (.A1(_00752_),
    .A2(_05787_),
    .B(_05908_),
    .Y(_05909_));
 AO221x1_ASAP7_75t_R _12810_ (.A1(_05041_),
    .A2(_05907_),
    .B1(_05909_),
    .B2(_04856_),
    .C(_05798_),
    .Y(_05910_));
 AND2x2_ASAP7_75t_R _12811_ (.A(_03087_),
    .B(_00750_),
    .Y(_05911_));
 AO21x1_ASAP7_75t_R _12812_ (.A1(_03161_),
    .A2(_00748_),
    .B(_05911_),
    .Y(_05912_));
 AO21x1_ASAP7_75t_R _12813_ (.A1(_00749_),
    .A2(_04861_),
    .B(_04862_),
    .Y(_05913_));
 AO221x1_ASAP7_75t_R _12814_ (.A1(_00751_),
    .A2(_04413_),
    .B1(_05912_),
    .B2(_05814_),
    .C(_05913_),
    .Y(_05914_));
 AND3x1_ASAP7_75t_R _12815_ (.A(_05034_),
    .B(_05910_),
    .C(_05914_),
    .Y(_05915_));
 OR3x1_ASAP7_75t_R _12816_ (.A(_04423_),
    .B(_05905_),
    .C(_05915_),
    .Y(_05916_));
 AO21x2_ASAP7_75t_R _12817_ (.A1(_05895_),
    .A2(_05916_),
    .B(_04163_),
    .Y(_05917_));
 AND3x2_ASAP7_75t_R _12818_ (.A(net89),
    .B(net22),
    .C(_03777_),
    .Y(_09736_));
 NAND2x1_ASAP7_75t_R _12819_ (.A(_03707_),
    .B(_09736_),
    .Y(_05918_));
 OA21x2_ASAP7_75t_R _12820_ (.A1(_03780_),
    .A2(_05917_),
    .B(_05918_),
    .Y(_05919_));
 XNOR2x1_ASAP7_75t_R _12821_ (.B(_05919_),
    .Y(_09666_),
    .A(_03556_));
 INVx1_ASAP7_75t_R _12822_ (.A(_09666_),
    .Y(_09668_));
 AND2x2_ASAP7_75t_R _12823_ (.A(_00749_),
    .B(_03401_),
    .Y(_05920_));
 AO21x1_ASAP7_75t_R _12824_ (.A1(_00748_),
    .A2(_05557_),
    .B(_05920_),
    .Y(_05921_));
 OA22x2_ASAP7_75t_R _12825_ (.A1(_00752_),
    .A2(_03429_),
    .B1(_03432_),
    .B2(_00753_),
    .Y(_05922_));
 OA211x2_ASAP7_75t_R _12826_ (.A1(_03284_),
    .A2(_03288_),
    .B(_04885_),
    .C(_05922_),
    .Y(_05923_));
 AO21x1_ASAP7_75t_R _12827_ (.A1(_05444_),
    .A2(_05921_),
    .B(_05923_),
    .Y(_05924_));
 OA22x2_ASAP7_75t_R _12828_ (.A1(_00750_),
    .A2(_03350_),
    .B1(_03383_),
    .B2(_00751_),
    .Y(_05925_));
 OA222x2_ASAP7_75t_R _12829_ (.A1(_00754_),
    .A2(_05106_),
    .B1(_04445_),
    .B2(_00755_),
    .C1(_03470_),
    .C2(_05314_),
    .Y(_05926_));
 AO21x1_ASAP7_75t_R _12830_ (.A1(_05318_),
    .A2(_05925_),
    .B(_05926_),
    .Y(_05927_));
 OA21x2_ASAP7_75t_R _12831_ (.A1(_04214_),
    .A2(_05927_),
    .B(_03406_),
    .Y(_05928_));
 OAI21x1_ASAP7_75t_R _12832_ (.A1(_03444_),
    .A2(_05924_),
    .B(_05928_),
    .Y(_05929_));
 AND2x2_ASAP7_75t_R _12833_ (.A(_00757_),
    .B(_03409_),
    .Y(_05930_));
 AO21x1_ASAP7_75t_R _12834_ (.A1(_00756_),
    .A2(_05241_),
    .B(_05930_),
    .Y(_05931_));
 OA22x2_ASAP7_75t_R _12835_ (.A1(_00761_),
    .A2(_03335_),
    .B1(_04132_),
    .B2(_00760_),
    .Y(_05932_));
 OA211x2_ASAP7_75t_R _12836_ (.A1(_03284_),
    .A2(_03288_),
    .B(_04885_),
    .C(_05932_),
    .Y(_05933_));
 AO221x1_ASAP7_75t_R _12837_ (.A1(_03412_),
    .A2(_05195_),
    .B1(_05444_),
    .B2(_05931_),
    .C(_05933_),
    .Y(_05934_));
 OA22x2_ASAP7_75t_R _12838_ (.A1(_00758_),
    .A2(_03350_),
    .B1(_03357_),
    .B2(_00759_),
    .Y(_05935_));
 OA222x2_ASAP7_75t_R _12839_ (.A1(_00762_),
    .A2(_05106_),
    .B1(_04445_),
    .B2(_00763_),
    .C1(_03470_),
    .C2(_05314_),
    .Y(_05936_));
 AO21x1_ASAP7_75t_R _12840_ (.A1(_05318_),
    .A2(_05935_),
    .B(_05936_),
    .Y(_05937_));
 OA21x2_ASAP7_75t_R _12841_ (.A1(_04214_),
    .A2(_05937_),
    .B(_04791_),
    .Y(_05938_));
 AOI21x1_ASAP7_75t_R _12842_ (.A1(_05934_),
    .A2(_05938_),
    .B(_04003_),
    .Y(_05939_));
 OAI22x1_ASAP7_75t_R _12843_ (.A1(_00745_),
    .A2(_03377_),
    .B1(_04768_),
    .B2(_00744_),
    .Y(_05940_));
 NAND2x1_ASAP7_75t_R _12844_ (.A(_03362_),
    .B(_05940_),
    .Y(_05941_));
 OA22x2_ASAP7_75t_R _12845_ (.A1(_00742_),
    .A2(_03429_),
    .B1(_03432_),
    .B2(_00743_),
    .Y(_05942_));
 OA222x2_ASAP7_75t_R _12846_ (.A1(_00746_),
    .A2(_04560_),
    .B1(_04005_),
    .B2(_00747_),
    .C1(_03470_),
    .C2(_03468_),
    .Y(_05943_));
 AO221x1_ASAP7_75t_R _12847_ (.A1(_03326_),
    .A2(_03988_),
    .B1(_03394_),
    .B2(_05942_),
    .C(_05943_),
    .Y(_05944_));
 AO21x1_ASAP7_75t_R _12848_ (.A1(_05941_),
    .A2(_05944_),
    .B(_03345_),
    .Y(_05945_));
 AND2x2_ASAP7_75t_R _12849_ (.A(_00741_),
    .B(_03401_),
    .Y(_05946_));
 AO21x1_ASAP7_75t_R _12850_ (.A1(_00740_),
    .A2(_05847_),
    .B(_05946_),
    .Y(_05947_));
 OA21x2_ASAP7_75t_R _12851_ (.A1(_04450_),
    .A2(_05947_),
    .B(_04791_),
    .Y(_05948_));
 OAI22x1_ASAP7_75t_R _12852_ (.A1(_00736_),
    .A2(_05227_),
    .B1(_05241_),
    .B2(_00737_),
    .Y(_05949_));
 NAND2x1_ASAP7_75t_R _12853_ (.A(_03362_),
    .B(_05949_),
    .Y(_05950_));
 OA22x2_ASAP7_75t_R _12854_ (.A1(_00734_),
    .A2(_04023_),
    .B1(_03432_),
    .B2(_00735_),
    .Y(_05951_));
 OA222x2_ASAP7_75t_R _12855_ (.A1(_00738_),
    .A2(_04560_),
    .B1(_03450_),
    .B2(_00739_),
    .C1(_03277_),
    .C2(_03468_),
    .Y(_05952_));
 AO221x1_ASAP7_75t_R _12856_ (.A1(_03326_),
    .A2(_03988_),
    .B1(_03394_),
    .B2(_05951_),
    .C(_05952_),
    .Y(_05953_));
 AO21x1_ASAP7_75t_R _12857_ (.A1(_05950_),
    .A2(_05953_),
    .B(_03345_),
    .Y(_05954_));
 AND2x2_ASAP7_75t_R _12858_ (.A(_00733_),
    .B(_03541_),
    .Y(_05955_));
 AO21x1_ASAP7_75t_R _12859_ (.A1(_00732_),
    .A2(_05847_),
    .B(_05955_),
    .Y(_05956_));
 OA21x2_ASAP7_75t_R _12860_ (.A1(_04450_),
    .A2(_05956_),
    .B(_03406_),
    .Y(_05957_));
 AOI22x1_ASAP7_75t_R _12861_ (.A1(_05945_),
    .A2(_05948_),
    .B1(_05954_),
    .B2(_05957_),
    .Y(_05958_));
 AO22x1_ASAP7_75t_R _12862_ (.A1(_05929_),
    .A2(_05939_),
    .B1(_05958_),
    .B2(_04484_),
    .Y(_05959_));
 BUFx6f_ASAP7_75t_R _12863_ (.A(_05959_),
    .Y(_09665_));
 INVx2_ASAP7_75t_R _12864_ (.A(_09665_),
    .Y(_09667_));
 AND2x2_ASAP7_75t_R _12865_ (.A(_03092_),
    .B(_00768_),
    .Y(_05960_));
 AO21x2_ASAP7_75t_R _12866_ (.A1(_04748_),
    .A2(_00767_),
    .B(_05960_),
    .Y(_05961_));
 AO21x1_ASAP7_75t_R _12867_ (.A1(_05041_),
    .A2(_05961_),
    .B(_05474_),
    .Y(_05962_));
 AO22x1_ASAP7_75t_R _12868_ (.A1(_03566_),
    .A2(_00765_),
    .B1(_00766_),
    .B2(_03906_),
    .Y(_05963_));
 AO22x1_ASAP7_75t_R _12869_ (.A1(_03131_),
    .A2(_00765_),
    .B1(_05963_),
    .B2(_03904_),
    .Y(_05964_));
 AO21x1_ASAP7_75t_R _12870_ (.A1(_03216_),
    .A2(_05962_),
    .B(_05964_),
    .Y(_05965_));
 AND2x2_ASAP7_75t_R _12871_ (.A(_05070_),
    .B(_00772_),
    .Y(_05966_));
 AO21x1_ASAP7_75t_R _12872_ (.A1(_04528_),
    .A2(_00771_),
    .B(_05966_),
    .Y(_05967_));
 AND3x1_ASAP7_75t_R _12873_ (.A(_03041_),
    .B(_03200_),
    .C(_00770_),
    .Y(_05968_));
 AO21x1_ASAP7_75t_R _12874_ (.A1(_00769_),
    .A2(_05073_),
    .B(_05968_),
    .Y(_05969_));
 AO221x1_ASAP7_75t_R _12875_ (.A1(_05069_),
    .A2(_05967_),
    .B1(_05969_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_05970_));
 AND3x1_ASAP7_75t_R _12876_ (.A(_05034_),
    .B(_05965_),
    .C(_05970_),
    .Y(_05971_));
 AND2x2_ASAP7_75t_R _12877_ (.A(_05070_),
    .B(_00780_),
    .Y(_05972_));
 AO21x1_ASAP7_75t_R _12878_ (.A1(_04528_),
    .A2(_00779_),
    .B(_05972_),
    .Y(_05973_));
 AND3x1_ASAP7_75t_R _12879_ (.A(_05070_),
    .B(_03200_),
    .C(_00778_),
    .Y(_05974_));
 AO21x1_ASAP7_75t_R _12880_ (.A1(_00777_),
    .A2(_05073_),
    .B(_05974_),
    .Y(_05975_));
 AO221x1_ASAP7_75t_R _12881_ (.A1(_05364_),
    .A2(_05973_),
    .B1(_05975_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_05976_));
 AO22x1_ASAP7_75t_R _12882_ (.A1(_04401_),
    .A2(_00773_),
    .B1(_00774_),
    .B2(_05370_),
    .Y(_05977_));
 AND2x2_ASAP7_75t_R _12883_ (.A(_03092_),
    .B(_00776_),
    .Y(_05978_));
 AO21x1_ASAP7_75t_R _12884_ (.A1(_04748_),
    .A2(_00775_),
    .B(_05978_),
    .Y(_05979_));
 AO21x1_ASAP7_75t_R _12885_ (.A1(_04850_),
    .A2(_05979_),
    .B(_05474_),
    .Y(_05980_));
 AO21x1_ASAP7_75t_R _12886_ (.A1(_05372_),
    .A2(_05977_),
    .B(_05980_),
    .Y(_05981_));
 AND3x1_ASAP7_75t_R _12887_ (.A(_05793_),
    .B(_05976_),
    .C(_05981_),
    .Y(_05982_));
 NOR3x1_ASAP7_75t_R _12888_ (.A(_04486_),
    .B(_05971_),
    .C(_05982_),
    .Y(_05983_));
 AND2x2_ASAP7_75t_R _12889_ (.A(_03071_),
    .B(_00796_),
    .Y(_05984_));
 AO21x1_ASAP7_75t_R _12890_ (.A1(_04860_),
    .A2(_00795_),
    .B(_05984_),
    .Y(_05985_));
 AND3x1_ASAP7_75t_R _12891_ (.A(_03049_),
    .B(_05229_),
    .C(_00794_),
    .Y(_05986_));
 AO21x1_ASAP7_75t_R _12892_ (.A1(_00793_),
    .A2(_05073_),
    .B(_05986_),
    .Y(_05987_));
 AO221x1_ASAP7_75t_R _12893_ (.A1(_05069_),
    .A2(_05985_),
    .B1(_05987_),
    .B2(_04764_),
    .C(_04657_),
    .Y(_05988_));
 AND2x2_ASAP7_75t_R _12894_ (.A(_04722_),
    .B(_00791_),
    .Y(_05989_));
 AO21x1_ASAP7_75t_R _12895_ (.A1(_03029_),
    .A2(_00789_),
    .B(_05989_),
    .Y(_05990_));
 AO21x1_ASAP7_75t_R _12896_ (.A1(_00790_),
    .A2(_05066_),
    .B(_05474_),
    .Y(_05991_));
 AO221x1_ASAP7_75t_R _12897_ (.A1(_00792_),
    .A2(_05061_),
    .B1(_05990_),
    .B2(_05375_),
    .C(_05991_),
    .Y(_05992_));
 AO21x1_ASAP7_75t_R _12898_ (.A1(_05988_),
    .A2(_05992_),
    .B(_04545_),
    .Y(_05993_));
 AND2x2_ASAP7_75t_R _12899_ (.A(_03049_),
    .B(_00788_),
    .Y(_05994_));
 AO21x1_ASAP7_75t_R _12900_ (.A1(_04860_),
    .A2(_00787_),
    .B(_05994_),
    .Y(_05995_));
 AND3x1_ASAP7_75t_R _12901_ (.A(_03049_),
    .B(_05229_),
    .C(_00786_),
    .Y(_05996_));
 AO21x1_ASAP7_75t_R _12902_ (.A1(_00785_),
    .A2(_03291_),
    .B(_05996_),
    .Y(_05997_));
 AO221x1_ASAP7_75t_R _12903_ (.A1(_05069_),
    .A2(_05995_),
    .B1(_05997_),
    .B2(_04764_),
    .C(_04657_),
    .Y(_05998_));
 AND2x2_ASAP7_75t_R _12904_ (.A(_04722_),
    .B(_00783_),
    .Y(_05999_));
 AO21x1_ASAP7_75t_R _12905_ (.A1(_03029_),
    .A2(_00781_),
    .B(_05999_),
    .Y(_06000_));
 AO21x1_ASAP7_75t_R _12906_ (.A1(_00782_),
    .A2(_05066_),
    .B(_05474_),
    .Y(_06001_));
 AO221x1_ASAP7_75t_R _12907_ (.A1(_00784_),
    .A2(_05061_),
    .B1(_06000_),
    .B2(_05375_),
    .C(_06001_),
    .Y(_06002_));
 AO21x1_ASAP7_75t_R _12908_ (.A1(_05998_),
    .A2(_06002_),
    .B(_03175_),
    .Y(_06003_));
 AOI21x1_ASAP7_75t_R _12909_ (.A1(_05993_),
    .A2(_06003_),
    .B(_04423_),
    .Y(_06004_));
 OAI21x1_ASAP7_75t_R _12910_ (.A1(_05983_),
    .A2(_06004_),
    .B(_03705_),
    .Y(_06005_));
 AND3x2_ASAP7_75t_R _12911_ (.A(net89),
    .B(net20),
    .C(_03777_),
    .Y(_09734_));
 NAND2x1_ASAP7_75t_R _12912_ (.A(_03707_),
    .B(_09734_),
    .Y(_06006_));
 OA21x2_ASAP7_75t_R _12913_ (.A1(_03780_),
    .A2(_06005_),
    .B(_06006_),
    .Y(_06007_));
 XNOR2x1_ASAP7_75t_R _12914_ (.B(_06007_),
    .Y(_09671_),
    .A(_03556_));
 INVx1_ASAP7_75t_R _12915_ (.A(_09671_),
    .Y(_09673_));
 NAND2x1_ASAP7_75t_R _12916_ (.A(_00765_),
    .B(_03529_),
    .Y(_06008_));
 NAND2x1_ASAP7_75t_R _12917_ (.A(_00766_),
    .B(_04466_),
    .Y(_06009_));
 OAI22x1_ASAP7_75t_R _12918_ (.A1(_00769_),
    .A2(_04023_),
    .B1(_04005_),
    .B2(_00770_),
    .Y(_06010_));
 AO32x1_ASAP7_75t_R _12919_ (.A1(_03520_),
    .A2(_06008_),
    .A3(_06009_),
    .B1(_03516_),
    .B2(_06010_),
    .Y(_06011_));
 AND3x1_ASAP7_75t_R _12920_ (.A(_03117_),
    .B(_03970_),
    .C(_00772_),
    .Y(_06012_));
 AOI221x1_ASAP7_75t_R _12921_ (.A1(_03316_),
    .A2(_04460_),
    .B1(_03975_),
    .B2(_00771_),
    .C(_06012_),
    .Y(_06013_));
 INVx1_ASAP7_75t_R _12922_ (.A(_00768_),
    .Y(_06014_));
 OA211x2_ASAP7_75t_R _12923_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03327_),
    .C(_06014_),
    .Y(_06015_));
 NOR2x1_ASAP7_75t_R _12924_ (.A(_00767_),
    .B(_03348_),
    .Y(_06016_));
 OA211x2_ASAP7_75t_R _12925_ (.A1(_06015_),
    .A2(_06016_),
    .B(_03250_),
    .C(_03387_),
    .Y(_06017_));
 OA21x2_ASAP7_75t_R _12926_ (.A1(_06013_),
    .A2(_06017_),
    .B(_03340_),
    .Y(_06018_));
 OA21x2_ASAP7_75t_R _12927_ (.A1(_03997_),
    .A2(_06018_),
    .B(_03521_),
    .Y(_06019_));
 OR3x1_ASAP7_75t_R _12928_ (.A(_03096_),
    .B(_03749_),
    .C(_00776_),
    .Y(_06020_));
 OA22x2_ASAP7_75t_R _12929_ (.A1(_00775_),
    .A2(_03428_),
    .B1(_03748_),
    .B2(_06020_),
    .Y(_06021_));
 AND3x1_ASAP7_75t_R _12930_ (.A(_03860_),
    .B(_03970_),
    .C(_00780_),
    .Y(_06022_));
 AO221x1_ASAP7_75t_R _12931_ (.A1(_03316_),
    .A2(_03321_),
    .B1(_03975_),
    .B2(_00779_),
    .C(_06022_),
    .Y(_06023_));
 OA21x2_ASAP7_75t_R _12932_ (.A1(_04444_),
    .A2(_06021_),
    .B(_06023_),
    .Y(_06024_));
 AND2x2_ASAP7_75t_R _12933_ (.A(_00774_),
    .B(_03400_),
    .Y(_06025_));
 AO21x1_ASAP7_75t_R _12934_ (.A1(_00773_),
    .A2(_04445_),
    .B(_06025_),
    .Y(_06026_));
 OAI22x1_ASAP7_75t_R _12935_ (.A1(_04786_),
    .A2(_06024_),
    .B1(_06026_),
    .B2(_03411_),
    .Y(_06027_));
 OAI22x1_ASAP7_75t_R _12936_ (.A1(_00778_),
    .A2(_04480_),
    .B1(_03409_),
    .B2(_00777_),
    .Y(_06028_));
 AO21x1_ASAP7_75t_R _12937_ (.A1(_03540_),
    .A2(_06028_),
    .B(_03405_),
    .Y(_06029_));
 OA221x2_ASAP7_75t_R _12938_ (.A1(_06011_),
    .A2(_06019_),
    .B1(_06027_),
    .B2(_06029_),
    .C(_03498_),
    .Y(_06030_));
 OA22x2_ASAP7_75t_R _12939_ (.A1(_00794_),
    .A2(_03334_),
    .B1(_03408_),
    .B2(_00793_),
    .Y(_06031_));
 AO221x1_ASAP7_75t_R _12940_ (.A1(_04784_),
    .A2(_04783_),
    .B1(_04441_),
    .B2(_03325_),
    .C(_06031_),
    .Y(_06032_));
 AND2x2_ASAP7_75t_R _12941_ (.A(_00789_),
    .B(_03449_),
    .Y(_06033_));
 AND2x2_ASAP7_75t_R _12942_ (.A(_00790_),
    .B(_03408_),
    .Y(_06034_));
 OR3x1_ASAP7_75t_R _12943_ (.A(_03747_),
    .B(_06033_),
    .C(_06034_),
    .Y(_06035_));
 AND3x1_ASAP7_75t_R _12944_ (.A(_00791_),
    .B(_03250_),
    .C(_03736_),
    .Y(_06036_));
 AO221x1_ASAP7_75t_R _12945_ (.A1(_03064_),
    .A2(_05124_),
    .B1(_00795_),
    .B2(_03504_),
    .C(_06036_),
    .Y(_06037_));
 OR3x1_ASAP7_75t_R _12946_ (.A(_00792_),
    .B(_03359_),
    .C(_03485_),
    .Y(_06038_));
 OA211x2_ASAP7_75t_R _12947_ (.A1(_00796_),
    .A2(_03732_),
    .B(_06038_),
    .C(_03501_),
    .Y(_06039_));
 AO32x2_ASAP7_75t_R _12948_ (.A1(_03855_),
    .A2(_06032_),
    .A3(_06035_),
    .B1(_06037_),
    .B2(_06039_),
    .Y(_06040_));
 OA22x2_ASAP7_75t_R _12949_ (.A1(_00783_),
    .A2(_04022_),
    .B1(_04153_),
    .B2(_00784_),
    .Y(_06041_));
 AND2x2_ASAP7_75t_R _12950_ (.A(_00787_),
    .B(_03465_),
    .Y(_06042_));
 AO221x2_ASAP7_75t_R _12951_ (.A1(_03316_),
    .A2(_03321_),
    .B1(_03313_),
    .B2(_00788_),
    .C(_06042_),
    .Y(_06043_));
 OA21x2_ASAP7_75t_R _12952_ (.A1(_04444_),
    .A2(_06041_),
    .B(_06043_),
    .Y(_06044_));
 AO21x1_ASAP7_75t_R _12953_ (.A1(_04771_),
    .A2(_06044_),
    .B(_03836_),
    .Y(_06045_));
 OA22x2_ASAP7_75t_R _12954_ (.A1(_00785_),
    .A2(_04560_),
    .B1(_04005_),
    .B2(_00786_),
    .Y(_06046_));
 AND2x2_ASAP7_75t_R _12955_ (.A(_00782_),
    .B(_03467_),
    .Y(_06047_));
 AO21x1_ASAP7_75t_R _12956_ (.A1(_00781_),
    .A2(_03529_),
    .B(_06047_),
    .Y(_06048_));
 OA22x2_ASAP7_75t_R _12957_ (.A1(_04107_),
    .A2(_06046_),
    .B1(_06048_),
    .B2(_03845_),
    .Y(_06049_));
 AOI221x1_ASAP7_75t_R _12958_ (.A1(_04791_),
    .A2(_06040_),
    .B1(_06045_),
    .B2(_06049_),
    .C(_04003_),
    .Y(_06050_));
 OR2x2_ASAP7_75t_R _12959_ (.A(_06030_),
    .B(_06050_),
    .Y(_06051_));
 BUFx2_ASAP7_75t_R _12960_ (.A(_06051_),
    .Y(_09670_));
 INVx1_ASAP7_75t_R _12961_ (.A(_09670_),
    .Y(_09672_));
 AND2x2_ASAP7_75t_R _12962_ (.A(_04502_),
    .B(_00830_),
    .Y(_06052_));
 AO21x1_ASAP7_75t_R _12963_ (.A1(_03905_),
    .A2(_00829_),
    .B(_06052_),
    .Y(_06053_));
 AND3x1_ASAP7_75t_R _12964_ (.A(_03048_),
    .B(_03034_),
    .C(_00828_),
    .Y(_06054_));
 AO21x1_ASAP7_75t_R _12965_ (.A1(_00827_),
    .A2(_04393_),
    .B(_06054_),
    .Y(_06055_));
 AO221x1_ASAP7_75t_R _12966_ (.A1(_04389_),
    .A2(_06053_),
    .B1(_06055_),
    .B2(_04396_),
    .C(_05260_),
    .Y(_06056_));
 AND2x2_ASAP7_75t_R _12967_ (.A(_04502_),
    .B(_00822_),
    .Y(_06057_));
 AO21x1_ASAP7_75t_R _12968_ (.A1(_03112_),
    .A2(_00821_),
    .B(_06057_),
    .Y(_06058_));
 AND3x1_ASAP7_75t_R _12969_ (.A(_03048_),
    .B(_03034_),
    .C(_00820_),
    .Y(_06059_));
 AO21x1_ASAP7_75t_R _12970_ (.A1(_00819_),
    .A2(_04393_),
    .B(_06059_),
    .Y(_06060_));
 AO221x1_ASAP7_75t_R _12971_ (.A1(_04497_),
    .A2(_06058_),
    .B1(_06060_),
    .B2(_04396_),
    .C(_05253_),
    .Y(_06061_));
 AND3x1_ASAP7_75t_R _12972_ (.A(_03143_),
    .B(_06056_),
    .C(_06061_),
    .Y(_06062_));
 AND2x2_ASAP7_75t_R _12973_ (.A(_03806_),
    .B(_00817_),
    .Y(_06063_));
 AO21x1_ASAP7_75t_R _12974_ (.A1(_03589_),
    .A2(_00815_),
    .B(_06063_),
    .Y(_06064_));
 AO221x1_ASAP7_75t_R _12975_ (.A1(_03109_),
    .A2(_00818_),
    .B1(_05269_),
    .B2(_00816_),
    .C(_05153_),
    .Y(_06065_));
 OA211x2_ASAP7_75t_R _12976_ (.A1(_05366_),
    .A2(_06064_),
    .B(_06065_),
    .C(_03585_),
    .Y(_06066_));
 AND2x2_ASAP7_75t_R _12977_ (.A(_03806_),
    .B(_00825_),
    .Y(_06067_));
 AO21x1_ASAP7_75t_R _12978_ (.A1(_03589_),
    .A2(_00823_),
    .B(_06067_),
    .Y(_06068_));
 AO221x1_ASAP7_75t_R _12979_ (.A1(_03109_),
    .A2(_00826_),
    .B1(_05269_),
    .B2(_00824_),
    .C(_05153_),
    .Y(_06069_));
 OA211x2_ASAP7_75t_R _12980_ (.A1(_05366_),
    .A2(_06068_),
    .B(_06069_),
    .C(_03173_),
    .Y(_06070_));
 OR3x1_ASAP7_75t_R _12981_ (.A(_05067_),
    .B(_06066_),
    .C(_06070_),
    .Y(_06071_));
 AND2x2_ASAP7_75t_R _12982_ (.A(_03073_),
    .B(_00809_),
    .Y(_06072_));
 AO21x1_ASAP7_75t_R _12983_ (.A1(_03589_),
    .A2(_00807_),
    .B(_06072_),
    .Y(_06073_));
 AO21x1_ASAP7_75t_R _12984_ (.A1(_00810_),
    .A2(_03697_),
    .B(_03623_),
    .Y(_06074_));
 AO221x1_ASAP7_75t_R _12985_ (.A1(_00808_),
    .A2(_04861_),
    .B1(_06073_),
    .B2(_03139_),
    .C(_06074_),
    .Y(_06075_));
 AND2x2_ASAP7_75t_R _12986_ (.A(_03898_),
    .B(_00814_),
    .Y(_06076_));
 AO21x1_ASAP7_75t_R _12987_ (.A1(_03112_),
    .A2(_00813_),
    .B(_06076_),
    .Y(_06077_));
 AND3x1_ASAP7_75t_R _12988_ (.A(_03048_),
    .B(_03034_),
    .C(_00812_),
    .Y(_06078_));
 AO21x1_ASAP7_75t_R _12989_ (.A1(_00811_),
    .A2(_04393_),
    .B(_06078_),
    .Y(_06079_));
 AO221x1_ASAP7_75t_R _12990_ (.A1(_04497_),
    .A2(_06077_),
    .B1(_06079_),
    .B2(_03922_),
    .C(_04397_),
    .Y(_06080_));
 AND2x2_ASAP7_75t_R _12991_ (.A(_04488_),
    .B(_00802_),
    .Y(_06081_));
 AO21x1_ASAP7_75t_R _12992_ (.A1(_03062_),
    .A2(_00801_),
    .B(_06081_),
    .Y(_06082_));
 AO21x1_ASAP7_75t_R _12993_ (.A1(_04487_),
    .A2(_06082_),
    .B(_04416_),
    .Y(_06083_));
 AO22x1_ASAP7_75t_R _12994_ (.A1(_03573_),
    .A2(_00799_),
    .B1(_00800_),
    .B2(_03946_),
    .Y(_06084_));
 AO22x1_ASAP7_75t_R _12995_ (.A1(_04493_),
    .A2(_00799_),
    .B1(_06084_),
    .B2(_03028_),
    .Y(_06085_));
 AO21x1_ASAP7_75t_R _12996_ (.A1(_03201_),
    .A2(_06083_),
    .B(_06085_),
    .Y(_06086_));
 AND2x2_ASAP7_75t_R _12997_ (.A(_03675_),
    .B(_00806_),
    .Y(_06087_));
 AO21x1_ASAP7_75t_R _12998_ (.A1(_03625_),
    .A2(_00805_),
    .B(_06087_),
    .Y(_06088_));
 AND3x1_ASAP7_75t_R _12999_ (.A(_03678_),
    .B(_03117_),
    .C(_00804_),
    .Y(_06089_));
 AO21x1_ASAP7_75t_R _13000_ (.A1(_00803_),
    .A2(_03289_),
    .B(_06089_),
    .Y(_06090_));
 AO221x1_ASAP7_75t_R _13001_ (.A1(_03674_),
    .A2(_06088_),
    .B1(_06090_),
    .B2(_03681_),
    .C(_03636_),
    .Y(_06091_));
 AND2x2_ASAP7_75t_R _13002_ (.A(_03586_),
    .B(_06091_),
    .Y(_06092_));
 AO32x1_ASAP7_75t_R _13003_ (.A1(_03174_),
    .A2(_06075_),
    .A3(_06080_),
    .B1(_06086_),
    .B2(_06092_),
    .Y(_06093_));
 AO221x2_ASAP7_75t_R _13004_ (.A1(_06062_),
    .A2(_06071_),
    .B1(_06093_),
    .B2(_04100_),
    .C(_03127_),
    .Y(_06094_));
 AND3x2_ASAP7_75t_R _13005_ (.A(net89),
    .B(net19),
    .C(_03715_),
    .Y(_09732_));
 NAND2x1_ASAP7_75t_R _13006_ (.A(_03707_),
    .B(_09732_),
    .Y(_06095_));
 OA21x2_ASAP7_75t_R _13007_ (.A1(_03780_),
    .A2(_06094_),
    .B(_06095_),
    .Y(_06096_));
 XNOR2x1_ASAP7_75t_R _13008_ (.B(_06096_),
    .Y(_09676_),
    .A(_03556_));
 INVx1_ASAP7_75t_R _13009_ (.A(_09676_),
    .Y(_09678_));
 AND3x1_ASAP7_75t_R _13010_ (.A(_03215_),
    .B(_05335_),
    .C(_00814_),
    .Y(_06097_));
 AO21x1_ASAP7_75t_R _13011_ (.A1(_00813_),
    .A2(_04550_),
    .B(_06097_),
    .Y(_06098_));
 OA21x2_ASAP7_75t_R _13012_ (.A1(_00809_),
    .A2(_03329_),
    .B(_03388_),
    .Y(_06099_));
 OA21x2_ASAP7_75t_R _13013_ (.A1(_00810_),
    .A2(_04473_),
    .B(_06099_),
    .Y(_06100_));
 OA21x2_ASAP7_75t_R _13014_ (.A1(_03988_),
    .A2(_06100_),
    .B(_03210_),
    .Y(_06101_));
 AO21x1_ASAP7_75t_R _13015_ (.A1(_05093_),
    .A2(_06098_),
    .B(_06101_),
    .Y(_06102_));
 AND2x2_ASAP7_75t_R _13016_ (.A(_00808_),
    .B(_03409_),
    .Y(_06103_));
 AO21x1_ASAP7_75t_R _13017_ (.A1(_00807_),
    .A2(_03451_),
    .B(_06103_),
    .Y(_06104_));
 OAI22x1_ASAP7_75t_R _13018_ (.A1(_00812_),
    .A2(_03378_),
    .B1(_03479_),
    .B2(_00811_),
    .Y(_06105_));
 NAND2x1_ASAP7_75t_R _13019_ (.A(_03362_),
    .B(_06105_),
    .Y(_06106_));
 OA211x2_ASAP7_75t_R _13020_ (.A1(_04450_),
    .A2(_06104_),
    .B(_06106_),
    .C(_04791_),
    .Y(_06107_));
 OR3x1_ASAP7_75t_R _13021_ (.A(_04493_),
    .B(_04561_),
    .C(_00806_),
    .Y(_06108_));
 OR3x1_ASAP7_75t_R _13022_ (.A(_00802_),
    .B(_03468_),
    .C(_03722_),
    .Y(_06109_));
 OA211x2_ASAP7_75t_R _13023_ (.A1(_05318_),
    .A2(_06108_),
    .B(_06109_),
    .C(_04771_),
    .Y(_06110_));
 AND3x1_ASAP7_75t_R _13024_ (.A(_00801_),
    .B(_03317_),
    .C(_03322_),
    .Y(_06111_));
 AO221x1_ASAP7_75t_R _13025_ (.A1(_03201_),
    .A2(_05335_),
    .B1(_00805_),
    .B2(_04885_),
    .C(_06111_),
    .Y(_06112_));
 AO21x2_ASAP7_75t_R _13026_ (.A1(_06110_),
    .A2(_06112_),
    .B(_04458_),
    .Y(_06113_));
 OA22x2_ASAP7_75t_R _13027_ (.A1(_00803_),
    .A2(_05227_),
    .B1(_03451_),
    .B2(_00804_),
    .Y(_06114_));
 AND2x2_ASAP7_75t_R _13028_ (.A(_00800_),
    .B(_03541_),
    .Y(_06115_));
 AO21x1_ASAP7_75t_R _13029_ (.A1(_00799_),
    .A2(_05241_),
    .B(_06115_),
    .Y(_06116_));
 OA22x2_ASAP7_75t_R _13030_ (.A1(_04107_),
    .A2(_06114_),
    .B1(_06116_),
    .B2(_04450_),
    .Y(_06117_));
 AOI22x1_ASAP7_75t_R _13031_ (.A1(_06102_),
    .A2(_06107_),
    .B1(_06113_),
    .B2(_06117_),
    .Y(_06118_));
 INVx1_ASAP7_75t_R _13032_ (.A(_00815_),
    .Y(_06119_));
 NAND2x1_ASAP7_75t_R _13033_ (.A(_00816_),
    .B(_03455_),
    .Y(_06120_));
 OA211x2_ASAP7_75t_R _13034_ (.A1(_06119_),
    .A2(_03410_),
    .B(_03448_),
    .C(_06120_),
    .Y(_06121_));
 NOR2x1_ASAP7_75t_R _13035_ (.A(_00817_),
    .B(_03428_),
    .Y(_06122_));
 INVx1_ASAP7_75t_R _13036_ (.A(_00818_),
    .Y(_06123_));
 OA211x2_ASAP7_75t_R _13037_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03328_),
    .C(_06123_),
    .Y(_06124_));
 OA211x2_ASAP7_75t_R _13038_ (.A1(_06122_),
    .A2(_06124_),
    .B(_03325_),
    .C(_04441_),
    .Y(_06125_));
 AND2x2_ASAP7_75t_R _13039_ (.A(_00821_),
    .B(_03466_),
    .Y(_06126_));
 AOI221x1_ASAP7_75t_R _13040_ (.A1(_03317_),
    .A2(_04020_),
    .B1(_04023_),
    .B2(_00822_),
    .C(_06126_),
    .Y(_06127_));
 OA21x2_ASAP7_75t_R _13041_ (.A1(_06125_),
    .A2(_06127_),
    .B(_04026_),
    .Y(_06128_));
 OR3x1_ASAP7_75t_R _13042_ (.A(_03597_),
    .B(_04561_),
    .C(_00820_),
    .Y(_06129_));
 OAI22x1_ASAP7_75t_R _13043_ (.A1(_00819_),
    .A2(_05106_),
    .B1(_03748_),
    .B2(_06129_),
    .Y(_06130_));
 AO21x1_ASAP7_75t_R _13044_ (.A1(_03457_),
    .A2(_06130_),
    .B(_03461_),
    .Y(_06131_));
 OA21x2_ASAP7_75t_R _13045_ (.A1(_06128_),
    .A2(_06131_),
    .B(_03412_),
    .Y(_06132_));
 INVx1_ASAP7_75t_R _13046_ (.A(_00825_),
    .Y(_06133_));
 INVx1_ASAP7_75t_R _13047_ (.A(_00826_),
    .Y(_06134_));
 AO221x1_ASAP7_75t_R _13048_ (.A1(_06133_),
    .A2(_03466_),
    .B1(_03467_),
    .B2(_06134_),
    .C(_03468_),
    .Y(_06135_));
 AO21x1_ASAP7_75t_R _13049_ (.A1(_03382_),
    .A2(_06135_),
    .B(_03470_),
    .Y(_06136_));
 AND3x1_ASAP7_75t_R _13050_ (.A(_03473_),
    .B(_03475_),
    .C(_00830_),
    .Y(_06137_));
 AO21x1_ASAP7_75t_R _13051_ (.A1(_00829_),
    .A2(_03437_),
    .B(_06137_),
    .Y(_06138_));
 NAND2x1_ASAP7_75t_R _13052_ (.A(_03472_),
    .B(_06138_),
    .Y(_06139_));
 OAI22x1_ASAP7_75t_R _13053_ (.A1(_00828_),
    .A2(_03378_),
    .B1(_03479_),
    .B2(_00827_),
    .Y(_06140_));
 OA211x2_ASAP7_75t_R _13054_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03313_),
    .C(_00824_),
    .Y(_06141_));
 AOI21x1_ASAP7_75t_R _13055_ (.A1(_00823_),
    .A2(_03529_),
    .B(_06141_),
    .Y(_06142_));
 AO21x1_ASAP7_75t_R _13056_ (.A1(_03484_),
    .A2(_06142_),
    .B(_03299_),
    .Y(_06143_));
 AO221x1_ASAP7_75t_R _13057_ (.A1(_06136_),
    .A2(_06139_),
    .B1(_06140_),
    .B2(_04891_),
    .C(_06143_),
    .Y(_06144_));
 OA211x2_ASAP7_75t_R _13058_ (.A1(_06121_),
    .A2(_06132_),
    .B(_06144_),
    .C(_03495_),
    .Y(_06145_));
 AO21x1_ASAP7_75t_R _13059_ (.A1(_04484_),
    .A2(_06118_),
    .B(_06145_),
    .Y(_06146_));
 BUFx3_ASAP7_75t_R _13060_ (.A(_06146_),
    .Y(_09675_));
 INVx1_ASAP7_75t_R _13061_ (.A(_09675_),
    .Y(_09677_));
 AND2x2_ASAP7_75t_R _13062_ (.A(_04390_),
    .B(_00839_),
    .Y(_06147_));
 AO21x1_ASAP7_75t_R _13063_ (.A1(_03566_),
    .A2(_00838_),
    .B(_06147_),
    .Y(_06148_));
 AND3x1_ASAP7_75t_R _13064_ (.A(_04408_),
    .B(_03149_),
    .C(_00837_),
    .Y(_06149_));
 AO21x1_ASAP7_75t_R _13065_ (.A1(_00836_),
    .A2(_03290_),
    .B(_06149_),
    .Y(_06150_));
 AO221x2_ASAP7_75t_R _13066_ (.A1(_04389_),
    .A2(_06148_),
    .B1(_06150_),
    .B2(_04396_),
    .C(_04397_),
    .Y(_06151_));
 AO22x1_ASAP7_75t_R _13067_ (.A1(_04748_),
    .A2(_00832_),
    .B1(_00833_),
    .B2(_04513_),
    .Y(_06152_));
 AND2x2_ASAP7_75t_R _13068_ (.A(_04267_),
    .B(_00835_),
    .Y(_06153_));
 AO21x2_ASAP7_75t_R _13069_ (.A1(_03945_),
    .A2(_00834_),
    .B(_06153_),
    .Y(_06154_));
 AO221x1_ASAP7_75t_R _13070_ (.A1(_04493_),
    .A2(_00832_),
    .B1(_03925_),
    .B2(_06154_),
    .C(_03914_),
    .Y(_06155_));
 AO21x1_ASAP7_75t_R _13071_ (.A1(_03137_),
    .A2(_06152_),
    .B(_06155_),
    .Y(_06156_));
 AND3x1_ASAP7_75t_R _13072_ (.A(_03703_),
    .B(_06151_),
    .C(_06156_),
    .Y(_06157_));
 AND2x2_ASAP7_75t_R _13073_ (.A(_04390_),
    .B(_00855_),
    .Y(_06158_));
 AO21x1_ASAP7_75t_R _13074_ (.A1(_03566_),
    .A2(_00854_),
    .B(_06158_),
    .Y(_06159_));
 AND3x1_ASAP7_75t_R _13075_ (.A(_04390_),
    .B(_03149_),
    .C(_00853_),
    .Y(_06160_));
 AO21x1_ASAP7_75t_R _13076_ (.A1(_00852_),
    .A2(_04393_),
    .B(_06160_),
    .Y(_06161_));
 AO221x1_ASAP7_75t_R _13077_ (.A1(_04389_),
    .A2(_06159_),
    .B1(_06161_),
    .B2(_04396_),
    .C(_04397_),
    .Y(_06162_));
 AND2x2_ASAP7_75t_R _13078_ (.A(_03806_),
    .B(_00850_),
    .Y(_06163_));
 AO21x1_ASAP7_75t_R _13079_ (.A1(_03028_),
    .A2(_00848_),
    .B(_06163_),
    .Y(_06164_));
 AO21x1_ASAP7_75t_R _13080_ (.A1(_00849_),
    .A2(_03561_),
    .B(_04416_),
    .Y(_06165_));
 AO221x1_ASAP7_75t_R _13081_ (.A1(_00851_),
    .A2(_04413_),
    .B1(_06164_),
    .B2(_04401_),
    .C(_06165_),
    .Y(_06166_));
 AND3x1_ASAP7_75t_R _13082_ (.A(_03143_),
    .B(_06162_),
    .C(_06166_),
    .Y(_06167_));
 OR4x1_ASAP7_75t_R _13083_ (.A(_03175_),
    .B(_03781_),
    .C(_06157_),
    .D(_06167_),
    .Y(_06168_));
 AND2x2_ASAP7_75t_R _13084_ (.A(_03092_),
    .B(_00847_),
    .Y(_06169_));
 AO21x1_ASAP7_75t_R _13085_ (.A1(_04080_),
    .A2(_00846_),
    .B(_06169_),
    .Y(_06170_));
 AND3x1_ASAP7_75t_R _13086_ (.A(_05044_),
    .B(_03045_),
    .C(_00845_),
    .Y(_06171_));
 AO21x1_ASAP7_75t_R _13087_ (.A1(_00844_),
    .A2(_03290_),
    .B(_06171_),
    .Y(_06172_));
 AO221x1_ASAP7_75t_R _13088_ (.A1(_05041_),
    .A2(_06170_),
    .B1(_06172_),
    .B2(_04856_),
    .C(_04411_),
    .Y(_06173_));
 AO22x1_ASAP7_75t_R _13089_ (.A1(_04528_),
    .A2(_00840_),
    .B1(_00841_),
    .B2(_04513_),
    .Y(_06174_));
 AND2x2_ASAP7_75t_R _13090_ (.A(_03155_),
    .B(_00843_),
    .Y(_06175_));
 AO21x1_ASAP7_75t_R _13091_ (.A1(_03056_),
    .A2(_00842_),
    .B(_06175_),
    .Y(_06176_));
 AO221x1_ASAP7_75t_R _13092_ (.A1(_03098_),
    .A2(_00840_),
    .B1(_03925_),
    .B2(_06176_),
    .C(_03914_),
    .Y(_06177_));
 AO21x1_ASAP7_75t_R _13093_ (.A1(_03137_),
    .A2(_06174_),
    .B(_06177_),
    .Y(_06178_));
 AND3x1_ASAP7_75t_R _13094_ (.A(_03703_),
    .B(_06173_),
    .C(_06178_),
    .Y(_06179_));
 AND2x2_ASAP7_75t_R _13095_ (.A(_03092_),
    .B(_00863_),
    .Y(_06180_));
 AO21x1_ASAP7_75t_R _13096_ (.A1(_04080_),
    .A2(_00862_),
    .B(_06180_),
    .Y(_06181_));
 AND3x1_ASAP7_75t_R _13097_ (.A(_05044_),
    .B(_03045_),
    .C(_00861_),
    .Y(_06182_));
 AO21x1_ASAP7_75t_R _13098_ (.A1(_00860_),
    .A2(_03290_),
    .B(_06182_),
    .Y(_06183_));
 AO221x1_ASAP7_75t_R _13099_ (.A1(_05041_),
    .A2(_06181_),
    .B1(_06183_),
    .B2(_04856_),
    .C(_04411_),
    .Y(_06184_));
 AND2x2_ASAP7_75t_R _13100_ (.A(_03087_),
    .B(_00858_),
    .Y(_06185_));
 AO21x2_ASAP7_75t_R _13101_ (.A1(_03161_),
    .A2(_00856_),
    .B(_06185_),
    .Y(_06186_));
 AO21x1_ASAP7_75t_R _13102_ (.A1(_00857_),
    .A2(_04861_),
    .B(_04862_),
    .Y(_06187_));
 AO221x1_ASAP7_75t_R _13103_ (.A1(_00859_),
    .A2(_04413_),
    .B1(_06186_),
    .B2(_05814_),
    .C(_06187_),
    .Y(_06188_));
 AND3x1_ASAP7_75t_R _13104_ (.A(_04043_),
    .B(_06184_),
    .C(_06188_),
    .Y(_06189_));
 OR3x1_ASAP7_75t_R _13105_ (.A(_04545_),
    .B(_06179_),
    .C(_06189_),
    .Y(_06190_));
 AND2x6_ASAP7_75t_R _13106_ (.A(_06168_),
    .B(_06190_),
    .Y(_06191_));
 CKINVDCx20_ASAP7_75t_R _13107_ (.A(_06191_),
    .Y(net128));
 AND3x2_ASAP7_75t_R _13108_ (.A(net89),
    .B(net18),
    .C(_03715_),
    .Y(_09730_));
 NAND2x1_ASAP7_75t_R _13109_ (.A(_03707_),
    .B(_09730_),
    .Y(_06192_));
 OA21x2_ASAP7_75t_R _13110_ (.A1(_03780_),
    .A2(_06191_),
    .B(_06192_),
    .Y(_06193_));
 XNOR2x1_ASAP7_75t_R _13111_ (.B(_06193_),
    .Y(_09681_),
    .A(_03556_));
 INVx1_ASAP7_75t_R _13112_ (.A(_09681_),
    .Y(_09683_));
 INVx3_ASAP7_75t_R _13113_ (.A(_00841_),
    .Y(_06194_));
 NAND2x1_ASAP7_75t_R _13114_ (.A(_00840_),
    .B(_05241_),
    .Y(_06195_));
 OA211x2_ASAP7_75t_R _13115_ (.A1(_06194_),
    .A2(_05557_),
    .B(_04881_),
    .C(_06195_),
    .Y(_06196_));
 OA22x2_ASAP7_75t_R _13116_ (.A1(_00842_),
    .A2(_03429_),
    .B1(_04445_),
    .B2(_00843_),
    .Y(_06197_));
 AND2x2_ASAP7_75t_R _13117_ (.A(_00846_),
    .B(_03466_),
    .Y(_06198_));
 AO221x1_ASAP7_75t_R _13118_ (.A1(_03209_),
    .A2(_04020_),
    .B1(_04023_),
    .B2(_00847_),
    .C(_06198_),
    .Y(_06199_));
 OAI21x1_ASAP7_75t_R _13119_ (.A1(_04885_),
    .A2(_06197_),
    .B(_06199_),
    .Y(_06200_));
 OAI22x1_ASAP7_75t_R _13120_ (.A1(_00845_),
    .A2(_03377_),
    .B1(_04768_),
    .B2(_00844_),
    .Y(_06201_));
 AO221x1_ASAP7_75t_R _13121_ (.A1(_03341_),
    .A2(_06200_),
    .B1(_06201_),
    .B2(_04891_),
    .C(_04552_),
    .Y(_06202_));
 OR2x2_ASAP7_75t_R _13122_ (.A(_06196_),
    .B(_06202_),
    .Y(_06203_));
 NAND2x1_ASAP7_75t_R _13123_ (.A(_00832_),
    .B(_05341_),
    .Y(_06204_));
 NAND2x1_ASAP7_75t_R _13124_ (.A(_00833_),
    .B(_04882_),
    .Y(_06205_));
 OR3x1_ASAP7_75t_R _13125_ (.A(_03097_),
    .B(_04561_),
    .C(_00835_),
    .Y(_06206_));
 OA22x2_ASAP7_75t_R _13126_ (.A1(_00834_),
    .A2(_05106_),
    .B1(_03748_),
    .B2(_06206_),
    .Y(_06207_));
 AND2x2_ASAP7_75t_R _13127_ (.A(_00838_),
    .B(_03847_),
    .Y(_06208_));
 AO221x1_ASAP7_75t_R _13128_ (.A1(_03317_),
    .A2(_03322_),
    .B1(_03429_),
    .B2(_00839_),
    .C(_06208_),
    .Y(_06209_));
 OAI21x1_ASAP7_75t_R _13129_ (.A1(_05127_),
    .A2(_06207_),
    .B(_06209_),
    .Y(_06210_));
 OAI22x1_ASAP7_75t_R _13130_ (.A1(_00836_),
    .A2(_04440_),
    .B1(_05847_),
    .B2(_00837_),
    .Y(_06211_));
 AO221x1_ASAP7_75t_R _13131_ (.A1(_03341_),
    .A2(_06210_),
    .B1(_06211_),
    .B2(_03362_),
    .C(_04899_),
    .Y(_06212_));
 AO32x1_ASAP7_75t_R _13132_ (.A1(_04881_),
    .A2(_06204_),
    .A3(_06205_),
    .B1(_06212_),
    .B2(_03247_),
    .Y(_06213_));
 OA22x2_ASAP7_75t_R _13133_ (.A1(_00850_),
    .A2(_03330_),
    .B1(_03415_),
    .B2(_00851_),
    .Y(_06214_));
 AND2x2_ASAP7_75t_R _13134_ (.A(_00854_),
    .B(_03396_),
    .Y(_06215_));
 AO221x2_ASAP7_75t_R _13135_ (.A1(_03317_),
    .A2(_03322_),
    .B1(_05106_),
    .B2(_00855_),
    .C(_06215_),
    .Y(_06216_));
 OAI21x1_ASAP7_75t_R _13136_ (.A1(_05127_),
    .A2(_06214_),
    .B(_06216_),
    .Y(_06217_));
 AO21x1_ASAP7_75t_R _13137_ (.A1(_05195_),
    .A2(_06217_),
    .B(_04899_),
    .Y(_06218_));
 INVx1_ASAP7_75t_R _13138_ (.A(_00849_),
    .Y(_06219_));
 NAND2x1_ASAP7_75t_R _13139_ (.A(_00848_),
    .B(_05241_),
    .Y(_06220_));
 OA211x2_ASAP7_75t_R _13140_ (.A1(_06219_),
    .A2(_05557_),
    .B(_04881_),
    .C(_06220_),
    .Y(_06221_));
 OAI22x1_ASAP7_75t_R _13141_ (.A1(_00852_),
    .A2(_04440_),
    .B1(_05847_),
    .B2(_00853_),
    .Y(_06222_));
 AND2x2_ASAP7_75t_R _13142_ (.A(_04891_),
    .B(_06222_),
    .Y(_06223_));
 NAND2x1_ASAP7_75t_R _13143_ (.A(_00856_),
    .B(_05847_),
    .Y(_06224_));
 NAND2x1_ASAP7_75t_R _13144_ (.A(_00857_),
    .B(_04768_),
    .Y(_06225_));
 OAI22x1_ASAP7_75t_R _13145_ (.A1(_00861_),
    .A2(_04550_),
    .B1(_04768_),
    .B2(_00860_),
    .Y(_06226_));
 AO32x1_ASAP7_75t_R _13146_ (.A1(_03484_),
    .A2(_06224_),
    .A3(_06225_),
    .B1(_03362_),
    .B2(_06226_),
    .Y(_06227_));
 AND3x1_ASAP7_75t_R _13147_ (.A(_00858_),
    .B(_03317_),
    .C(_03322_),
    .Y(_06228_));
 AOI211x1_ASAP7_75t_R _13148_ (.A1(_00862_),
    .A2(_05127_),
    .B(_04440_),
    .C(_06228_),
    .Y(_06229_));
 INVx2_ASAP7_75t_R _13149_ (.A(_00863_),
    .Y(_06230_));
 AND2x2_ASAP7_75t_R _13150_ (.A(_04020_),
    .B(_04132_),
    .Y(_06231_));
 INVx1_ASAP7_75t_R _13151_ (.A(_00859_),
    .Y(_06232_));
 AO32x1_ASAP7_75t_R _13152_ (.A1(_06230_),
    .A2(_04885_),
    .A3(_05227_),
    .B1(_06231_),
    .B2(_06232_),
    .Y(_06233_));
 OA21x2_ASAP7_75t_R _13153_ (.A1(_06229_),
    .A2(_06233_),
    .B(_05195_),
    .Y(_06234_));
 OA33x2_ASAP7_75t_R _13154_ (.A1(_06218_),
    .A2(_06221_),
    .A3(_06223_),
    .B1(_06227_),
    .B2(_06234_),
    .B3(_03406_),
    .Y(_06235_));
 AO32x2_ASAP7_75t_R _13155_ (.A1(_04484_),
    .A2(_06203_),
    .A3(_06213_),
    .B1(_06235_),
    .B2(_05032_),
    .Y(_06236_));
 INVx1_ASAP7_75t_R _13156_ (.A(_06236_),
    .Y(_09682_));
 AND2x2_ASAP7_75t_R _13157_ (.A(_05044_),
    .B(_00881_),
    .Y(_06237_));
 AO21x1_ASAP7_75t_R _13158_ (.A1(_04095_),
    .A2(_00880_),
    .B(_06237_),
    .Y(_06238_));
 AND3x1_ASAP7_75t_R _13159_ (.A(_05266_),
    .B(_03145_),
    .C(_00879_),
    .Y(_06239_));
 AO21x1_ASAP7_75t_R _13160_ (.A1(_00878_),
    .A2(_05787_),
    .B(_06239_),
    .Y(_06240_));
 AO221x1_ASAP7_75t_R _13161_ (.A1(_05410_),
    .A2(_06238_),
    .B1(_06240_),
    .B2(_05790_),
    .C(_05798_),
    .Y(_06241_));
 AO22x1_ASAP7_75t_R _13162_ (.A1(_03139_),
    .A2(_00874_),
    .B1(_00875_),
    .B2(_04513_),
    .Y(_06242_));
 AND2x2_ASAP7_75t_R _13163_ (.A(_04499_),
    .B(_00877_),
    .Y(_06243_));
 AO21x1_ASAP7_75t_R _13164_ (.A1(_04498_),
    .A2(_00876_),
    .B(_06243_),
    .Y(_06244_));
 AO221x1_ASAP7_75t_R _13165_ (.A1(_03098_),
    .A2(_00874_),
    .B1(_03925_),
    .B2(_06244_),
    .C(_03914_),
    .Y(_06245_));
 AO21x1_ASAP7_75t_R _13166_ (.A1(_03137_),
    .A2(_06242_),
    .B(_06245_),
    .Y(_06246_));
 AND3x1_ASAP7_75t_R _13167_ (.A(_05793_),
    .B(_06241_),
    .C(_06246_),
    .Y(_06247_));
 AND2x2_ASAP7_75t_R _13168_ (.A(_05272_),
    .B(_00873_),
    .Y(_06248_));
 AO21x1_ASAP7_75t_R _13169_ (.A1(_03082_),
    .A2(_00872_),
    .B(_06248_),
    .Y(_06249_));
 AND3x1_ASAP7_75t_R _13170_ (.A(_05266_),
    .B(_03145_),
    .C(_00871_),
    .Y(_06250_));
 AO21x1_ASAP7_75t_R _13171_ (.A1(_00870_),
    .A2(_05787_),
    .B(_06250_),
    .Y(_06251_));
 AO221x1_ASAP7_75t_R _13172_ (.A1(_05410_),
    .A2(_06249_),
    .B1(_06251_),
    .B2(_05790_),
    .C(_05798_),
    .Y(_06252_));
 AO22x1_ASAP7_75t_R _13173_ (.A1(_03139_),
    .A2(_00866_),
    .B1(_00867_),
    .B2(_05370_),
    .Y(_06253_));
 AND2x2_ASAP7_75t_R _13174_ (.A(_03898_),
    .B(_00869_),
    .Y(_06254_));
 AO21x2_ASAP7_75t_R _13175_ (.A1(_04498_),
    .A2(_00868_),
    .B(_06254_),
    .Y(_06255_));
 AO221x1_ASAP7_75t_R _13176_ (.A1(_03098_),
    .A2(_00866_),
    .B1(_03925_),
    .B2(_06255_),
    .C(_03914_),
    .Y(_06256_));
 AO21x1_ASAP7_75t_R _13177_ (.A1(_05372_),
    .A2(_06253_),
    .B(_06256_),
    .Y(_06257_));
 AND3x1_ASAP7_75t_R _13178_ (.A(_05034_),
    .B(_06252_),
    .C(_06257_),
    .Y(_06258_));
 OR2x2_ASAP7_75t_R _13179_ (.A(_04043_),
    .B(_03127_),
    .Y(_06259_));
 AND2x2_ASAP7_75t_R _13180_ (.A(_05266_),
    .B(_00889_),
    .Y(_06260_));
 AO21x1_ASAP7_75t_R _13181_ (.A1(_03082_),
    .A2(_00888_),
    .B(_06260_),
    .Y(_06261_));
 AND3x1_ASAP7_75t_R _13182_ (.A(_05070_),
    .B(_03200_),
    .C(_00887_),
    .Y(_06262_));
 AO21x1_ASAP7_75t_R _13183_ (.A1(_00886_),
    .A2(_05073_),
    .B(_06262_),
    .Y(_06263_));
 AO221x1_ASAP7_75t_R _13184_ (.A1(_05410_),
    .A2(_06261_),
    .B1(_06263_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_06264_));
 AND2x2_ASAP7_75t_R _13185_ (.A(_03674_),
    .B(_00884_),
    .Y(_06265_));
 AO21x1_ASAP7_75t_R _13186_ (.A1(_03161_),
    .A2(_00882_),
    .B(_06265_),
    .Y(_06266_));
 AO21x1_ASAP7_75t_R _13187_ (.A1(_00883_),
    .A2(_04861_),
    .B(_04862_),
    .Y(_06267_));
 AO221x1_ASAP7_75t_R _13188_ (.A1(_00885_),
    .A2(_04413_),
    .B1(_06266_),
    .B2(_05814_),
    .C(_06267_),
    .Y(_06268_));
 AND3x1_ASAP7_75t_R _13189_ (.A(_05034_),
    .B(_06264_),
    .C(_06268_),
    .Y(_06269_));
 AND2x2_ASAP7_75t_R _13190_ (.A(_05266_),
    .B(_00897_),
    .Y(_06270_));
 AO21x1_ASAP7_75t_R _13191_ (.A1(_03082_),
    .A2(_00896_),
    .B(_06270_),
    .Y(_06271_));
 AND3x1_ASAP7_75t_R _13192_ (.A(_05070_),
    .B(_03200_),
    .C(_00895_),
    .Y(_06272_));
 AO21x1_ASAP7_75t_R _13193_ (.A1(_00894_),
    .A2(_05073_),
    .B(_06272_),
    .Y(_06273_));
 AO221x1_ASAP7_75t_R _13194_ (.A1(_05364_),
    .A2(_06271_),
    .B1(_06273_),
    .B2(_05076_),
    .C(_05077_),
    .Y(_06274_));
 AND2x2_ASAP7_75t_R _13195_ (.A(_03674_),
    .B(_00892_),
    .Y(_06275_));
 AO21x1_ASAP7_75t_R _13196_ (.A1(_04381_),
    .A2(_00890_),
    .B(_06275_),
    .Y(_06276_));
 AO21x1_ASAP7_75t_R _13197_ (.A1(_00891_),
    .A2(_04861_),
    .B(_03078_),
    .Y(_06277_));
 AO221x1_ASAP7_75t_R _13198_ (.A1(_00893_),
    .A2(_05061_),
    .B1(_06276_),
    .B2(_05814_),
    .C(_06277_),
    .Y(_06278_));
 AND3x1_ASAP7_75t_R _13199_ (.A(_05793_),
    .B(_06274_),
    .C(_06278_),
    .Y(_06279_));
 OA33x2_ASAP7_75t_R _13200_ (.A1(_06247_),
    .A2(_06258_),
    .A3(_06259_),
    .B1(_06269_),
    .B2(_06279_),
    .B3(_04423_),
    .Y(_06280_));
 CKINVDCx20_ASAP7_75t_R _13201_ (.A(_06280_),
    .Y(net127));
 AND3x2_ASAP7_75t_R _13202_ (.A(net89),
    .B(net17),
    .C(_03715_),
    .Y(_09728_));
 NAND2x1_ASAP7_75t_R _13203_ (.A(_03707_),
    .B(_09728_),
    .Y(_06281_));
 OA21x2_ASAP7_75t_R _13204_ (.A1(_03780_),
    .A2(_06280_),
    .B(_06281_),
    .Y(_06282_));
 XNOR2x1_ASAP7_75t_R _13205_ (.B(_06282_),
    .Y(_09686_),
    .A(_03556_));
 INVx1_ASAP7_75t_R _13206_ (.A(_09686_),
    .Y(_09688_));
 INVx1_ASAP7_75t_R _13207_ (.A(_00875_),
    .Y(_06283_));
 NAND2x1_ASAP7_75t_R _13208_ (.A(_00874_),
    .B(_04473_),
    .Y(_06284_));
 OA211x2_ASAP7_75t_R _13209_ (.A1(_06283_),
    .A2(_04472_),
    .B(_04469_),
    .C(_06284_),
    .Y(_06285_));
 OAI22x1_ASAP7_75t_R _13210_ (.A1(_00879_),
    .A2(_04480_),
    .B1(_03541_),
    .B2(_00878_),
    .Y(_06286_));
 OA22x2_ASAP7_75t_R _13211_ (.A1(_00876_),
    .A2(_03994_),
    .B1(_03765_),
    .B2(_00877_),
    .Y(_06287_));
 AND2x2_ASAP7_75t_R _13212_ (.A(_00880_),
    .B(_03395_),
    .Y(_06288_));
 AO221x1_ASAP7_75t_R _13213_ (.A1(_04574_),
    .A2(_04575_),
    .B1(_03428_),
    .B2(_00881_),
    .C(_06288_),
    .Y(_06289_));
 OAI21x1_ASAP7_75t_R _13214_ (.A1(_03441_),
    .A2(_06287_),
    .B(_06289_),
    .Y(_06290_));
 AO221x1_ASAP7_75t_R _13215_ (.A1(_03540_),
    .A2(_06286_),
    .B1(_06290_),
    .B2(_04026_),
    .C(_03405_),
    .Y(_06291_));
 OAI22x1_ASAP7_75t_R _13216_ (.A1(_00870_),
    .A2(_03330_),
    .B1(_04676_),
    .B2(_00871_),
    .Y(_06292_));
 AND2x2_ASAP7_75t_R _13217_ (.A(_03483_),
    .B(_06292_),
    .Y(_06293_));
 OA22x2_ASAP7_75t_R _13218_ (.A1(_00868_),
    .A2(_03994_),
    .B1(_03418_),
    .B2(_00869_),
    .Y(_06294_));
 AND2x2_ASAP7_75t_R _13219_ (.A(_00872_),
    .B(_03465_),
    .Y(_06295_));
 AO221x1_ASAP7_75t_R _13220_ (.A1(_03316_),
    .A2(_04460_),
    .B1(_04022_),
    .B2(_00873_),
    .C(_06295_),
    .Y(_06296_));
 OA211x2_ASAP7_75t_R _13221_ (.A1(_03441_),
    .A2(_06294_),
    .B(_06296_),
    .C(_03550_),
    .Y(_06297_));
 AND2x2_ASAP7_75t_R _13222_ (.A(_00867_),
    .B(_03454_),
    .Y(_06298_));
 AO21x1_ASAP7_75t_R _13223_ (.A1(_00866_),
    .A2(_03415_),
    .B(_06298_),
    .Y(_06299_));
 OAI22x1_ASAP7_75t_R _13224_ (.A1(_04458_),
    .A2(_06297_),
    .B1(_06299_),
    .B2(_04450_),
    .Y(_06300_));
 OA22x2_ASAP7_75t_R _13225_ (.A1(_06285_),
    .A2(_06291_),
    .B1(_06293_),
    .B2(_06300_),
    .Y(_06301_));
 OA22x2_ASAP7_75t_R _13226_ (.A1(_00892_),
    .A2(_03994_),
    .B1(_03765_),
    .B2(_00893_),
    .Y(_06302_));
 AND2x2_ASAP7_75t_R _13227_ (.A(_00896_),
    .B(_03334_),
    .Y(_06303_));
 AO221x1_ASAP7_75t_R _13228_ (.A1(_03261_),
    .A2(_04018_),
    .B1(_03349_),
    .B2(_00897_),
    .C(_06303_),
    .Y(_06304_));
 OA21x2_ASAP7_75t_R _13229_ (.A1(_03441_),
    .A2(_06302_),
    .B(_06304_),
    .Y(_06305_));
 OA21x2_ASAP7_75t_R _13230_ (.A1(_04786_),
    .A2(_06305_),
    .B(_04791_),
    .Y(_06306_));
 OA22x2_ASAP7_75t_R _13231_ (.A1(_00895_),
    .A2(_04480_),
    .B1(_03541_),
    .B2(_00894_),
    .Y(_06307_));
 AND2x2_ASAP7_75t_R _13232_ (.A(_00891_),
    .B(_03511_),
    .Y(_06308_));
 AO21x1_ASAP7_75t_R _13233_ (.A1(_00890_),
    .A2(_04676_),
    .B(_06308_),
    .Y(_06309_));
 OA22x2_ASAP7_75t_R _13234_ (.A1(_04107_),
    .A2(_06307_),
    .B1(_06309_),
    .B2(_03845_),
    .Y(_06310_));
 OA22x2_ASAP7_75t_R _13235_ (.A1(_00886_),
    .A2(_05106_),
    .B1(_04473_),
    .B2(_00887_),
    .Y(_06311_));
 AND2x2_ASAP7_75t_R _13236_ (.A(_00883_),
    .B(_03454_),
    .Y(_06312_));
 AO21x1_ASAP7_75t_R _13237_ (.A1(_00882_),
    .A2(_04676_),
    .B(_06312_),
    .Y(_06313_));
 OA22x2_ASAP7_75t_R _13238_ (.A1(_04107_),
    .A2(_06311_),
    .B1(_06313_),
    .B2(_04450_),
    .Y(_06314_));
 AO21x1_ASAP7_75t_R _13239_ (.A1(_03045_),
    .A2(_05124_),
    .B(_00888_),
    .Y(_06315_));
 OR3x1_ASAP7_75t_R _13240_ (.A(_00885_),
    .B(_03468_),
    .C(_03356_),
    .Y(_06316_));
 OA211x2_ASAP7_75t_R _13241_ (.A1(_04447_),
    .A2(_06315_),
    .B(_06316_),
    .C(_03299_),
    .Y(_06317_));
 OR4x1_ASAP7_75t_R _13242_ (.A(_00884_),
    .B(_03277_),
    .C(_03468_),
    .D(_03349_),
    .Y(_06318_));
 OA21x2_ASAP7_75t_R _13243_ (.A1(_00889_),
    .A2(_03732_),
    .B(_06318_),
    .Y(_06319_));
 AO21x1_ASAP7_75t_R _13244_ (.A1(_06317_),
    .A2(_06319_),
    .B(_04458_),
    .Y(_06320_));
 AOI221x1_ASAP7_75t_R _13245_ (.A1(_06306_),
    .A2(_06310_),
    .B1(_06314_),
    .B2(_06320_),
    .C(_04003_),
    .Y(_06321_));
 AO21x1_ASAP7_75t_R _13246_ (.A1(_04484_),
    .A2(_06301_),
    .B(_06321_),
    .Y(_06322_));
 BUFx6f_ASAP7_75t_R _13247_ (.A(_06322_),
    .Y(_09685_));
 INVx1_ASAP7_75t_R _13248_ (.A(_09685_),
    .Y(_09687_));
 AND2x2_ASAP7_75t_R _13249_ (.A(_03926_),
    .B(_00902_),
    .Y(_06323_));
 AO21x2_ASAP7_75t_R _13250_ (.A1(_03932_),
    .A2(_00901_),
    .B(_06323_),
    .Y(_06324_));
 AO21x1_ASAP7_75t_R _13251_ (.A1(_03107_),
    .A2(_06324_),
    .B(_04529_),
    .Y(_06325_));
 AO22x1_ASAP7_75t_R _13252_ (.A1(_03111_),
    .A2(_00899_),
    .B1(_00900_),
    .B2(_03626_),
    .Y(_06326_));
 AO22x1_ASAP7_75t_R _13253_ (.A1(_03130_),
    .A2(_00899_),
    .B1(_06326_),
    .B2(_03665_),
    .Y(_06327_));
 AO21x1_ASAP7_75t_R _13254_ (.A1(_03215_),
    .A2(_06325_),
    .B(_06327_),
    .Y(_06328_));
 AND2x2_ASAP7_75t_R _13255_ (.A(_03040_),
    .B(_00906_),
    .Y(_06329_));
 AO21x1_ASAP7_75t_R _13256_ (.A1(_05153_),
    .A2(_00905_),
    .B(_06329_),
    .Y(_06330_));
 AND3x1_ASAP7_75t_R _13257_ (.A(_03065_),
    .B(_04692_),
    .C(_00904_),
    .Y(_06331_));
 AO21x1_ASAP7_75t_R _13258_ (.A1(_00903_),
    .A2(_04376_),
    .B(_06331_),
    .Y(_06332_));
 AO221x1_ASAP7_75t_R _13259_ (.A1(_04487_),
    .A2(_06330_),
    .B1(_06332_),
    .B2(_03582_),
    .C(_04379_),
    .Y(_06333_));
 AND3x1_ASAP7_75t_R _13260_ (.A(_04085_),
    .B(_06328_),
    .C(_06333_),
    .Y(_06334_));
 AND2x2_ASAP7_75t_R _13261_ (.A(_04488_),
    .B(_00914_),
    .Y(_06335_));
 AO21x1_ASAP7_75t_R _13262_ (.A1(_05153_),
    .A2(_00913_),
    .B(_06335_),
    .Y(_06336_));
 AND3x1_ASAP7_75t_R _13263_ (.A(_03065_),
    .B(_04692_),
    .C(_00912_),
    .Y(_06337_));
 AO21x1_ASAP7_75t_R _13264_ (.A1(_00911_),
    .A2(_04376_),
    .B(_06337_),
    .Y(_06338_));
 AO221x1_ASAP7_75t_R _13265_ (.A1(_04722_),
    .A2(_06336_),
    .B1(_06338_),
    .B2(_03582_),
    .C(_04379_),
    .Y(_06339_));
 AO22x1_ASAP7_75t_R _13266_ (.A1(_03685_),
    .A2(_00907_),
    .B1(_00908_),
    .B2(_04361_),
    .Y(_06340_));
 AND2x2_ASAP7_75t_R _13267_ (.A(_03091_),
    .B(_00910_),
    .Y(_06341_));
 AO21x1_ASAP7_75t_R _13268_ (.A1(_03932_),
    .A2(_00909_),
    .B(_06341_),
    .Y(_06342_));
 AO21x1_ASAP7_75t_R _13269_ (.A1(_03107_),
    .A2(_06342_),
    .B(_04529_),
    .Y(_06343_));
 AO21x1_ASAP7_75t_R _13270_ (.A1(_04381_),
    .A2(_06340_),
    .B(_06343_),
    .Y(_06344_));
 AND3x2_ASAP7_75t_R _13271_ (.A(_03119_),
    .B(_06339_),
    .C(_06344_),
    .Y(_06345_));
 OR3x1_ASAP7_75t_R _13272_ (.A(_04043_),
    .B(_06334_),
    .C(_06345_),
    .Y(_06346_));
 AND2x2_ASAP7_75t_R _13273_ (.A(_03065_),
    .B(_00930_),
    .Y(_06347_));
 AO21x1_ASAP7_75t_R _13274_ (.A1(_03138_),
    .A2(_00929_),
    .B(_06347_),
    .Y(_06348_));
 AND3x1_ASAP7_75t_R _13275_ (.A(_04087_),
    .B(_04009_),
    .C(_00928_),
    .Y(_06349_));
 AO21x1_ASAP7_75t_R _13276_ (.A1(_00927_),
    .A2(_04376_),
    .B(_06349_),
    .Y(_06350_));
 AO221x1_ASAP7_75t_R _13277_ (.A1(_04068_),
    .A2(_06348_),
    .B1(_06350_),
    .B2(_04074_),
    .C(_04379_),
    .Y(_06351_));
 AND2x2_ASAP7_75t_R _13278_ (.A(_03088_),
    .B(_00925_),
    .Y(_06352_));
 AO21x1_ASAP7_75t_R _13279_ (.A1(_03160_),
    .A2(_00923_),
    .B(_06352_),
    .Y(_06353_));
 AO21x1_ASAP7_75t_R _13280_ (.A1(_00924_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_06354_));
 AO221x1_ASAP7_75t_R _13281_ (.A1(_00926_),
    .A2(_04077_),
    .B1(_06353_),
    .B2(_04080_),
    .C(_06354_),
    .Y(_06355_));
 AND3x1_ASAP7_75t_R _13282_ (.A(_04098_),
    .B(_06351_),
    .C(_06355_),
    .Y(_06356_));
 AND2x2_ASAP7_75t_R _13283_ (.A(_03065_),
    .B(_00922_),
    .Y(_06357_));
 AO21x1_ASAP7_75t_R _13284_ (.A1(_03138_),
    .A2(_00921_),
    .B(_06357_),
    .Y(_06358_));
 AND3x1_ASAP7_75t_R _13285_ (.A(_04087_),
    .B(_04692_),
    .C(_00920_),
    .Y(_06359_));
 AO21x1_ASAP7_75t_R _13286_ (.A1(_00919_),
    .A2(_04376_),
    .B(_06359_),
    .Y(_06360_));
 AO221x1_ASAP7_75t_R _13287_ (.A1(_04068_),
    .A2(_06358_),
    .B1(_06360_),
    .B2(_04074_),
    .C(_04379_),
    .Y(_06361_));
 AND2x2_ASAP7_75t_R _13288_ (.A(_03647_),
    .B(_00917_),
    .Y(_06362_));
 AO21x1_ASAP7_75t_R _13289_ (.A1(_03160_),
    .A2(_00915_),
    .B(_06362_),
    .Y(_06363_));
 AO21x1_ASAP7_75t_R _13290_ (.A1(_00916_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_06364_));
 AO221x2_ASAP7_75t_R _13291_ (.A1(_00918_),
    .A2(_03697_),
    .B1(_06363_),
    .B2(_04080_),
    .C(_06364_),
    .Y(_06365_));
 AND3x1_ASAP7_75t_R _13292_ (.A(_04085_),
    .B(_06361_),
    .C(_06365_),
    .Y(_06366_));
 OR3x1_ASAP7_75t_R _13293_ (.A(_04100_),
    .B(_06356_),
    .C(_06366_),
    .Y(_06367_));
 AOI21x1_ASAP7_75t_R _13294_ (.A1(_06346_),
    .A2(_06367_),
    .B(_03781_),
    .Y(net3));
 AND3x1_ASAP7_75t_R _13295_ (.A(net89),
    .B(net16),
    .C(_03715_),
    .Y(_09726_));
 AND2x2_ASAP7_75t_R _13296_ (.A(_03707_),
    .B(_09726_),
    .Y(_06368_));
 AOI21x1_ASAP7_75t_R _13297_ (.A1(_04159_),
    .A2(net126),
    .B(_06368_),
    .Y(_06369_));
 XNOR2x1_ASAP7_75t_R _13298_ (.B(_06369_),
    .Y(_09691_),
    .A(_03556_));
 INVx1_ASAP7_75t_R _13299_ (.A(_09691_),
    .Y(_09693_));
 OA22x2_ASAP7_75t_R _13300_ (.A1(_00903_),
    .A2(_03348_),
    .B1(_03355_),
    .B2(_00904_),
    .Y(_06370_));
 AND2x2_ASAP7_75t_R _13301_ (.A(_00899_),
    .B(_03355_),
    .Y(_06371_));
 AND2x2_ASAP7_75t_R _13302_ (.A(_00900_),
    .B(_03453_),
    .Y(_06372_));
 OA33x2_ASAP7_75t_R _13303_ (.A1(_03343_),
    .A2(_03865_),
    .A3(_06370_),
    .B1(_06371_),
    .B2(_06372_),
    .B3(_03844_),
    .Y(_06373_));
 AND3x1_ASAP7_75t_R _13304_ (.A(_03043_),
    .B(_03474_),
    .C(_00906_),
    .Y(_06374_));
 AOI221x1_ASAP7_75t_R _13305_ (.A1(_03324_),
    .A2(_03506_),
    .B1(_03395_),
    .B2(_00905_),
    .C(_06374_),
    .Y(_06375_));
 INVx1_ASAP7_75t_R _13306_ (.A(_00902_),
    .Y(_06376_));
 OA211x2_ASAP7_75t_R _13307_ (.A1(_03197_),
    .A2(_03309_),
    .B(_03303_),
    .C(_06376_),
    .Y(_06377_));
 NOR2x1_ASAP7_75t_R _13308_ (.A(_00901_),
    .B(_03312_),
    .Y(_06378_));
 OA211x2_ASAP7_75t_R _13309_ (.A1(_06377_),
    .A2(_06378_),
    .B(_03260_),
    .C(_03320_),
    .Y(_06379_));
 OAI21x1_ASAP7_75t_R _13310_ (.A1(_06375_),
    .A2(_06379_),
    .B(_03501_),
    .Y(_06380_));
 AO21x1_ASAP7_75t_R _13311_ (.A1(_03298_),
    .A2(_06380_),
    .B(_03344_),
    .Y(_06381_));
 AND2x2_ASAP7_75t_R _13312_ (.A(_00908_),
    .B(_03399_),
    .Y(_06382_));
 AO21x1_ASAP7_75t_R _13313_ (.A1(_00907_),
    .A2(_03413_),
    .B(_06382_),
    .Y(_06383_));
 OA21x2_ASAP7_75t_R _13314_ (.A1(_00909_),
    .A2(_03303_),
    .B(_03319_),
    .Y(_06384_));
 OA21x2_ASAP7_75t_R _13315_ (.A1(_00910_),
    .A2(_03354_),
    .B(_06384_),
    .Y(_06385_));
 OA21x2_ASAP7_75t_R _13316_ (.A1(_03338_),
    .A2(_06385_),
    .B(_03324_),
    .Y(_06386_));
 AND3x1_ASAP7_75t_R _13317_ (.A(_03018_),
    .B(_03301_),
    .C(_00914_),
    .Y(_06387_));
 AO21x1_ASAP7_75t_R _13318_ (.A1(_00913_),
    .A2(_03333_),
    .B(_06387_),
    .Y(_06388_));
 AND2x2_ASAP7_75t_R _13319_ (.A(_03503_),
    .B(_06388_),
    .Y(_06389_));
 OA22x2_ASAP7_75t_R _13320_ (.A1(_00912_),
    .A2(_03465_),
    .B1(_03399_),
    .B2(_00911_),
    .Y(_06390_));
 OA222x2_ASAP7_75t_R _13321_ (.A1(_03844_),
    .A2(_06383_),
    .B1(_06386_),
    .B2(_06389_),
    .C1(_06390_),
    .C2(_03865_),
    .Y(_06391_));
 AOI221x1_ASAP7_75t_R _13322_ (.A1(_06373_),
    .A2(_06381_),
    .B1(_06391_),
    .B2(_03888_),
    .C(_03425_),
    .Y(_06392_));
 INVx1_ASAP7_75t_R _13323_ (.A(_00916_),
    .Y(_06393_));
 NAND2x1_ASAP7_75t_R _13324_ (.A(_00915_),
    .B(_03449_),
    .Y(_06394_));
 OA211x2_ASAP7_75t_R _13325_ (.A1(_06393_),
    .A2(_04153_),
    .B(_03446_),
    .C(_06394_),
    .Y(_06395_));
 OAI22x1_ASAP7_75t_R _13326_ (.A1(_00919_),
    .A2(_03304_),
    .B1(_03430_),
    .B2(_00920_),
    .Y(_06396_));
 AND2x2_ASAP7_75t_R _13327_ (.A(_03360_),
    .B(_06396_),
    .Y(_06397_));
 AND3x1_ASAP7_75t_R _13328_ (.A(_03116_),
    .B(_03474_),
    .C(_00922_),
    .Y(_06398_));
 AOI221x1_ASAP7_75t_R _13329_ (.A1(_03207_),
    .A2(_03386_),
    .B1(_03435_),
    .B2(_00921_),
    .C(_06398_),
    .Y(_06399_));
 INVx1_ASAP7_75t_R _13330_ (.A(_00918_),
    .Y(_06400_));
 OA211x2_ASAP7_75t_R _13331_ (.A1(net24),
    .A2(_03309_),
    .B(_03302_),
    .C(_06400_),
    .Y(_06401_));
 NOR2x1_ASAP7_75t_R _13332_ (.A(_00917_),
    .B(_03303_),
    .Y(_06402_));
 OA211x2_ASAP7_75t_R _13333_ (.A1(_06401_),
    .A2(_06402_),
    .B(_03206_),
    .C(_03319_),
    .Y(_06403_));
 OA21x2_ASAP7_75t_R _13334_ (.A1(_06399_),
    .A2(_06403_),
    .B(_03339_),
    .Y(_06404_));
 OA31x2_ASAP7_75t_R _13335_ (.A1(_03460_),
    .A2(_06397_),
    .A3(_06404_),
    .B1(_03244_),
    .Y(_06405_));
 OA21x2_ASAP7_75t_R _13336_ (.A1(_00925_),
    .A2(_03303_),
    .B(_03319_),
    .Y(_06406_));
 OAI21x1_ASAP7_75t_R _13337_ (.A1(_00926_),
    .A2(_03430_),
    .B(_06406_),
    .Y(_06407_));
 AO21x1_ASAP7_75t_R _13338_ (.A1(_03381_),
    .A2(_06407_),
    .B(_03276_),
    .Y(_06408_));
 AND3x1_ASAP7_75t_R _13339_ (.A(_03018_),
    .B(_03301_),
    .C(_00930_),
    .Y(_06409_));
 AO21x1_ASAP7_75t_R _13340_ (.A1(_00929_),
    .A2(_03435_),
    .B(_06409_),
    .Y(_06410_));
 NAND2x1_ASAP7_75t_R _13341_ (.A(_03503_),
    .B(_06410_),
    .Y(_06411_));
 OAI22x1_ASAP7_75t_R _13342_ (.A1(_00928_),
    .A2(_03395_),
    .B1(_03453_),
    .B2(_00927_),
    .Y(_06412_));
 OA211x2_ASAP7_75t_R _13343_ (.A1(_03197_),
    .A2(_03309_),
    .B(_03303_),
    .C(_00924_),
    .Y(_06413_));
 AOI21x1_ASAP7_75t_R _13344_ (.A1(_00923_),
    .A2(_03430_),
    .B(_06413_),
    .Y(_06414_));
 AO21x1_ASAP7_75t_R _13345_ (.A1(_03420_),
    .A2(_06414_),
    .B(_03298_),
    .Y(_06415_));
 AO221x1_ASAP7_75t_R _13346_ (.A1(_06408_),
    .A2(_06411_),
    .B1(_06412_),
    .B2(_03482_),
    .C(_06415_),
    .Y(_06416_));
 OA211x2_ASAP7_75t_R _13347_ (.A1(_06395_),
    .A2(_06405_),
    .B(_06416_),
    .C(_03424_),
    .Y(_06417_));
 OR2x2_ASAP7_75t_R _13348_ (.A(_06392_),
    .B(_06417_),
    .Y(_06418_));
 BUFx3_ASAP7_75t_R _13349_ (.A(_06418_),
    .Y(_09690_));
 INVx2_ASAP7_75t_R _13350_ (.A(_09690_),
    .Y(_09692_));
 AOI21x1_ASAP7_75t_R _13351_ (.A1(_03210_),
    .A2(_03227_),
    .B(_03249_),
    .Y(_06419_));
 AO21x2_ASAP7_75t_R _13352_ (.A1(_03708_),
    .A2(_03275_),
    .B(_04979_),
    .Y(_06420_));
 AO22x2_ASAP7_75t_R _13353_ (.A1(net5),
    .A2(_06419_),
    .B1(_06420_),
    .B2(_03033_),
    .Y(_06421_));
 AND2x2_ASAP7_75t_R _13354_ (.A(net89),
    .B(_06421_),
    .Y(_09724_));
 AND2x2_ASAP7_75t_R _13355_ (.A(_03692_),
    .B(_00956_),
    .Y(_06422_));
 AO21x1_ASAP7_75t_R _13356_ (.A1(_03565_),
    .A2(_00955_),
    .B(_06422_),
    .Y(_06423_));
 AND3x1_ASAP7_75t_R _13357_ (.A(_03926_),
    .B(_03860_),
    .C(_00954_),
    .Y(_06424_));
 AO21x1_ASAP7_75t_R _13358_ (.A1(_00953_),
    .A2(_03289_),
    .B(_06424_),
    .Y(_06425_));
 AO221x2_ASAP7_75t_R _13359_ (.A1(_03689_),
    .A2(_06423_),
    .B1(_06425_),
    .B2(_03681_),
    .C(_03695_),
    .Y(_06426_));
 AO22x1_ASAP7_75t_R _13360_ (.A1(_03945_),
    .A2(_00949_),
    .B1(_00950_),
    .B2(_03946_),
    .Y(_06427_));
 AND2x2_ASAP7_75t_R _13361_ (.A(_03807_),
    .B(_00952_),
    .Y(_06428_));
 AO21x1_ASAP7_75t_R _13362_ (.A1(_03061_),
    .A2(_00951_),
    .B(_06428_),
    .Y(_06429_));
 AO221x1_ASAP7_75t_R _13363_ (.A1(_03597_),
    .A2(_00949_),
    .B1(_03909_),
    .B2(_06429_),
    .C(_03936_),
    .Y(_06430_));
 AO21x1_ASAP7_75t_R _13364_ (.A1(_03068_),
    .A2(_06427_),
    .B(_06430_),
    .Y(_06431_));
 AO21x1_ASAP7_75t_R _13365_ (.A1(_06426_),
    .A2(_06431_),
    .B(_03154_),
    .Y(_06432_));
 AND2x2_ASAP7_75t_R _13366_ (.A(_03692_),
    .B(_00940_),
    .Y(_06433_));
 AO21x1_ASAP7_75t_R _13367_ (.A1(_03565_),
    .A2(_00939_),
    .B(_06433_),
    .Y(_06434_));
 AND3x1_ASAP7_75t_R _13368_ (.A(_03926_),
    .B(_03860_),
    .C(_00938_),
    .Y(_06435_));
 AO21x1_ASAP7_75t_R _13369_ (.A1(_00937_),
    .A2(_03289_),
    .B(_06435_),
    .Y(_06436_));
 AO221x2_ASAP7_75t_R _13370_ (.A1(_03689_),
    .A2(_06434_),
    .B1(_06436_),
    .B2(_03681_),
    .C(_03695_),
    .Y(_06437_));
 AO22x1_ASAP7_75t_R _13371_ (.A1(_03620_),
    .A2(_00933_),
    .B1(_00934_),
    .B2(_03946_),
    .Y(_06438_));
 AND2x2_ASAP7_75t_R _13372_ (.A(_03807_),
    .B(_00936_),
    .Y(_06439_));
 AO21x1_ASAP7_75t_R _13373_ (.A1(_03061_),
    .A2(_00935_),
    .B(_06439_),
    .Y(_06440_));
 AO221x1_ASAP7_75t_R _13374_ (.A1(_03597_),
    .A2(_00933_),
    .B1(_03909_),
    .B2(_06440_),
    .C(_03936_),
    .Y(_06441_));
 AO21x1_ASAP7_75t_R _13375_ (.A1(_03068_),
    .A2(_06438_),
    .B(_06441_),
    .Y(_06442_));
 AO21x1_ASAP7_75t_R _13376_ (.A1(_06437_),
    .A2(_06442_),
    .B(_03142_),
    .Y(_06443_));
 AO21x1_ASAP7_75t_R _13377_ (.A1(_06432_),
    .A2(_06443_),
    .B(_03127_),
    .Y(_06444_));
 AO22x1_ASAP7_75t_R _13378_ (.A1(_03062_),
    .A2(_00957_),
    .B1(_00958_),
    .B2(_04361_),
    .Y(_06445_));
 AND2x2_ASAP7_75t_R _13379_ (.A(_03039_),
    .B(_00960_),
    .Y(_06446_));
 AO21x1_ASAP7_75t_R _13380_ (.A1(_03055_),
    .A2(_00959_),
    .B(_06446_),
    .Y(_06447_));
 AO221x1_ASAP7_75t_R _13381_ (.A1(_03597_),
    .A2(_00957_),
    .B1(_03909_),
    .B2(_06447_),
    .C(_03936_),
    .Y(_06448_));
 AO21x1_ASAP7_75t_R _13382_ (.A1(_03161_),
    .A2(_06445_),
    .B(_06448_),
    .Y(_06449_));
 AND2x2_ASAP7_75t_R _13383_ (.A(_03091_),
    .B(_00964_),
    .Y(_06450_));
 AO21x1_ASAP7_75t_R _13384_ (.A1(_03932_),
    .A2(_00963_),
    .B(_06450_),
    .Y(_06451_));
 AND3x1_ASAP7_75t_R _13385_ (.A(_03578_),
    .B(_03063_),
    .C(_00962_),
    .Y(_06452_));
 AO21x1_ASAP7_75t_R _13386_ (.A1(_00961_),
    .A2(_03577_),
    .B(_06452_),
    .Y(_06453_));
 AO221x1_ASAP7_75t_R _13387_ (.A1(_03571_),
    .A2(_06451_),
    .B1(_06453_),
    .B2(_03604_),
    .C(_03583_),
    .Y(_06454_));
 AO21x1_ASAP7_75t_R _13388_ (.A1(_06449_),
    .A2(_06454_),
    .B(_03154_),
    .Y(_06455_));
 AO22x1_ASAP7_75t_R _13389_ (.A1(_03062_),
    .A2(_00941_),
    .B1(_00942_),
    .B2(_04361_),
    .Y(_06456_));
 AND2x2_ASAP7_75t_R _13390_ (.A(_03039_),
    .B(_00944_),
    .Y(_06457_));
 AO21x2_ASAP7_75t_R _13391_ (.A1(_03080_),
    .A2(_00943_),
    .B(_06457_),
    .Y(_06458_));
 AO221x1_ASAP7_75t_R _13392_ (.A1(_03597_),
    .A2(_00941_),
    .B1(_03909_),
    .B2(_06458_),
    .C(_03936_),
    .Y(_06459_));
 AO21x1_ASAP7_75t_R _13393_ (.A1(_03161_),
    .A2(_06456_),
    .B(_06459_),
    .Y(_06460_));
 AND2x2_ASAP7_75t_R _13394_ (.A(_03091_),
    .B(_00948_),
    .Y(_06461_));
 AO21x1_ASAP7_75t_R _13395_ (.A1(_03932_),
    .A2(_00947_),
    .B(_06461_),
    .Y(_06462_));
 AND3x1_ASAP7_75t_R _13396_ (.A(_03578_),
    .B(_03063_),
    .C(_00946_),
    .Y(_06463_));
 AO21x1_ASAP7_75t_R _13397_ (.A1(_00945_),
    .A2(_03577_),
    .B(_06463_),
    .Y(_06464_));
 AO221x2_ASAP7_75t_R _13398_ (.A1(_03571_),
    .A2(_06462_),
    .B1(_06464_),
    .B2(_03604_),
    .C(_03583_),
    .Y(_06465_));
 AO21x1_ASAP7_75t_R _13399_ (.A1(_06460_),
    .A2(_06465_),
    .B(_03142_),
    .Y(_06466_));
 AO21x2_ASAP7_75t_R _13400_ (.A1(_06455_),
    .A2(_06466_),
    .B(_04404_),
    .Y(_06467_));
 OAI21x1_ASAP7_75t_R _13401_ (.A1(_06444_),
    .A2(_05793_),
    .B(_06467_),
    .Y(net125));
 AND3x1_ASAP7_75t_R _13402_ (.A(_03024_),
    .B(_03270_),
    .C(_06421_),
    .Y(_06468_));
 AOI21x1_ASAP7_75t_R _13403_ (.A1(_03558_),
    .A2(net125),
    .B(_06468_),
    .Y(_06469_));
 BUFx4f_ASAP7_75t_R _13404_ (.A(_06469_),
    .Y(_06470_));
 BUFx4f_ASAP7_75t_R _13405_ (.A(_06470_),
    .Y(_06471_));
 BUFx6f_ASAP7_75t_R _13406_ (.A(_06471_),
    .Y(_06472_));
 XNOR2x1_ASAP7_75t_R _13407_ (.B(_06472_),
    .Y(_09696_),
    .A(_03556_));
 INVx1_ASAP7_75t_R _13408_ (.A(_09696_),
    .Y(_09698_));
 OR3x1_ASAP7_75t_R _13409_ (.A(_03597_),
    .B(_04561_),
    .C(_00936_),
    .Y(_06473_));
 OA22x2_ASAP7_75t_R _13410_ (.A1(_00935_),
    .A2(_04023_),
    .B1(_03748_),
    .B2(_06473_),
    .Y(_06474_));
 AND3x1_ASAP7_75t_R _13411_ (.A(_04503_),
    .B(_03475_),
    .C(_00940_),
    .Y(_06475_));
 AO221x1_ASAP7_75t_R _13412_ (.A1(_03251_),
    .A2(_03388_),
    .B1(_03335_),
    .B2(_00939_),
    .C(_06475_),
    .Y(_06476_));
 OAI21x1_ASAP7_75t_R _13413_ (.A1(_04885_),
    .A2(_06474_),
    .B(_06476_),
    .Y(_06477_));
 INVx1_ASAP7_75t_R _13414_ (.A(_00933_),
    .Y(_01248_));
 INVx1_ASAP7_75t_R _13415_ (.A(_00934_),
    .Y(_06478_));
 AND2x2_ASAP7_75t_R _13416_ (.A(_06478_),
    .B(_04132_),
    .Y(_06479_));
 AO21x1_ASAP7_75t_R _13417_ (.A1(_01248_),
    .A2(_04451_),
    .B(_06479_),
    .Y(_06480_));
 OR3x1_ASAP7_75t_R _13418_ (.A(_03096_),
    .B(_03749_),
    .C(_00938_),
    .Y(_06481_));
 AO21x1_ASAP7_75t_R _13419_ (.A1(_03351_),
    .A2(_03352_),
    .B(_06481_),
    .Y(_06482_));
 AO21x1_ASAP7_75t_R _13420_ (.A1(_03149_),
    .A2(_05124_),
    .B(_00937_),
    .Y(_06483_));
 AO21x2_ASAP7_75t_R _13421_ (.A1(_06482_),
    .A2(_06483_),
    .B(_03979_),
    .Y(_06484_));
 AOI22x1_ASAP7_75t_R _13422_ (.A1(_04784_),
    .A2(_04783_),
    .B1(_04771_),
    .B2(_06484_),
    .Y(_06485_));
 AOI221x1_ASAP7_75t_R _13423_ (.A1(_03444_),
    .A2(_06477_),
    .B1(_06480_),
    .B2(_03448_),
    .C(_06485_),
    .Y(_06486_));
 AND2x2_ASAP7_75t_R _13424_ (.A(_00942_),
    .B(_03511_),
    .Y(_06487_));
 AO21x2_ASAP7_75t_R _13425_ (.A1(_00941_),
    .A2(_03357_),
    .B(_06487_),
    .Y(_06488_));
 OAI22x1_ASAP7_75t_R _13426_ (.A1(_00946_),
    .A2(_03976_),
    .B1(_04466_),
    .B2(_00945_),
    .Y(_06489_));
 AOI221x1_ASAP7_75t_R _13427_ (.A1(_04784_),
    .A2(_04783_),
    .B1(_03457_),
    .B2(_06489_),
    .C(_03299_),
    .Y(_06490_));
 INVx1_ASAP7_75t_R _13428_ (.A(_00944_),
    .Y(_06491_));
 OA211x2_ASAP7_75t_R _13429_ (.A1(_03488_),
    .A2(_03490_),
    .B(_03522_),
    .C(_06491_),
    .Y(_06492_));
 OAI21x1_ASAP7_75t_R _13430_ (.A1(_00943_),
    .A2(_03428_),
    .B(_04018_),
    .Y(_06493_));
 OA21x2_ASAP7_75t_R _13431_ (.A1(_06492_),
    .A2(_06493_),
    .B(_03382_),
    .Y(_06494_));
 AND3x1_ASAP7_75t_R _13432_ (.A(_03034_),
    .B(_03475_),
    .C(_00948_),
    .Y(_06495_));
 AOI21x1_ASAP7_75t_R _13433_ (.A1(_00947_),
    .A2(_03976_),
    .B(_06495_),
    .Y(_06496_));
 OAI22x1_ASAP7_75t_R _13434_ (.A1(_03278_),
    .A2(_06494_),
    .B1(_06496_),
    .B2(_03394_),
    .Y(_06497_));
 OA211x2_ASAP7_75t_R _13435_ (.A1(_03845_),
    .A2(_06488_),
    .B(_06490_),
    .C(_06497_),
    .Y(_06498_));
 OR3x4_ASAP7_75t_R _13436_ (.A(_03426_),
    .B(_06486_),
    .C(_06498_),
    .Y(_06499_));
 INVx1_ASAP7_75t_R _13437_ (.A(_00952_),
    .Y(_06500_));
 OA211x2_ASAP7_75t_R _13438_ (.A1(_03488_),
    .A2(_03311_),
    .B(_03313_),
    .C(_06500_),
    .Y(_06501_));
 NOR2x1_ASAP7_75t_R _13439_ (.A(_00951_),
    .B(_03385_),
    .Y(_06502_));
 OA211x2_ASAP7_75t_R _13440_ (.A1(_06501_),
    .A2(_06502_),
    .B(_03209_),
    .C(_04020_),
    .Y(_06503_));
 AND2x2_ASAP7_75t_R _13441_ (.A(_00955_),
    .B(_03396_),
    .Y(_06504_));
 AOI221x1_ASAP7_75t_R _13442_ (.A1(_03317_),
    .A2(_03322_),
    .B1(_03330_),
    .B2(_00956_),
    .C(_06504_),
    .Y(_06505_));
 OA21x2_ASAP7_75t_R _13443_ (.A1(_06503_),
    .A2(_06505_),
    .B(_03341_),
    .Y(_06506_));
 OA21x2_ASAP7_75t_R _13444_ (.A1(_04899_),
    .A2(_06506_),
    .B(_03412_),
    .Y(_06507_));
 OA211x2_ASAP7_75t_R _13445_ (.A1(_03226_),
    .A2(_03311_),
    .B(_04022_),
    .C(_00950_),
    .Y(_06508_));
 AOI21x1_ASAP7_75t_R _13446_ (.A1(_00949_),
    .A2(_04473_),
    .B(_06508_),
    .Y(_06509_));
 AND2x2_ASAP7_75t_R _13447_ (.A(_04786_),
    .B(_06509_),
    .Y(_06510_));
 OAI22x1_ASAP7_75t_R _13448_ (.A1(_00953_),
    .A2(_05106_),
    .B1(_04473_),
    .B2(_00954_),
    .Y(_06511_));
 AND3x1_ASAP7_75t_R _13449_ (.A(_04786_),
    .B(_05314_),
    .C(_06511_),
    .Y(_06512_));
 AND3x1_ASAP7_75t_R _13450_ (.A(_04784_),
    .B(_04783_),
    .C(_06509_),
    .Y(_06513_));
 AO221x2_ASAP7_75t_R _13451_ (.A1(_05842_),
    .A2(_06510_),
    .B1(_06512_),
    .B2(_03412_),
    .C(_06513_),
    .Y(_06514_));
 INVx1_ASAP7_75t_R _13452_ (.A(_00960_),
    .Y(_06515_));
 OA211x2_ASAP7_75t_R _13453_ (.A1(_03226_),
    .A2(_03311_),
    .B(_03313_),
    .C(_06515_),
    .Y(_06516_));
 OAI21x1_ASAP7_75t_R _13454_ (.A1(_00959_),
    .A2(_03306_),
    .B(_03388_),
    .Y(_06517_));
 OA21x2_ASAP7_75t_R _13455_ (.A1(_06516_),
    .A2(_06517_),
    .B(_03382_),
    .Y(_06518_));
 AND3x1_ASAP7_75t_R _13456_ (.A(_03045_),
    .B(_05124_),
    .C(_00964_),
    .Y(_06519_));
 AOI21x1_ASAP7_75t_R _13457_ (.A1(_00963_),
    .A2(_03378_),
    .B(_06519_),
    .Y(_06520_));
 OA22x2_ASAP7_75t_R _13458_ (.A1(_03278_),
    .A2(_06518_),
    .B1(_06520_),
    .B2(_05318_),
    .Y(_06521_));
 OA211x2_ASAP7_75t_R _13459_ (.A1(_03226_),
    .A2(_03311_),
    .B(_03428_),
    .C(_00958_),
    .Y(_06522_));
 AOI21x1_ASAP7_75t_R _13460_ (.A1(_00957_),
    .A2(_03357_),
    .B(_06522_),
    .Y(_06523_));
 AO221x1_ASAP7_75t_R _13461_ (.A1(_04784_),
    .A2(_04783_),
    .B1(_03484_),
    .B2(_06523_),
    .C(_04771_),
    .Y(_06524_));
 OAI22x1_ASAP7_75t_R _13462_ (.A1(_00962_),
    .A2(_03397_),
    .B1(_03541_),
    .B2(_00961_),
    .Y(_06525_));
 OA211x2_ASAP7_75t_R _13463_ (.A1(_03284_),
    .A2(_03288_),
    .B(_03362_),
    .C(_06525_),
    .Y(_06526_));
 OA31x2_ASAP7_75t_R _13464_ (.A1(_06521_),
    .A2(_06524_),
    .A3(_06526_),
    .B1(_03495_),
    .Y(_06527_));
 OAI21x1_ASAP7_75t_R _13465_ (.A1(_06507_),
    .A2(_06514_),
    .B(_06527_),
    .Y(_06528_));
 NAND2x1_ASAP7_75t_R _13466_ (.A(_06499_),
    .B(_06528_),
    .Y(_09695_));
 INVx1_ASAP7_75t_R _13467_ (.A(_09695_),
    .Y(_09697_));
 AO32x1_ASAP7_75t_R _13468_ (.A1(_03023_),
    .A2(net2),
    .A3(_06419_),
    .B1(_06420_),
    .B2(_03175_),
    .Y(_06529_));
 BUFx3_ASAP7_75t_R _13469_ (.A(_06529_),
    .Y(_09722_));
 AND2x2_ASAP7_75t_R _13470_ (.A(_05366_),
    .B(_00997_),
    .Y(_06530_));
 AO21x1_ASAP7_75t_R _13471_ (.A1(_05064_),
    .A2(_00996_),
    .B(_06530_),
    .Y(_06531_));
 AND3x1_ASAP7_75t_R _13472_ (.A(_05366_),
    .B(_03201_),
    .C(_00995_),
    .Y(_06532_));
 AO21x1_ASAP7_75t_R _13473_ (.A1(_00994_),
    .A2(_03291_),
    .B(_06532_),
    .Y(_06533_));
 AO221x1_ASAP7_75t_R _13474_ (.A1(_05365_),
    .A2(_06531_),
    .B1(_06533_),
    .B2(_04764_),
    .C(_05260_),
    .Y(_06534_));
 AND2x2_ASAP7_75t_R _13475_ (.A(_05366_),
    .B(_00989_),
    .Y(_06535_));
 AO21x1_ASAP7_75t_R _13476_ (.A1(_05064_),
    .A2(_00988_),
    .B(_06535_),
    .Y(_06536_));
 AND3x1_ASAP7_75t_R _13477_ (.A(_05366_),
    .B(_03215_),
    .C(_00987_),
    .Y(_06537_));
 AO21x1_ASAP7_75t_R _13478_ (.A1(_00986_),
    .A2(_03291_),
    .B(_06537_),
    .Y(_06538_));
 AO221x1_ASAP7_75t_R _13479_ (.A1(_05365_),
    .A2(_06536_),
    .B1(_06538_),
    .B2(_04764_),
    .C(_05253_),
    .Y(_06539_));
 AND3x1_ASAP7_75t_R _13480_ (.A(_04486_),
    .B(_06534_),
    .C(_06539_),
    .Y(_06540_));
 AND2x2_ASAP7_75t_R _13481_ (.A(_04389_),
    .B(_00984_),
    .Y(_06541_));
 AO21x1_ASAP7_75t_R _13482_ (.A1(_03137_),
    .A2(_00982_),
    .B(_06541_),
    .Y(_06542_));
 AO221x1_ASAP7_75t_R _13483_ (.A1(_05041_),
    .A2(_00985_),
    .B1(_05269_),
    .B2(_00983_),
    .C(_05814_),
    .Y(_06543_));
 OA211x2_ASAP7_75t_R _13484_ (.A1(_05376_),
    .A2(_06542_),
    .B(_06543_),
    .C(_05034_),
    .Y(_06544_));
 AND2x2_ASAP7_75t_R _13485_ (.A(_04389_),
    .B(_00992_),
    .Y(_06545_));
 AO21x1_ASAP7_75t_R _13486_ (.A1(_03137_),
    .A2(_00990_),
    .B(_06545_),
    .Y(_06546_));
 AO221x1_ASAP7_75t_R _13487_ (.A1(_05041_),
    .A2(_00993_),
    .B1(_05269_),
    .B2(_00991_),
    .C(_05814_),
    .Y(_06547_));
 OA211x2_ASAP7_75t_R _13488_ (.A1(_05376_),
    .A2(_06546_),
    .B(_06547_),
    .C(_03174_),
    .Y(_06548_));
 OR3x1_ASAP7_75t_R _13489_ (.A(_05067_),
    .B(_06544_),
    .C(_06548_),
    .Y(_06549_));
 AND2x2_ASAP7_75t_R _13490_ (.A(_04389_),
    .B(_00976_),
    .Y(_06550_));
 AO21x1_ASAP7_75t_R _13491_ (.A1(_03137_),
    .A2(_00974_),
    .B(_06550_),
    .Y(_06551_));
 AO21x1_ASAP7_75t_R _13492_ (.A1(_00977_),
    .A2(_05061_),
    .B(_05067_),
    .Y(_06552_));
 AO221x1_ASAP7_75t_R _13493_ (.A1(_00975_),
    .A2(_05066_),
    .B1(_06551_),
    .B2(_05375_),
    .C(_06552_),
    .Y(_06553_));
 AND2x2_ASAP7_75t_R _13494_ (.A(_03049_),
    .B(_00981_),
    .Y(_06554_));
 AO21x1_ASAP7_75t_R _13495_ (.A1(_05064_),
    .A2(_00980_),
    .B(_06554_),
    .Y(_06555_));
 AND3x1_ASAP7_75t_R _13496_ (.A(_05366_),
    .B(_03215_),
    .C(_00979_),
    .Y(_06556_));
 AO21x1_ASAP7_75t_R _13497_ (.A1(_00978_),
    .A2(_03291_),
    .B(_06556_),
    .Y(_06557_));
 AO221x1_ASAP7_75t_R _13498_ (.A1(_05365_),
    .A2(_06555_),
    .B1(_06557_),
    .B2(_04764_),
    .C(_04657_),
    .Y(_06558_));
 AO22x1_ASAP7_75t_R _13499_ (.A1(_05814_),
    .A2(_00966_),
    .B1(_00967_),
    .B2(_05370_),
    .Y(_06559_));
 AND2x2_ASAP7_75t_R _13500_ (.A(_03041_),
    .B(_00969_),
    .Y(_06560_));
 AO21x1_ASAP7_75t_R _13501_ (.A1(_03139_),
    .A2(_00968_),
    .B(_06560_),
    .Y(_06561_));
 AO21x1_ASAP7_75t_R _13502_ (.A1(_05069_),
    .A2(_06561_),
    .B(_05474_),
    .Y(_06562_));
 AND2x2_ASAP7_75t_R _13503_ (.A(_03099_),
    .B(_00966_),
    .Y(_06563_));
 AO221x1_ASAP7_75t_R _13504_ (.A1(_05372_),
    .A2(_06559_),
    .B1(_06562_),
    .B2(_03023_),
    .C(_06563_),
    .Y(_06564_));
 AND2x2_ASAP7_75t_R _13505_ (.A(_03071_),
    .B(_00973_),
    .Y(_06565_));
 AO21x1_ASAP7_75t_R _13506_ (.A1(_04860_),
    .A2(_00972_),
    .B(_06565_),
    .Y(_06566_));
 AO21x1_ASAP7_75t_R _13507_ (.A1(_05069_),
    .A2(_06566_),
    .B(_04657_),
    .Y(_06567_));
 AND3x1_ASAP7_75t_R _13508_ (.A(_05366_),
    .B(_03201_),
    .C(_00971_),
    .Y(_06568_));
 OA21x2_ASAP7_75t_R _13509_ (.A1(_04401_),
    .A2(_03131_),
    .B(_00970_),
    .Y(_06569_));
 OA21x2_ASAP7_75t_R _13510_ (.A1(_06568_),
    .A2(_06569_),
    .B(_05076_),
    .Y(_06570_));
 OA21x2_ASAP7_75t_R _13511_ (.A1(_06567_),
    .A2(_06570_),
    .B(_04545_),
    .Y(_06571_));
 AO32x1_ASAP7_75t_R _13512_ (.A1(_03175_),
    .A2(_06553_),
    .A3(_06558_),
    .B1(_06564_),
    .B2(_06571_),
    .Y(_06572_));
 AO221x2_ASAP7_75t_R _13513_ (.A1(_06540_),
    .A2(_06549_),
    .B1(_06572_),
    .B2(_04423_),
    .C(_04163_),
    .Y(_06573_));
 CKINVDCx20_ASAP7_75t_R _13514_ (.A(_06573_),
    .Y(net124));
 NAND2x1_ASAP7_75t_R _13515_ (.A(_03558_),
    .B(_06573_),
    .Y(_06574_));
 OA21x2_ASAP7_75t_R _13516_ (.A1(_03558_),
    .A2(_09722_),
    .B(_06574_),
    .Y(_06575_));
 BUFx4f_ASAP7_75t_R _13517_ (.A(_06575_),
    .Y(_06576_));
 BUFx4f_ASAP7_75t_R _13518_ (.A(_06576_),
    .Y(_06577_));
 BUFx4f_ASAP7_75t_R _13519_ (.A(_06577_),
    .Y(_06578_));
 XNOR2x1_ASAP7_75t_R _13520_ (.B(_06578_),
    .Y(_09701_),
    .A(_03259_));
 INVx1_ASAP7_75t_R _13521_ (.A(_09701_),
    .Y(_09703_));
 OR3x1_ASAP7_75t_R _13522_ (.A(_03130_),
    .B(_04561_),
    .C(_00985_),
    .Y(_06579_));
 OA22x2_ASAP7_75t_R _13523_ (.A1(_00984_),
    .A2(_04896_),
    .B1(_03748_),
    .B2(_06579_),
    .Y(_06580_));
 AND3x1_ASAP7_75t_R _13524_ (.A(_03200_),
    .B(_05335_),
    .C(_00989_),
    .Y(_06581_));
 AO221x1_ASAP7_75t_R _13525_ (.A1(_03326_),
    .A2(_05842_),
    .B1(_03378_),
    .B2(_00988_),
    .C(_06581_),
    .Y(_06582_));
 OA21x2_ASAP7_75t_R _13526_ (.A1(_05093_),
    .A2(_06580_),
    .B(_06582_),
    .Y(_06583_));
 AO21x1_ASAP7_75t_R _13527_ (.A1(_03300_),
    .A2(_06583_),
    .B(_04458_),
    .Y(_06584_));
 OA22x2_ASAP7_75t_R _13528_ (.A1(_00986_),
    .A2(_04440_),
    .B1(_05847_),
    .B2(_00987_),
    .Y(_06585_));
 AND2x2_ASAP7_75t_R _13529_ (.A(_00982_),
    .B(_05847_),
    .Y(_06586_));
 AND2x2_ASAP7_75t_R _13530_ (.A(_00983_),
    .B(_03410_),
    .Y(_06587_));
 OA33x2_ASAP7_75t_R _13531_ (.A1(_03345_),
    .A2(_03979_),
    .A3(_06585_),
    .B1(_06586_),
    .B2(_06587_),
    .B3(_04450_),
    .Y(_06588_));
 AND2x2_ASAP7_75t_R _13532_ (.A(_00990_),
    .B(_05557_),
    .Y(_06589_));
 AO221x1_ASAP7_75t_R _13533_ (.A1(_00991_),
    .A2(_04882_),
    .B1(_03411_),
    .B2(_03247_),
    .C(_06589_),
    .Y(_06590_));
 OAI22x1_ASAP7_75t_R _13534_ (.A1(_00995_),
    .A2(_04550_),
    .B1(_04882_),
    .B2(_00994_),
    .Y(_06591_));
 OA22x2_ASAP7_75t_R _13535_ (.A1(_00992_),
    .A2(_04440_),
    .B1(_05847_),
    .B2(_00993_),
    .Y(_06592_));
 AND2x2_ASAP7_75t_R _13536_ (.A(_00996_),
    .B(_04480_),
    .Y(_06593_));
 AO221x1_ASAP7_75t_R _13537_ (.A1(_03210_),
    .A2(_05842_),
    .B1(_05227_),
    .B2(_00997_),
    .C(_06593_),
    .Y(_06594_));
 OAI21x1_ASAP7_75t_R _13538_ (.A1(_05093_),
    .A2(_06592_),
    .B(_06594_),
    .Y(_06595_));
 AOI221x1_ASAP7_75t_R _13539_ (.A1(_04549_),
    .A2(_06591_),
    .B1(_06595_),
    .B2(_05195_),
    .C(_03406_),
    .Y(_06596_));
 AOI22x1_ASAP7_75t_R _13540_ (.A1(_06584_),
    .A2(_06588_),
    .B1(_06590_),
    .B2(_06596_),
    .Y(_06597_));
 AND2x2_ASAP7_75t_R _13541_ (.A(_00974_),
    .B(_05557_),
    .Y(_06598_));
 AO221x1_ASAP7_75t_R _13542_ (.A1(_00975_),
    .A2(_04882_),
    .B1(_03411_),
    .B2(_03247_),
    .C(_06598_),
    .Y(_06599_));
 OAI22x1_ASAP7_75t_R _13543_ (.A1(_00979_),
    .A2(_04550_),
    .B1(_04882_),
    .B2(_00978_),
    .Y(_06600_));
 OA22x2_ASAP7_75t_R _13544_ (.A1(_00976_),
    .A2(_04440_),
    .B1(_05241_),
    .B2(_00977_),
    .Y(_06601_));
 AND2x2_ASAP7_75t_R _13545_ (.A(_00980_),
    .B(_04480_),
    .Y(_06602_));
 AO221x1_ASAP7_75t_R _13546_ (.A1(_03326_),
    .A2(_05842_),
    .B1(_05227_),
    .B2(_00981_),
    .C(_06602_),
    .Y(_06603_));
 OAI21x1_ASAP7_75t_R _13547_ (.A1(_05093_),
    .A2(_06601_),
    .B(_06603_),
    .Y(_06604_));
 AOI221x1_ASAP7_75t_R _13548_ (.A1(_04549_),
    .A2(_06600_),
    .B1(_06604_),
    .B2(_05195_),
    .C(_03406_),
    .Y(_06605_));
 OR3x1_ASAP7_75t_R _13549_ (.A(_03098_),
    .B(_04561_),
    .C(_00973_),
    .Y(_06606_));
 OR4x1_ASAP7_75t_R _13550_ (.A(_00969_),
    .B(_03470_),
    .C(_05314_),
    .D(_03432_),
    .Y(_06607_));
 OA211x2_ASAP7_75t_R _13551_ (.A1(_05318_),
    .A2(_06606_),
    .B(_06607_),
    .C(_04771_),
    .Y(_06608_));
 AND3x1_ASAP7_75t_R _13552_ (.A(_00968_),
    .B(_03326_),
    .C(_05842_),
    .Y(_06609_));
 AO221x1_ASAP7_75t_R _13553_ (.A1(_03022_),
    .A2(_05335_),
    .B1(_00972_),
    .B2(_05127_),
    .C(_06609_),
    .Y(_06610_));
 AO21x1_ASAP7_75t_R _13554_ (.A1(_06608_),
    .A2(_06610_),
    .B(_04458_),
    .Y(_06611_));
 OA22x2_ASAP7_75t_R _13555_ (.A1(_00970_),
    .A2(_04440_),
    .B1(_05241_),
    .B2(_00971_),
    .Y(_06612_));
 AND2x2_ASAP7_75t_R _13556_ (.A(_00966_),
    .B(_05847_),
    .Y(_06613_));
 AND2x2_ASAP7_75t_R _13557_ (.A(_00967_),
    .B(_04768_),
    .Y(_06614_));
 OA33x2_ASAP7_75t_R _13558_ (.A1(_03345_),
    .A2(_03979_),
    .A3(_06612_),
    .B1(_06613_),
    .B2(_06614_),
    .B3(_04450_),
    .Y(_06615_));
 AOI22x1_ASAP7_75t_R _13559_ (.A1(_06599_),
    .A2(_06605_),
    .B1(_06611_),
    .B2(_06615_),
    .Y(_06616_));
 AO32x1_ASAP7_75t_R _13560_ (.A1(_03247_),
    .A2(_03539_),
    .A3(_06597_),
    .B1(_06616_),
    .B2(_04484_),
    .Y(_06617_));
 BUFx4f_ASAP7_75t_R _13561_ (.A(_06617_),
    .Y(_09700_));
 INVx2_ASAP7_75t_R _13562_ (.A(_09700_),
    .Y(_09702_));
 AO21x2_ASAP7_75t_R _13563_ (.A1(_03023_),
    .A2(net30),
    .B(_03238_),
    .Y(_06618_));
 AO32x1_ASAP7_75t_R _13564_ (.A1(_05067_),
    .A2(_03023_),
    .A3(_06420_),
    .B1(_06618_),
    .B2(_06419_),
    .Y(_06619_));
 BUFx2_ASAP7_75t_R _13565_ (.A(_06619_),
    .Y(_09716_));
 AND2x2_ASAP7_75t_R _13566_ (.A(_05272_),
    .B(_01014_),
    .Y(_06620_));
 AO21x1_ASAP7_75t_R _13567_ (.A1(_03082_),
    .A2(_01013_),
    .B(_06620_),
    .Y(_06621_));
 AO21x1_ASAP7_75t_R _13568_ (.A1(_05364_),
    .A2(_06621_),
    .B(_04411_),
    .Y(_06622_));
 AND3x1_ASAP7_75t_R _13569_ (.A(_03049_),
    .B(_05229_),
    .C(_01012_),
    .Y(_06623_));
 OA21x2_ASAP7_75t_R _13570_ (.A1(_04748_),
    .A2(_04493_),
    .B(_01011_),
    .Y(_06624_));
 OA21x2_ASAP7_75t_R _13571_ (.A1(_06623_),
    .A2(_06624_),
    .B(_04856_),
    .Y(_06625_));
 AND2x2_ASAP7_75t_R _13572_ (.A(_03593_),
    .B(_01009_),
    .Y(_06626_));
 AO21x1_ASAP7_75t_R _13573_ (.A1(_03132_),
    .A2(_01007_),
    .B(_06626_),
    .Y(_06627_));
 AO21x1_ASAP7_75t_R _13574_ (.A1(_01010_),
    .A2(_03697_),
    .B(_04862_),
    .Y(_06628_));
 AO221x1_ASAP7_75t_R _13575_ (.A1(_01008_),
    .A2(_05066_),
    .B1(_06627_),
    .B2(_04860_),
    .C(_06628_),
    .Y(_06629_));
 OA21x2_ASAP7_75t_R _13576_ (.A1(_06622_),
    .A2(_06625_),
    .B(_06629_),
    .Y(_06630_));
 AO22x1_ASAP7_75t_R _13577_ (.A1(_04401_),
    .A2(_00999_),
    .B1(_01000_),
    .B2(_05370_),
    .Y(_06631_));
 AND2x2_ASAP7_75t_R _13578_ (.A(_04408_),
    .B(_01002_),
    .Y(_06632_));
 AO21x1_ASAP7_75t_R _13579_ (.A1(_04748_),
    .A2(_01001_),
    .B(_06632_),
    .Y(_06633_));
 AO21x1_ASAP7_75t_R _13580_ (.A1(_04850_),
    .A2(_06633_),
    .B(_05474_),
    .Y(_06634_));
 AND2x2_ASAP7_75t_R _13581_ (.A(_03131_),
    .B(_00999_),
    .Y(_06635_));
 AO221x1_ASAP7_75t_R _13582_ (.A1(_05372_),
    .A2(_06631_),
    .B1(_06634_),
    .B2(_03216_),
    .C(_06635_),
    .Y(_06636_));
 AND2x2_ASAP7_75t_R _13583_ (.A(_05070_),
    .B(_01006_),
    .Y(_06637_));
 AO21x1_ASAP7_75t_R _13584_ (.A1(_04528_),
    .A2(_01005_),
    .B(_06637_),
    .Y(_06638_));
 AO21x1_ASAP7_75t_R _13585_ (.A1(_05364_),
    .A2(_06638_),
    .B(_05798_),
    .Y(_06639_));
 AND3x1_ASAP7_75t_R _13586_ (.A(_03049_),
    .B(_05229_),
    .C(_01004_),
    .Y(_06640_));
 OA21x2_ASAP7_75t_R _13587_ (.A1(_04080_),
    .A2(_03098_),
    .B(_01003_),
    .Y(_06641_));
 OA21x2_ASAP7_75t_R _13588_ (.A1(_06640_),
    .A2(_06641_),
    .B(_05790_),
    .Y(_06642_));
 OA21x2_ASAP7_75t_R _13589_ (.A1(_06639_),
    .A2(_06642_),
    .B(_05034_),
    .Y(_06643_));
 AO221x1_ASAP7_75t_R _13590_ (.A1(_05793_),
    .A2(_06630_),
    .B1(_06636_),
    .B2(_06643_),
    .C(_04486_),
    .Y(_06644_));
 AND2x2_ASAP7_75t_R _13591_ (.A(_05272_),
    .B(_01030_),
    .Y(_06645_));
 AO21x1_ASAP7_75t_R _13592_ (.A1(_04095_),
    .A2(_01029_),
    .B(_06645_),
    .Y(_06646_));
 AO21x1_ASAP7_75t_R _13593_ (.A1(_05364_),
    .A2(_06646_),
    .B(_04411_),
    .Y(_06647_));
 AND3x1_ASAP7_75t_R _13594_ (.A(_03049_),
    .B(_05229_),
    .C(_01028_),
    .Y(_06648_));
 OA21x2_ASAP7_75t_R _13595_ (.A1(_04851_),
    .A2(_04493_),
    .B(_01027_),
    .Y(_06649_));
 OA21x2_ASAP7_75t_R _13596_ (.A1(_06648_),
    .A2(_06649_),
    .B(_04856_),
    .Y(_06650_));
 AND2x2_ASAP7_75t_R _13597_ (.A(_03593_),
    .B(_01025_),
    .Y(_06651_));
 AO21x1_ASAP7_75t_R _13598_ (.A1(_03132_),
    .A2(_01023_),
    .B(_06651_),
    .Y(_06652_));
 AO21x1_ASAP7_75t_R _13599_ (.A1(_01026_),
    .A2(_03697_),
    .B(_04416_),
    .Y(_06653_));
 AO221x1_ASAP7_75t_R _13600_ (.A1(_01024_),
    .A2(_04861_),
    .B1(_06652_),
    .B2(_04860_),
    .C(_06653_),
    .Y(_06654_));
 OA21x2_ASAP7_75t_R _13601_ (.A1(_06647_),
    .A2(_06650_),
    .B(_06654_),
    .Y(_06655_));
 AO22x1_ASAP7_75t_R _13602_ (.A1(_04401_),
    .A2(_01015_),
    .B1(_01016_),
    .B2(_05370_),
    .Y(_06656_));
 AND2x2_ASAP7_75t_R _13603_ (.A(_04408_),
    .B(_01018_),
    .Y(_06657_));
 AO21x1_ASAP7_75t_R _13604_ (.A1(_04748_),
    .A2(_01017_),
    .B(_06657_),
    .Y(_06658_));
 AO21x1_ASAP7_75t_R _13605_ (.A1(_04850_),
    .A2(_06658_),
    .B(_03078_),
    .Y(_06659_));
 AND2x2_ASAP7_75t_R _13606_ (.A(_03131_),
    .B(_01015_),
    .Y(_06660_));
 AO221x1_ASAP7_75t_R _13607_ (.A1(_05372_),
    .A2(_06656_),
    .B1(_06659_),
    .B2(_03216_),
    .C(_06660_),
    .Y(_06661_));
 AND2x2_ASAP7_75t_R _13608_ (.A(_05266_),
    .B(_01022_),
    .Y(_06662_));
 AO21x1_ASAP7_75t_R _13609_ (.A1(_04528_),
    .A2(_01021_),
    .B(_06662_),
    .Y(_06663_));
 AO21x1_ASAP7_75t_R _13610_ (.A1(_05364_),
    .A2(_06663_),
    .B(_05798_),
    .Y(_06664_));
 AND3x1_ASAP7_75t_R _13611_ (.A(_03049_),
    .B(_05229_),
    .C(_01020_),
    .Y(_06665_));
 OA21x2_ASAP7_75t_R _13612_ (.A1(_04748_),
    .A2(_03098_),
    .B(_01019_),
    .Y(_06666_));
 OA21x2_ASAP7_75t_R _13613_ (.A1(_06665_),
    .A2(_06666_),
    .B(_05790_),
    .Y(_06667_));
 OA21x2_ASAP7_75t_R _13614_ (.A1(_06664_),
    .A2(_06667_),
    .B(_04404_),
    .Y(_06668_));
 AO221x1_ASAP7_75t_R _13615_ (.A1(_05793_),
    .A2(_06655_),
    .B1(_06661_),
    .B2(_06668_),
    .C(_04423_),
    .Y(_06669_));
 AO21x2_ASAP7_75t_R _13616_ (.A1(_06644_),
    .A2(_06669_),
    .B(_04163_),
    .Y(_06670_));
 CKINVDCx20_ASAP7_75t_R _13617_ (.A(_06670_),
    .Y(net121));
 NAND2x1_ASAP7_75t_R _13618_ (.A(_03283_),
    .B(_06670_),
    .Y(_06671_));
 OA21x2_ASAP7_75t_R _13619_ (.A1(_03558_),
    .A2(_09716_),
    .B(_06671_),
    .Y(_06672_));
 BUFx4f_ASAP7_75t_R _13620_ (.A(_06672_),
    .Y(_06673_));
 BUFx4f_ASAP7_75t_R _13621_ (.A(_06673_),
    .Y(_06674_));
 BUFx6f_ASAP7_75t_R _13622_ (.A(_06674_),
    .Y(_06675_));
 XNOR2x1_ASAP7_75t_R _13623_ (.B(_06675_),
    .Y(_09706_),
    .A(_03259_));
 INVx1_ASAP7_75t_R _13624_ (.A(_09706_),
    .Y(_09708_));
 OAI22x1_ASAP7_75t_R _13625_ (.A1(_01019_),
    .A2(_05248_),
    .B1(_05341_),
    .B2(_01020_),
    .Y(_06676_));
 OR2x2_ASAP7_75t_R _13626_ (.A(_01015_),
    .B(_03410_),
    .Y(_06677_));
 OAI21x1_ASAP7_75t_R _13627_ (.A1(_01016_),
    .A2(_05341_),
    .B(_06677_),
    .Y(_06678_));
 OA222x2_ASAP7_75t_R _13628_ (.A1(_03099_),
    .A2(_03965_),
    .B1(_01022_),
    .B2(_03732_),
    .C1(_03733_),
    .C2(_01018_),
    .Y(_06679_));
 AND3x1_ASAP7_75t_R _13629_ (.A(_01017_),
    .B(_03326_),
    .C(_05842_),
    .Y(_06680_));
 AO221x1_ASAP7_75t_R _13630_ (.A1(_03216_),
    .A2(_05335_),
    .B1(_01021_),
    .B2(_05093_),
    .C(_06680_),
    .Y(_06681_));
 AOI21x1_ASAP7_75t_R _13631_ (.A1(_06679_),
    .A2(_06681_),
    .B(_04458_),
    .Y(_06682_));
 AO221x1_ASAP7_75t_R _13632_ (.A1(_04549_),
    .A2(_06676_),
    .B1(_06678_),
    .B2(_04881_),
    .C(_06682_),
    .Y(_06683_));
 OAI22x1_ASAP7_75t_R _13633_ (.A1(_01028_),
    .A2(_04550_),
    .B1(_04882_),
    .B2(_01027_),
    .Y(_06684_));
 OR2x2_ASAP7_75t_R _13634_ (.A(_01023_),
    .B(_03455_),
    .Y(_06685_));
 OAI21x1_ASAP7_75t_R _13635_ (.A1(_01024_),
    .A2(_05341_),
    .B(_06685_),
    .Y(_06686_));
 OA22x2_ASAP7_75t_R _13636_ (.A1(_01025_),
    .A2(_05227_),
    .B1(_05241_),
    .B2(_01026_),
    .Y(_06687_));
 AND2x2_ASAP7_75t_R _13637_ (.A(_01029_),
    .B(_03976_),
    .Y(_06688_));
 AO221x1_ASAP7_75t_R _13638_ (.A1(_03326_),
    .A2(_05842_),
    .B1(_04896_),
    .B2(_01030_),
    .C(_06688_),
    .Y(_06689_));
 OAI21x1_ASAP7_75t_R _13639_ (.A1(_05093_),
    .A2(_06687_),
    .B(_06689_),
    .Y(_06690_));
 AO221x1_ASAP7_75t_R _13640_ (.A1(_04881_),
    .A2(_06686_),
    .B1(_06690_),
    .B2(_05195_),
    .C(_03406_),
    .Y(_06691_));
 AO21x1_ASAP7_75t_R _13641_ (.A1(_04549_),
    .A2(_06684_),
    .B(_06691_),
    .Y(_06692_));
 INVx1_ASAP7_75t_R _13642_ (.A(_01008_),
    .Y(_06693_));
 NAND2x1_ASAP7_75t_R _13643_ (.A(_01007_),
    .B(_05341_),
    .Y(_06694_));
 OA211x2_ASAP7_75t_R _13644_ (.A1(_06693_),
    .A2(_05341_),
    .B(_04881_),
    .C(_06694_),
    .Y(_06695_));
 OAI22x1_ASAP7_75t_R _13645_ (.A1(_01012_),
    .A2(_04550_),
    .B1(_03410_),
    .B2(_01011_),
    .Y(_06696_));
 OA22x2_ASAP7_75t_R _13646_ (.A1(_01009_),
    .A2(_04896_),
    .B1(_04472_),
    .B2(_01010_),
    .Y(_06697_));
 AND2x2_ASAP7_75t_R _13647_ (.A(_01013_),
    .B(_03335_),
    .Y(_06698_));
 AO221x1_ASAP7_75t_R _13648_ (.A1(_03326_),
    .A2(_05842_),
    .B1(_04896_),
    .B2(_01014_),
    .C(_06698_),
    .Y(_06699_));
 OAI21x1_ASAP7_75t_R _13649_ (.A1(_05093_),
    .A2(_06697_),
    .B(_06699_),
    .Y(_06700_));
 AO221x1_ASAP7_75t_R _13650_ (.A1(_04549_),
    .A2(_06696_),
    .B1(_06700_),
    .B2(_05195_),
    .C(_03406_),
    .Y(_06701_));
 OR3x1_ASAP7_75t_R _13651_ (.A(_03131_),
    .B(_04561_),
    .C(_01006_),
    .Y(_06702_));
 OR4x1_ASAP7_75t_R _13652_ (.A(_01002_),
    .B(_03470_),
    .C(_05314_),
    .D(_03383_),
    .Y(_06703_));
 OA211x2_ASAP7_75t_R _13653_ (.A1(_05318_),
    .A2(_06702_),
    .B(_06703_),
    .C(_03300_),
    .Y(_06704_));
 AND3x1_ASAP7_75t_R _13654_ (.A(_01001_),
    .B(_03210_),
    .C(_05842_),
    .Y(_06705_));
 AO221x1_ASAP7_75t_R _13655_ (.A1(_03216_),
    .A2(_05335_),
    .B1(_01005_),
    .B2(_05093_),
    .C(_06705_),
    .Y(_06706_));
 AOI21x1_ASAP7_75t_R _13656_ (.A1(_06704_),
    .A2(_06706_),
    .B(_04458_),
    .Y(_06707_));
 NAND2x1_ASAP7_75t_R _13657_ (.A(_00999_),
    .B(_05341_),
    .Y(_06708_));
 NAND2x1_ASAP7_75t_R _13658_ (.A(_01000_),
    .B(_04882_),
    .Y(_06709_));
 OAI22x1_ASAP7_75t_R _13659_ (.A1(_01003_),
    .A2(_05248_),
    .B1(_05341_),
    .B2(_01004_),
    .Y(_06710_));
 AO32x1_ASAP7_75t_R _13660_ (.A1(_04881_),
    .A2(_06708_),
    .A3(_06709_),
    .B1(_04549_),
    .B2(_06710_),
    .Y(_06711_));
 OA22x2_ASAP7_75t_R _13661_ (.A1(_06695_),
    .A2(_06701_),
    .B1(_06707_),
    .B2(_06711_),
    .Y(_06712_));
 BUFx4f_ASAP7_75t_R _13662_ (.A(_04484_),
    .Y(_06713_));
 AO32x2_ASAP7_75t_R _13663_ (.A1(_05032_),
    .A2(_06683_),
    .A3(_06692_),
    .B1(_06712_),
    .B2(_06713_),
    .Y(_06714_));
 BUFx6f_ASAP7_75t_R _13664_ (.A(_06714_),
    .Y(_09705_));
 INVx1_ASAP7_75t_R _13665_ (.A(_09705_),
    .Y(_09707_));
 AO21x2_ASAP7_75t_R _13666_ (.A1(_03022_),
    .A2(net29),
    .B(_03238_),
    .Y(_06715_));
 AO32x2_ASAP7_75t_R _13667_ (.A1(_05365_),
    .A2(net89),
    .A3(_06420_),
    .B1(_06715_),
    .B2(_06419_),
    .Y(_09553_));
 AO22x1_ASAP7_75t_R _13668_ (.A1(_03945_),
    .A2(_01032_),
    .B1(_01033_),
    .B2(_03946_),
    .Y(_06716_));
 AND2x2_ASAP7_75t_R _13669_ (.A(_03675_),
    .B(_01035_),
    .Y(_06717_));
 AO21x1_ASAP7_75t_R _13670_ (.A1(_03111_),
    .A2(_01034_),
    .B(_06717_),
    .Y(_06718_));
 AO21x1_ASAP7_75t_R _13671_ (.A1(_03087_),
    .A2(_06718_),
    .B(_03077_),
    .Y(_06719_));
 AND2x2_ASAP7_75t_R _13672_ (.A(_03097_),
    .B(_01032_),
    .Y(_06720_));
 AO221x1_ASAP7_75t_R _13673_ (.A1(_03068_),
    .A2(_06716_),
    .B1(_06719_),
    .B2(_03215_),
    .C(_06720_),
    .Y(_06721_));
 AND2x2_ASAP7_75t_R _13674_ (.A(_03692_),
    .B(_01039_),
    .Y(_06722_));
 AO21x1_ASAP7_75t_R _13675_ (.A1(_03565_),
    .A2(_01038_),
    .B(_06722_),
    .Y(_06723_));
 AO21x1_ASAP7_75t_R _13676_ (.A1(_03689_),
    .A2(_06723_),
    .B(_03695_),
    .Y(_06724_));
 AND3x1_ASAP7_75t_R _13677_ (.A(_03155_),
    .B(_03020_),
    .C(_01037_),
    .Y(_06725_));
 OA21x2_ASAP7_75t_R _13678_ (.A1(_03630_),
    .A2(_04492_),
    .B(_01036_),
    .Y(_06726_));
 OA21x2_ASAP7_75t_R _13679_ (.A1(_06725_),
    .A2(_06726_),
    .B(_03681_),
    .Y(_06727_));
 OA21x2_ASAP7_75t_R _13680_ (.A1(_06724_),
    .A2(_06727_),
    .B(_03586_),
    .Y(_06728_));
 AND2x2_ASAP7_75t_R _13681_ (.A(_03678_),
    .B(_01047_),
    .Y(_06729_));
 AO21x1_ASAP7_75t_R _13682_ (.A1(_03565_),
    .A2(_01046_),
    .B(_06729_),
    .Y(_06730_));
 AO21x1_ASAP7_75t_R _13683_ (.A1(_03689_),
    .A2(_06730_),
    .B(_03636_),
    .Y(_06731_));
 AND3x1_ASAP7_75t_R _13684_ (.A(_03058_),
    .B(_04009_),
    .C(_01045_),
    .Y(_06732_));
 OA21x2_ASAP7_75t_R _13685_ (.A1(_03630_),
    .A2(_04492_),
    .B(_01044_),
    .Y(_06733_));
 OA21x2_ASAP7_75t_R _13686_ (.A1(_06732_),
    .A2(_06733_),
    .B(_03681_),
    .Y(_06734_));
 AND2x2_ASAP7_75t_R _13687_ (.A(_03085_),
    .B(_01042_),
    .Y(_06735_));
 AO21x1_ASAP7_75t_R _13688_ (.A1(_03588_),
    .A2(_01040_),
    .B(_06735_),
    .Y(_06736_));
 AO21x1_ASAP7_75t_R _13689_ (.A1(_01043_),
    .A2(_03567_),
    .B(_03650_),
    .Y(_06737_));
 AO221x1_ASAP7_75t_R _13690_ (.A1(_01041_),
    .A2(_03560_),
    .B1(_06736_),
    .B2(_03620_),
    .C(_06737_),
    .Y(_06738_));
 OA211x2_ASAP7_75t_R _13691_ (.A1(_06731_),
    .A2(_06734_),
    .B(_03173_),
    .C(_06738_),
    .Y(_06739_));
 AOI211x1_ASAP7_75t_R _13692_ (.A1(_06721_),
    .A2(_06728_),
    .B(_06739_),
    .C(_03143_),
    .Y(_06740_));
 AND2x2_ASAP7_75t_R _13693_ (.A(_03692_),
    .B(_01063_),
    .Y(_06741_));
 AO21x1_ASAP7_75t_R _13694_ (.A1(_03910_),
    .A2(_01062_),
    .B(_06741_),
    .Y(_06742_));
 AO21x1_ASAP7_75t_R _13695_ (.A1(_03689_),
    .A2(_06742_),
    .B(_03695_),
    .Y(_06743_));
 AND3x1_ASAP7_75t_R _13696_ (.A(_03894_),
    .B(_03020_),
    .C(_01061_),
    .Y(_06744_));
 OA21x2_ASAP7_75t_R _13697_ (.A1(_03111_),
    .A2(_04492_),
    .B(_01060_),
    .Y(_06745_));
 OA21x2_ASAP7_75t_R _13698_ (.A1(_06744_),
    .A2(_06745_),
    .B(_03681_),
    .Y(_06746_));
 AND2x2_ASAP7_75t_R _13699_ (.A(_03072_),
    .B(_01058_),
    .Y(_06747_));
 AO21x1_ASAP7_75t_R _13700_ (.A1(_03027_),
    .A2(_01056_),
    .B(_06747_),
    .Y(_06748_));
 AO22x1_ASAP7_75t_R _13701_ (.A1(_01059_),
    .A2(_03568_),
    .B1(_06748_),
    .B2(_03056_),
    .Y(_06749_));
 AO21x1_ASAP7_75t_R _13702_ (.A1(_01057_),
    .A2(_04081_),
    .B(_04529_),
    .Y(_06750_));
 OA22x2_ASAP7_75t_R _13703_ (.A1(_06743_),
    .A2(_06746_),
    .B1(_06749_),
    .B2(_06750_),
    .Y(_06751_));
 AND2x2_ASAP7_75t_R _13704_ (.A(_03678_),
    .B(_01055_),
    .Y(_06752_));
 AO21x1_ASAP7_75t_R _13705_ (.A1(_03625_),
    .A2(_01054_),
    .B(_06752_),
    .Y(_06753_));
 AO21x2_ASAP7_75t_R _13706_ (.A1(_03689_),
    .A2(_06753_),
    .B(_03636_),
    .Y(_06754_));
 AND3x1_ASAP7_75t_R _13707_ (.A(_04087_),
    .B(_04692_),
    .C(_01053_),
    .Y(_06755_));
 OA21x2_ASAP7_75t_R _13708_ (.A1(_03630_),
    .A2(_04492_),
    .B(_01052_),
    .Y(_06756_));
 OA21x2_ASAP7_75t_R _13709_ (.A1(_06755_),
    .A2(_06756_),
    .B(_03635_),
    .Y(_06757_));
 AND2x2_ASAP7_75t_R _13710_ (.A(_03072_),
    .B(_01050_),
    .Y(_06758_));
 AO21x1_ASAP7_75t_R _13711_ (.A1(_03588_),
    .A2(_01048_),
    .B(_06758_),
    .Y(_06759_));
 AO22x1_ASAP7_75t_R _13712_ (.A1(_01051_),
    .A2(_03568_),
    .B1(_06759_),
    .B2(_05153_),
    .Y(_06760_));
 AO21x1_ASAP7_75t_R _13713_ (.A1(_01049_),
    .A2(_04081_),
    .B(_04082_),
    .Y(_06761_));
 OA222x2_ASAP7_75t_R _13714_ (.A1(_03959_),
    .A2(_03098_),
    .B1(_06754_),
    .B2(_06757_),
    .C1(_06760_),
    .C2(_06761_),
    .Y(_06762_));
 AOI211x1_ASAP7_75t_R _13715_ (.A1(_04098_),
    .A2(_06751_),
    .B(_06762_),
    .C(_03703_),
    .Y(_06763_));
 OAI21x1_ASAP7_75t_R _13716_ (.A1(_06740_),
    .A2(_06763_),
    .B(_03705_),
    .Y(_06764_));
 CKINVDCx20_ASAP7_75t_R _13717_ (.A(_06764_),
    .Y(net110));
 NAND2x2_ASAP7_75t_R _13718_ (.A(_03283_),
    .B(_06764_),
    .Y(_06765_));
 AO221x2_ASAP7_75t_R _13719_ (.A1(_03925_),
    .A2(_06420_),
    .B1(_06715_),
    .B2(_06419_),
    .C(_03283_),
    .Y(_06766_));
 BUFx6f_ASAP7_75t_R _13720_ (.A(_06766_),
    .Y(_06767_));
 AND2x2_ASAP7_75t_R _13721_ (.A(_06765_),
    .B(_06767_),
    .Y(_06768_));
 BUFx4f_ASAP7_75t_R _13722_ (.A(_06768_),
    .Y(_06769_));
 BUFx4f_ASAP7_75t_R _13723_ (.A(_06769_),
    .Y(_06770_));
 XNOR2x2_ASAP7_75t_R _13724_ (.A(_03259_),
    .B(_06770_),
    .Y(_09550_));
 INVx1_ASAP7_75t_R _13725_ (.A(_09550_),
    .Y(_09711_));
 INVx1_ASAP7_75t_R _13726_ (.A(_01049_),
    .Y(_06771_));
 NAND2x1_ASAP7_75t_R _13727_ (.A(_01048_),
    .B(_04005_),
    .Y(_06772_));
 OA211x2_ASAP7_75t_R _13728_ (.A1(_06771_),
    .A2(_03357_),
    .B(_03520_),
    .C(_06772_),
    .Y(_06773_));
 AND3x1_ASAP7_75t_R _13729_ (.A(_03860_),
    .B(_03970_),
    .C(_01055_),
    .Y(_06774_));
 AOI221x1_ASAP7_75t_R _13730_ (.A1(_04574_),
    .A2(_04460_),
    .B1(_03466_),
    .B2(_01054_),
    .C(_06774_),
    .Y(_06775_));
 INVx1_ASAP7_75t_R _13731_ (.A(_01051_),
    .Y(_06776_));
 OA211x2_ASAP7_75t_R _13732_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03312_),
    .C(_06776_),
    .Y(_06777_));
 NOR2x1_ASAP7_75t_R _13733_ (.A(_01050_),
    .B(_03348_),
    .Y(_06778_));
 OA211x2_ASAP7_75t_R _13734_ (.A1(_06777_),
    .A2(_06778_),
    .B(_03250_),
    .C(_03736_),
    .Y(_06779_));
 OA21x2_ASAP7_75t_R _13735_ (.A1(_06775_),
    .A2(_06779_),
    .B(_03340_),
    .Y(_06780_));
 OAI22x1_ASAP7_75t_R _13736_ (.A1(_01052_),
    .A2(_03349_),
    .B1(_03418_),
    .B2(_01053_),
    .Y(_06781_));
 AO21x1_ASAP7_75t_R _13737_ (.A1(_03361_),
    .A2(_06781_),
    .B(_03460_),
    .Y(_06782_));
 OA21x2_ASAP7_75t_R _13738_ (.A1(_06780_),
    .A2(_06782_),
    .B(_03521_),
    .Y(_06783_));
 INVx1_ASAP7_75t_R _13739_ (.A(_01057_),
    .Y(_06784_));
 NAND2x1_ASAP7_75t_R _13740_ (.A(_01056_),
    .B(_03485_),
    .Y(_06785_));
 OA211x2_ASAP7_75t_R _13741_ (.A1(_06784_),
    .A2(_04153_),
    .B(_03420_),
    .C(_06785_),
    .Y(_06786_));
 INVx1_ASAP7_75t_R _13742_ (.A(_01059_),
    .Y(_06787_));
 OA211x2_ASAP7_75t_R _13743_ (.A1(_03197_),
    .A2(_03489_),
    .B(_03347_),
    .C(_06787_),
    .Y(_06788_));
 OAI21x1_ASAP7_75t_R _13744_ (.A1(_01058_),
    .A2(_04021_),
    .B(_03320_),
    .Y(_06789_));
 OA21x2_ASAP7_75t_R _13745_ (.A1(_06788_),
    .A2(_06789_),
    .B(_03381_),
    .Y(_06790_));
 AND3x1_ASAP7_75t_R _13746_ (.A(_03031_),
    .B(_03474_),
    .C(_01063_),
    .Y(_06791_));
 AOI21x1_ASAP7_75t_R _13747_ (.A1(_01062_),
    .A2(_03436_),
    .B(_06791_),
    .Y(_06792_));
 OA22x2_ASAP7_75t_R _13748_ (.A1(_03277_),
    .A2(_06790_),
    .B1(_06792_),
    .B2(_03393_),
    .Y(_06793_));
 OAI22x1_ASAP7_75t_R _13749_ (.A1(_01061_),
    .A2(_03395_),
    .B1(_03453_),
    .B2(_01060_),
    .Y(_06794_));
 OA211x2_ASAP7_75t_R _13750_ (.A1(_03272_),
    .A2(_03286_),
    .B(_03361_),
    .C(_06794_),
    .Y(_06795_));
 OR4x1_ASAP7_75t_R _13751_ (.A(_03405_),
    .B(_06786_),
    .C(_06793_),
    .D(_06795_),
    .Y(_06796_));
 OA211x2_ASAP7_75t_R _13752_ (.A1(_06773_),
    .A2(_06783_),
    .B(_06796_),
    .C(_03495_),
    .Y(_06797_));
 NAND2x1_ASAP7_75t_R _13753_ (.A(_01032_),
    .B(_03529_),
    .Y(_06798_));
 NAND2x1_ASAP7_75t_R _13754_ (.A(_01033_),
    .B(_04466_),
    .Y(_06799_));
 OAI22x1_ASAP7_75t_R _13755_ (.A1(_01036_),
    .A2(_04023_),
    .B1(_03722_),
    .B2(_01037_),
    .Y(_06800_));
 AO32x1_ASAP7_75t_R _13756_ (.A1(_03520_),
    .A2(_06798_),
    .A3(_06799_),
    .B1(_03516_),
    .B2(_06800_),
    .Y(_06801_));
 AND3x1_ASAP7_75t_R _13757_ (.A(_03860_),
    .B(_03970_),
    .C(_01039_),
    .Y(_06802_));
 AOI221x1_ASAP7_75t_R _13758_ (.A1(_03316_),
    .A2(_04460_),
    .B1(_03466_),
    .B2(_01038_),
    .C(_06802_),
    .Y(_06803_));
 INVx1_ASAP7_75t_R _13759_ (.A(_01035_),
    .Y(_06804_));
 OA211x2_ASAP7_75t_R _13760_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03327_),
    .C(_06804_),
    .Y(_06805_));
 NOR2x1_ASAP7_75t_R _13761_ (.A(_01034_),
    .B(_03348_),
    .Y(_06806_));
 OA211x2_ASAP7_75t_R _13762_ (.A1(_06805_),
    .A2(_06806_),
    .B(_03250_),
    .C(_03387_),
    .Y(_06807_));
 OA21x2_ASAP7_75t_R _13763_ (.A1(_06803_),
    .A2(_06807_),
    .B(_03340_),
    .Y(_06808_));
 OA21x2_ASAP7_75t_R _13764_ (.A1(_03997_),
    .A2(_06808_),
    .B(_03521_),
    .Y(_06809_));
 INVx1_ASAP7_75t_R _13765_ (.A(_01041_),
    .Y(_06810_));
 NAND2x1_ASAP7_75t_R _13766_ (.A(_01040_),
    .B(_03722_),
    .Y(_06811_));
 OA211x2_ASAP7_75t_R _13767_ (.A1(_06810_),
    .A2(_04676_),
    .B(_03520_),
    .C(_06811_),
    .Y(_06812_));
 OA21x2_ASAP7_75t_R _13768_ (.A1(_01042_),
    .A2(_03507_),
    .B(_03387_),
    .Y(_06813_));
 OAI21x1_ASAP7_75t_R _13769_ (.A1(_01043_),
    .A2(_04153_),
    .B(_06813_),
    .Y(_06814_));
 AO21x1_ASAP7_75t_R _13770_ (.A1(_03381_),
    .A2(_06814_),
    .B(_03277_),
    .Y(_06815_));
 AND3x1_ASAP7_75t_R _13771_ (.A(_03860_),
    .B(_03970_),
    .C(_01047_),
    .Y(_06816_));
 AO21x1_ASAP7_75t_R _13772_ (.A1(_01046_),
    .A2(_03466_),
    .B(_06816_),
    .Y(_06817_));
 NAND2x1_ASAP7_75t_R _13773_ (.A(_03747_),
    .B(_06817_),
    .Y(_06818_));
 OAI22x1_ASAP7_75t_R _13774_ (.A1(_01045_),
    .A2(_03437_),
    .B1(_04132_),
    .B2(_01044_),
    .Y(_06819_));
 AO221x1_ASAP7_75t_R _13775_ (.A1(_06815_),
    .A2(_06818_),
    .B1(_06819_),
    .B2(_03457_),
    .C(_03405_),
    .Y(_06820_));
 OA221x2_ASAP7_75t_R _13776_ (.A1(_06801_),
    .A2(_06809_),
    .B1(_06812_),
    .B2(_06820_),
    .C(_03499_),
    .Y(_06821_));
 OR2x2_ASAP7_75t_R _13777_ (.A(_06797_),
    .B(_06821_),
    .Y(_06822_));
 BUFx4f_ASAP7_75t_R _13778_ (.A(_06822_),
    .Y(_09549_));
 INVx1_ASAP7_75t_R _13779_ (.A(_09549_),
    .Y(_09710_));
 OA22x2_ASAP7_75t_R _13780_ (.A1(_03176_),
    .A2(_03270_),
    .B1(_03281_),
    .B2(_03293_),
    .Y(_06823_));
 OR3x4_ASAP7_75t_R _13781_ (.A(_06823_),
    .B(_03427_),
    .C(_03496_),
    .Y(_06824_));
 OA21x2_ASAP7_75t_R _13782_ (.A1(_03557_),
    .A2(_03297_),
    .B(_06824_),
    .Y(_09548_));
 BUFx4f_ASAP7_75t_R _13783_ (.A(_06236_),
    .Y(_09680_));
 INVx1_ASAP7_75t_R _13784_ (.A(_09652_),
    .Y(_09650_));
 BUFx4f_ASAP7_75t_R _13785_ (.A(_05560_),
    .Y(_09645_));
 INVx1_ASAP7_75t_R _13786_ (.A(_09637_),
    .Y(_09635_));
 INVx1_ASAP7_75t_R _13787_ (.A(_09554_),
    .Y(_09551_));
 INVx2_ASAP7_75t_R _13788_ (.A(_09718_),
    .Y(net90));
 INVx4_ASAP7_75t_R _13789_ (.A(_09717_),
    .Y(net87));
 NAND2x1_ASAP7_75t_R _13790_ (.A(_03222_),
    .B(_03224_),
    .Y(_06825_));
 NOR2x2_ASAP7_75t_R _13791_ (.A(_03099_),
    .B(_03212_),
    .Y(_06826_));
 AND4x2_ASAP7_75t_R _13792_ (.A(_03217_),
    .B(_06825_),
    .C(_03229_),
    .D(_06826_),
    .Y(_06827_));
 OA21x2_ASAP7_75t_R _13793_ (.A1(_05358_),
    .A2(_03714_),
    .B(_03247_),
    .Y(_06828_));
 AND2x2_ASAP7_75t_R _13794_ (.A(_06827_),
    .B(_06828_),
    .Y(_06829_));
 BUFx6f_ASAP7_75t_R _13795_ (.A(_06829_),
    .Y(_06830_));
 BUFx6f_ASAP7_75t_R _13796_ (.A(_06830_),
    .Y(_06831_));
 AND2x2_ASAP7_75t_R _13797_ (.A(_05358_),
    .B(_06827_),
    .Y(_06832_));
 BUFx4f_ASAP7_75t_R _13798_ (.A(_06832_),
    .Y(_06833_));
 OAI21x1_ASAP7_75t_R _13799_ (.A1(_03558_),
    .A2(_09722_),
    .B(_06574_),
    .Y(_06834_));
 BUFx4f_ASAP7_75t_R _13800_ (.A(_06834_),
    .Y(_06835_));
 BUFx4f_ASAP7_75t_R _13801_ (.A(_06835_),
    .Y(_06836_));
 OAI21x1_ASAP7_75t_R _13802_ (.A1(_03558_),
    .A2(_09716_),
    .B(_06671_),
    .Y(_06837_));
 BUFx4f_ASAP7_75t_R _13803_ (.A(_06837_),
    .Y(_06838_));
 BUFx6f_ASAP7_75t_R _13804_ (.A(_06838_),
    .Y(_06839_));
 BUFx3_ASAP7_75t_R _13805_ (.A(_03295_),
    .Y(_06840_));
 NAND2x2_ASAP7_75t_R _13806_ (.A(_06765_),
    .B(_06767_),
    .Y(_06841_));
 AO221x1_ASAP7_75t_R _13807_ (.A1(_06713_),
    .A2(_04797_),
    .B1(_06765_),
    .B2(_06767_),
    .C(_04824_),
    .Y(_06842_));
 OA21x2_ASAP7_75t_R _13808_ (.A1(_09600_),
    .A2(_06841_),
    .B(_06842_),
    .Y(_06843_));
 AO221x2_ASAP7_75t_R _13809_ (.A1(_04893_),
    .A2(_04908_),
    .B1(_06765_),
    .B2(_06767_),
    .C(_04928_),
    .Y(_06844_));
 OA211x2_ASAP7_75t_R _13810_ (.A1(_09605_),
    .A2(_06841_),
    .B(_06844_),
    .C(_06823_),
    .Y(_06845_));
 AO21x1_ASAP7_75t_R _13811_ (.A1(_06840_),
    .A2(_06843_),
    .B(_06845_),
    .Y(_06846_));
 BUFx3_ASAP7_75t_R _13812_ (.A(_06841_),
    .Y(_06847_));
 BUFx4f_ASAP7_75t_R _13813_ (.A(_06765_),
    .Y(_06848_));
 BUFx4f_ASAP7_75t_R _13814_ (.A(_06767_),
    .Y(_06849_));
 AO211x2_ASAP7_75t_R _13815_ (.A1(_06848_),
    .A2(_06849_),
    .B(_05333_),
    .C(_05357_),
    .Y(_06850_));
 BUFx3_ASAP7_75t_R _13816_ (.A(_06823_),
    .Y(_06851_));
 OA211x2_ASAP7_75t_R _13817_ (.A1(_09625_),
    .A2(_06847_),
    .B(_06850_),
    .C(_06851_),
    .Y(_06852_));
 AOI221x1_ASAP7_75t_R _13818_ (.A1(_05202_),
    .A2(_05212_),
    .B1(_05214_),
    .B2(_05223_),
    .C(_04003_),
    .Y(_06853_));
 AND3x2_ASAP7_75t_R _13819_ (.A(_06713_),
    .B(_05234_),
    .C(_05246_),
    .Y(_06854_));
 AO211x2_ASAP7_75t_R _13820_ (.A1(_06848_),
    .A2(_06849_),
    .B(_06853_),
    .C(_06854_),
    .Y(_06855_));
 BUFx3_ASAP7_75t_R _13821_ (.A(_03294_),
    .Y(_06856_));
 OA211x2_ASAP7_75t_R _13822_ (.A1(_09620_),
    .A2(_06847_),
    .B(_06855_),
    .C(_06856_),
    .Y(_06857_));
 OR3x1_ASAP7_75t_R _13823_ (.A(_06673_),
    .B(_06852_),
    .C(_06857_),
    .Y(_06858_));
 OA21x2_ASAP7_75t_R _13824_ (.A1(_06839_),
    .A2(_06846_),
    .B(_06858_),
    .Y(_06859_));
 BUFx4f_ASAP7_75t_R _13825_ (.A(_06838_),
    .Y(_06860_));
 BUFx4f_ASAP7_75t_R _13826_ (.A(_06823_),
    .Y(_06861_));
 BUFx4f_ASAP7_75t_R _13827_ (.A(_06841_),
    .Y(_06862_));
 NAND2x1_ASAP7_75t_R _13828_ (.A(_09577_),
    .B(_06862_),
    .Y(_06863_));
 OR2x2_ASAP7_75t_R _13829_ (.A(_09565_),
    .B(_06841_),
    .Y(_06864_));
 AO211x2_ASAP7_75t_R _13830_ (.A1(_06765_),
    .A2(_06767_),
    .B(_03864_),
    .C(_03890_),
    .Y(_06865_));
 OA211x2_ASAP7_75t_R _13831_ (.A1(_03554_),
    .A2(_06841_),
    .B(_06865_),
    .C(_03295_),
    .Y(_06866_));
 AO31x2_ASAP7_75t_R _13832_ (.A1(_06861_),
    .A2(_06863_),
    .A3(_06864_),
    .B(_06866_),
    .Y(_06867_));
 BUFx4f_ASAP7_75t_R _13833_ (.A(_06673_),
    .Y(_06868_));
 BUFx4f_ASAP7_75t_R _13834_ (.A(_06768_),
    .Y(_06869_));
 AND2x4_ASAP7_75t_R _13835_ (.A(_03283_),
    .B(_06764_),
    .Y(_06870_));
 AOI221x1_ASAP7_75t_R _13836_ (.A1(_03925_),
    .A2(_06420_),
    .B1(_06715_),
    .B2(_06419_),
    .C(_03283_),
    .Y(_06871_));
 OR4x1_ASAP7_75t_R _13837_ (.A(_04239_),
    .B(_04265_),
    .C(_06870_),
    .D(_06871_),
    .Y(_06872_));
 OA211x2_ASAP7_75t_R _13838_ (.A1(_09595_),
    .A2(_06869_),
    .B(_06872_),
    .C(_06823_),
    .Y(_06873_));
 AO211x2_ASAP7_75t_R _13839_ (.A1(_06765_),
    .A2(_06767_),
    .B(_04338_),
    .C(_04359_),
    .Y(_06874_));
 OA211x2_ASAP7_75t_R _13840_ (.A1(_09580_),
    .A2(_06841_),
    .B(_06874_),
    .C(_03294_),
    .Y(_06875_));
 OR3x1_ASAP7_75t_R _13841_ (.A(_06868_),
    .B(_06873_),
    .C(_06875_),
    .Y(_06876_));
 OA211x2_ASAP7_75t_R _13842_ (.A1(_06860_),
    .A2(_06867_),
    .B(_06876_),
    .C(_06576_),
    .Y(_06877_));
 AO21x1_ASAP7_75t_R _13843_ (.A1(_06836_),
    .A2(_06859_),
    .B(_06877_),
    .Y(_06878_));
 AND2x2_ASAP7_75t_R _13844_ (.A(_06833_),
    .B(_06878_),
    .Y(_06879_));
 BUFx4f_ASAP7_75t_R _13845_ (.A(_06834_),
    .Y(_06880_));
 BUFx4f_ASAP7_75t_R _13846_ (.A(_06880_),
    .Y(_06881_));
 BUFx4f_ASAP7_75t_R _13847_ (.A(_06881_),
    .Y(_06882_));
 BUFx6f_ASAP7_75t_R _13848_ (.A(_06861_),
    .Y(_06883_));
 AO221x1_ASAP7_75t_R _13849_ (.A1(_05032_),
    .A2(_06597_),
    .B1(_06616_),
    .B2(_06713_),
    .C(_06883_),
    .Y(_06884_));
 OA21x2_ASAP7_75t_R _13850_ (.A1(_03297_),
    .A2(_09705_),
    .B(_06884_),
    .Y(_06885_));
 AND3x2_ASAP7_75t_R _13851_ (.A(_06840_),
    .B(_06847_),
    .C(_09549_),
    .Y(_06886_));
 AO21x1_ASAP7_75t_R _13852_ (.A1(_06770_),
    .A2(_06885_),
    .B(_06886_),
    .Y(_06887_));
 BUFx4f_ASAP7_75t_R _13853_ (.A(_06841_),
    .Y(_06888_));
 AND3x2_ASAP7_75t_R _13854_ (.A(_06861_),
    .B(_09555_),
    .C(_06888_),
    .Y(_06889_));
 AOI21x1_ASAP7_75t_R _13855_ (.A1(_06833_),
    .A2(_06887_),
    .B(_06889_),
    .Y(_06890_));
 BUFx4f_ASAP7_75t_R _13856_ (.A(_06860_),
    .Y(_06891_));
 NAND2x2_ASAP7_75t_R _13857_ (.A(_05358_),
    .B(_06827_),
    .Y(_06892_));
 BUFx4f_ASAP7_75t_R _13858_ (.A(_06892_),
    .Y(_06893_));
 BUFx4f_ASAP7_75t_R _13859_ (.A(_06869_),
    .Y(_06894_));
 AND2x2_ASAP7_75t_R _13860_ (.A(_09680_),
    .B(_06894_),
    .Y(_06895_));
 BUFx4f_ASAP7_75t_R _13861_ (.A(_06841_),
    .Y(_06896_));
 BUFx4f_ASAP7_75t_R _13862_ (.A(_06823_),
    .Y(_06897_));
 BUFx3_ASAP7_75t_R _13863_ (.A(_06897_),
    .Y(_06898_));
 AO21x1_ASAP7_75t_R _13864_ (.A1(_09690_),
    .A2(_06896_),
    .B(_06898_),
    .Y(_06899_));
 AOI22x1_ASAP7_75t_R _13865_ (.A1(_06499_),
    .A2(_06528_),
    .B1(_06848_),
    .B2(_06849_),
    .Y(_06900_));
 AO21x1_ASAP7_75t_R _13866_ (.A1(_09685_),
    .A2(_06894_),
    .B(_06900_),
    .Y(_06901_));
 BUFx4f_ASAP7_75t_R _13867_ (.A(_06840_),
    .Y(_06902_));
 OAI22x1_ASAP7_75t_R _13868_ (.A1(_06895_),
    .A2(_06899_),
    .B1(_06901_),
    .B2(_06902_),
    .Y(_06903_));
 OR3x1_ASAP7_75t_R _13869_ (.A(_06891_),
    .B(_06893_),
    .C(_06903_),
    .Y(_06904_));
 OAI21x1_ASAP7_75t_R _13870_ (.A1(_06675_),
    .A2(_06890_),
    .B(_06904_),
    .Y(_06905_));
 OR3x2_ASAP7_75t_R _13871_ (.A(_05442_),
    .B(_05465_),
    .C(_06847_),
    .Y(_06906_));
 NAND2x2_ASAP7_75t_R _13872_ (.A(_09652_),
    .B(_06896_),
    .Y(_06907_));
 AOI221x1_ASAP7_75t_R _13873_ (.A1(_05721_),
    .A2(_05728_),
    .B1(_05730_),
    .B2(_05742_),
    .C(_03426_),
    .Y(_06908_));
 AND3x1_ASAP7_75t_R _13874_ (.A(_05032_),
    .B(_05755_),
    .C(_05773_),
    .Y(_06909_));
 AO211x2_ASAP7_75t_R _13875_ (.A1(_06848_),
    .A2(_06849_),
    .B(_06908_),
    .C(_06909_),
    .Y(_06910_));
 OA211x2_ASAP7_75t_R _13876_ (.A1(_09645_),
    .A2(_06847_),
    .B(_06910_),
    .C(_06851_),
    .Y(_06911_));
 AO31x2_ASAP7_75t_R _13877_ (.A1(_06902_),
    .A2(_06906_),
    .A3(_06907_),
    .B(_06911_),
    .Y(_06912_));
 AO221x2_ASAP7_75t_R _13878_ (.A1(_06713_),
    .A2(_06118_),
    .B1(_06848_),
    .B2(_06849_),
    .C(_06145_),
    .Y(_06913_));
 OA211x2_ASAP7_75t_R _13879_ (.A1(_09665_),
    .A2(_06888_),
    .B(_06913_),
    .C(_06851_),
    .Y(_06914_));
 AO211x2_ASAP7_75t_R _13880_ (.A1(_06848_),
    .A2(_06849_),
    .B(_06030_),
    .C(_06050_),
    .Y(_06915_));
 OA211x2_ASAP7_75t_R _13881_ (.A1(_09660_),
    .A2(_06847_),
    .B(_06915_),
    .C(_06856_),
    .Y(_06916_));
 OR3x1_ASAP7_75t_R _13882_ (.A(_06673_),
    .B(_06914_),
    .C(_06916_),
    .Y(_06917_));
 OA21x2_ASAP7_75t_R _13883_ (.A1(_06839_),
    .A2(_06912_),
    .B(_06917_),
    .Y(_06918_));
 AND2x2_ASAP7_75t_R _13884_ (.A(_06576_),
    .B(_06832_),
    .Y(_06919_));
 AO21x2_ASAP7_75t_R _13885_ (.A1(_03558_),
    .A2(net125),
    .B(_06468_),
    .Y(_06920_));
 BUFx4f_ASAP7_75t_R _13886_ (.A(_06920_),
    .Y(_06921_));
 AO221x1_ASAP7_75t_R _13887_ (.A1(_06882_),
    .A2(_06905_),
    .B1(_06918_),
    .B2(_06919_),
    .C(_06921_),
    .Y(_06922_));
 OAI21x1_ASAP7_75t_R _13888_ (.A1(_06472_),
    .A2(_06879_),
    .B(_06922_),
    .Y(_06923_));
 NAND2x2_ASAP7_75t_R _13889_ (.A(_06827_),
    .B(_06828_),
    .Y(_06924_));
 BUFx4f_ASAP7_75t_R _13890_ (.A(_06924_),
    .Y(_06925_));
 AND3x2_ASAP7_75t_R _13891_ (.A(_03199_),
    .B(_03202_),
    .C(_03210_),
    .Y(_06926_));
 INVx1_ASAP7_75t_R _13892_ (.A(net6),
    .Y(_06927_));
 AND2x2_ASAP7_75t_R _13893_ (.A(_06927_),
    .B(_03217_),
    .Y(_06928_));
 INVx1_ASAP7_75t_R _13894_ (.A(_03217_),
    .Y(_06929_));
 AND2x2_ASAP7_75t_R _13895_ (.A(net6),
    .B(_06929_),
    .Y(_06930_));
 OR3x1_ASAP7_75t_R _13896_ (.A(_03212_),
    .B(_06928_),
    .C(_06930_),
    .Y(_06931_));
 OA211x2_ASAP7_75t_R _13897_ (.A1(net6),
    .A2(net22),
    .B(_06931_),
    .C(_03023_),
    .Y(_06932_));
 INVx1_ASAP7_75t_R _13898_ (.A(_06932_),
    .Y(_06933_));
 AO21x2_ASAP7_75t_R _13899_ (.A1(_06926_),
    .A2(_06933_),
    .B(_03257_),
    .Y(_06934_));
 BUFx4f_ASAP7_75t_R _13900_ (.A(_06825_),
    .Y(_06935_));
 AO21x1_ASAP7_75t_R _13901_ (.A1(_03217_),
    .A2(_03230_),
    .B(net6),
    .Y(_06936_));
 AO32x1_ASAP7_75t_R _13902_ (.A1(_06935_),
    .A2(_03229_),
    .A3(_06930_),
    .B1(_06936_),
    .B2(_03212_),
    .Y(_06937_));
 AOI21x1_ASAP7_75t_R _13903_ (.A1(_03024_),
    .A2(_06937_),
    .B(_06926_),
    .Y(_06938_));
 NOR2x2_ASAP7_75t_R _13904_ (.A(_06934_),
    .B(_06938_),
    .Y(_06939_));
 BUFx4f_ASAP7_75t_R _13905_ (.A(_06939_),
    .Y(_06940_));
 AO21x2_ASAP7_75t_R _13906_ (.A1(net22),
    .A2(_06926_),
    .B(_03230_),
    .Y(_06941_));
 NAND2x2_ASAP7_75t_R _13907_ (.A(_03023_),
    .B(_03212_),
    .Y(_06942_));
 AO21x2_ASAP7_75t_R _13908_ (.A1(_05358_),
    .A2(_03217_),
    .B(_06942_),
    .Y(_06943_));
 OR2x2_ASAP7_75t_R _13909_ (.A(_00499_),
    .B(_00532_),
    .Y(_06944_));
 INVx2_ASAP7_75t_R _13910_ (.A(_00932_),
    .Y(_06945_));
 INVx1_ASAP7_75t_R _13911_ (.A(_00965_),
    .Y(_06946_));
 INVx1_ASAP7_75t_R _13912_ (.A(_00998_),
    .Y(_06947_));
 OAI21x1_ASAP7_75t_R _13913_ (.A1(net163),
    .A2(_01158_),
    .B(_01212_),
    .Y(_06948_));
 INVx1_ASAP7_75t_R _13914_ (.A(_01210_),
    .Y(_06949_));
 AO21x1_ASAP7_75t_R _13915_ (.A1(_06947_),
    .A2(_06948_),
    .B(_06949_),
    .Y(_06950_));
 INVx1_ASAP7_75t_R _13916_ (.A(_01208_),
    .Y(_06951_));
 AO21x1_ASAP7_75t_R _13917_ (.A1(_06946_),
    .A2(_06950_),
    .B(_06951_),
    .Y(_06952_));
 INVx1_ASAP7_75t_R _13918_ (.A(_00931_),
    .Y(_06953_));
 AOI21x1_ASAP7_75t_R _13919_ (.A1(_06945_),
    .A2(_06952_),
    .B(_06953_),
    .Y(_06954_));
 OA21x2_ASAP7_75t_R _13920_ (.A1(_00898_),
    .A2(_06954_),
    .B(_01205_),
    .Y(_06955_));
 BUFx3_ASAP7_75t_R _13921_ (.A(_00764_),
    .Y(_06956_));
 OR3x4_ASAP7_75t_R _13922_ (.A(_00798_),
    .B(_00831_),
    .C(_00865_),
    .Y(_06957_));
 OR3x1_ASAP7_75t_R _13923_ (.A(_00731_),
    .B(_06956_),
    .C(_06957_),
    .Y(_06958_));
 OA21x2_ASAP7_75t_R _13924_ (.A1(_00831_),
    .A2(_00864_),
    .B(_01202_),
    .Y(_06959_));
 OA21x2_ASAP7_75t_R _13925_ (.A1(_00798_),
    .A2(_06959_),
    .B(_00797_),
    .Y(_06960_));
 OR3x1_ASAP7_75t_R _13926_ (.A(_00731_),
    .B(_06956_),
    .C(_06960_),
    .Y(_06961_));
 OA21x2_ASAP7_75t_R _13927_ (.A1(_00731_),
    .A2(_01199_),
    .B(_06961_),
    .Y(_06962_));
 OA21x2_ASAP7_75t_R _13928_ (.A1(_00632_),
    .A2(_01193_),
    .B(_01191_),
    .Y(_06963_));
 OA21x2_ASAP7_75t_R _13929_ (.A1(_00599_),
    .A2(_06963_),
    .B(_00598_),
    .Y(_06964_));
 AND3x1_ASAP7_75t_R _13930_ (.A(_01195_),
    .B(_01197_),
    .C(_06964_),
    .Y(_06965_));
 OA211x2_ASAP7_75t_R _13931_ (.A1(_06955_),
    .A2(_06958_),
    .B(_06962_),
    .C(_06965_),
    .Y(_06966_));
 OR3x1_ASAP7_75t_R _13932_ (.A(_00599_),
    .B(_00632_),
    .C(_00665_),
    .Y(_06967_));
 AND3x1_ASAP7_75t_R _13933_ (.A(_00698_),
    .B(_01195_),
    .C(_06964_),
    .Y(_06968_));
 AO21x1_ASAP7_75t_R _13934_ (.A1(_06964_),
    .A2(_06967_),
    .B(_06968_),
    .Y(_06969_));
 OR4x1_ASAP7_75t_R _13935_ (.A(_00565_),
    .B(_06944_),
    .C(_06966_),
    .D(_06969_),
    .Y(_06970_));
 OA21x2_ASAP7_75t_R _13936_ (.A1(_00499_),
    .A2(_01186_),
    .B(_01184_),
    .Y(_06971_));
 OA21x2_ASAP7_75t_R _13937_ (.A1(_01188_),
    .A2(_06944_),
    .B(_06971_),
    .Y(_06972_));
 OR2x2_ASAP7_75t_R _13938_ (.A(_00433_),
    .B(_00466_),
    .Y(_06973_));
 OR2x2_ASAP7_75t_R _13939_ (.A(_00367_),
    .B(_00400_),
    .Y(_06974_));
 OR2x2_ASAP7_75t_R _13940_ (.A(_06973_),
    .B(_06974_),
    .Y(_06975_));
 AO21x1_ASAP7_75t_R _13941_ (.A1(_06970_),
    .A2(_06972_),
    .B(_06975_),
    .Y(_06976_));
 OA21x2_ASAP7_75t_R _13942_ (.A1(_00433_),
    .A2(_01182_),
    .B(_01180_),
    .Y(_06977_));
 OA21x2_ASAP7_75t_R _13943_ (.A1(_00400_),
    .A2(_06977_),
    .B(_01178_),
    .Y(_06978_));
 OA21x2_ASAP7_75t_R _13944_ (.A1(_00367_),
    .A2(_06978_),
    .B(_01176_),
    .Y(_06979_));
 AND2x2_ASAP7_75t_R _13945_ (.A(_00333_),
    .B(_06979_),
    .Y(_06980_));
 AO221x1_ASAP7_75t_R _13946_ (.A1(_00334_),
    .A2(_00333_),
    .B1(_06976_),
    .B2(_06980_),
    .C(_00300_),
    .Y(_06981_));
 BUFx3_ASAP7_75t_R _13947_ (.A(_00167_),
    .Y(_06982_));
 OR3x1_ASAP7_75t_R _13948_ (.A(_00234_),
    .B(_00267_),
    .C(_01168_),
    .Y(_06983_));
 OR4x1_ASAP7_75t_R _13949_ (.A(_00100_),
    .B(_06982_),
    .C(_01165_),
    .D(_06983_),
    .Y(_06984_));
 OA21x2_ASAP7_75t_R _13950_ (.A1(_00267_),
    .A2(_01173_),
    .B(_01171_),
    .Y(_06985_));
 OA21x2_ASAP7_75t_R _13951_ (.A1(_00234_),
    .A2(_06985_),
    .B(_00233_),
    .Y(_06986_));
 OA21x2_ASAP7_75t_R _13952_ (.A1(_01168_),
    .A2(_06986_),
    .B(_00200_),
    .Y(_06987_));
 OR2x2_ASAP7_75t_R _13953_ (.A(_06982_),
    .B(_06987_),
    .Y(_06988_));
 AO21x1_ASAP7_75t_R _13954_ (.A1(_00166_),
    .A2(_06988_),
    .B(_01165_),
    .Y(_06989_));
 AO21x1_ASAP7_75t_R _13955_ (.A1(_00133_),
    .A2(_06989_),
    .B(_00100_),
    .Y(_06990_));
 OA211x2_ASAP7_75t_R _13956_ (.A1(_06981_),
    .A2(_06984_),
    .B(_06990_),
    .C(_00099_),
    .Y(_06991_));
 OA21x2_ASAP7_75t_R _13957_ (.A1(_01162_),
    .A2(_06991_),
    .B(_01161_),
    .Y(_06992_));
 NAND2x1_ASAP7_75t_R _13958_ (.A(_05468_),
    .B(_06928_),
    .Y(_06993_));
 XNOR2x1_ASAP7_75t_R _13959_ (.B(_03644_),
    .Y(_06994_),
    .A(_03554_));
 OA21x2_ASAP7_75t_R _13960_ (.A1(_06941_),
    .A2(_06993_),
    .B(_06994_),
    .Y(_06995_));
 XNOR2x1_ASAP7_75t_R _13961_ (.B(_06995_),
    .Y(_06996_),
    .A(_03556_));
 XNOR2x1_ASAP7_75t_R _13962_ (.B(_06996_),
    .Y(_06997_),
    .A(_06992_));
 OR5x1_ASAP7_75t_R _13963_ (.A(_03257_),
    .B(_06940_),
    .C(_06941_),
    .D(_06943_),
    .E(_06997_),
    .Y(_06998_));
 NOR3x2_ASAP7_75t_R _13964_ (.B(_06941_),
    .C(_06943_),
    .Y(_06999_),
    .A(_03257_));
 NAND2x2_ASAP7_75t_R _13965_ (.A(_06826_),
    .B(_06930_),
    .Y(_07000_));
 NOR3x2_ASAP7_75t_R _13966_ (.B(_06941_),
    .C(_07000_),
    .Y(_07001_),
    .A(_03257_));
 OR2x2_ASAP7_75t_R _13967_ (.A(_06999_),
    .B(_07001_),
    .Y(_07002_));
 NOR2x1_ASAP7_75t_R _13968_ (.A(_06939_),
    .B(_07002_),
    .Y(_07003_));
 BUFx4f_ASAP7_75t_R _13969_ (.A(_07003_),
    .Y(_07004_));
 BUFx4f_ASAP7_75t_R _13970_ (.A(_07001_),
    .Y(_07005_));
 AO21x1_ASAP7_75t_R _13971_ (.A1(_03259_),
    .A2(_07004_),
    .B(_07005_),
    .Y(_07006_));
 OR2x2_ASAP7_75t_R _13972_ (.A(_06939_),
    .B(_07002_),
    .Y(_07007_));
 BUFx3_ASAP7_75t_R _13973_ (.A(_07007_),
    .Y(_07008_));
 BUFx6f_ASAP7_75t_R _13974_ (.A(_07008_),
    .Y(_07009_));
 OAI21x1_ASAP7_75t_R _13975_ (.A1(_03259_),
    .A2(_07009_),
    .B(_00034_),
    .Y(_07010_));
 OAI21x1_ASAP7_75t_R _13976_ (.A1(_00034_),
    .A2(_07006_),
    .B(_07010_),
    .Y(_07011_));
 BUFx3_ASAP7_75t_R _13977_ (.A(_06999_),
    .Y(_07012_));
 NOR2x2_ASAP7_75t_R _13978_ (.A(_06999_),
    .B(_07001_),
    .Y(_07013_));
 BUFx3_ASAP7_75t_R _13979_ (.A(_07013_),
    .Y(_07014_));
 INVx1_ASAP7_75t_R _13980_ (.A(_01160_),
    .Y(_07015_));
 AO22x1_ASAP7_75t_R _13981_ (.A1(_01064_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07015_),
    .Y(_07016_));
 NAND2x1_ASAP7_75t_R _13982_ (.A(_06940_),
    .B(_07016_),
    .Y(_07017_));
 AND4x1_ASAP7_75t_R _13983_ (.A(_06925_),
    .B(_06998_),
    .C(_07011_),
    .D(_07017_),
    .Y(_07018_));
 AOI21x1_ASAP7_75t_R _13984_ (.A1(_06831_),
    .A2(_06923_),
    .B(_07018_),
    .Y(net32));
 BUFx6f_ASAP7_75t_R _13985_ (.A(_06924_),
    .Y(_07019_));
 BUFx4f_ASAP7_75t_R _13986_ (.A(_06920_),
    .Y(_07020_));
 BUFx4f_ASAP7_75t_R _13987_ (.A(_07020_),
    .Y(_07021_));
 BUFx4f_ASAP7_75t_R _13988_ (.A(_06837_),
    .Y(_07022_));
 BUFx4f_ASAP7_75t_R _13989_ (.A(_07022_),
    .Y(_07023_));
 AO221x2_ASAP7_75t_R _13990_ (.A1(_04673_),
    .A2(_04687_),
    .B1(_06765_),
    .B2(_06767_),
    .C(_04714_),
    .Y(_07024_));
 OA211x2_ASAP7_75t_R _13991_ (.A1(_09595_),
    .A2(_06888_),
    .B(_07024_),
    .C(_06840_),
    .Y(_07025_));
 AO21x1_ASAP7_75t_R _13992_ (.A1(_06883_),
    .A2(_06843_),
    .B(_07025_),
    .Y(_07026_));
 BUFx4f_ASAP7_75t_R _13993_ (.A(_06673_),
    .Y(_07027_));
 BUFx3_ASAP7_75t_R _13994_ (.A(_06862_),
    .Y(_07028_));
 BUFx4f_ASAP7_75t_R _13995_ (.A(_06851_),
    .Y(_07029_));
 OA211x2_ASAP7_75t_R _13996_ (.A1(_09620_),
    .A2(_07028_),
    .B(_06855_),
    .C(_07029_),
    .Y(_07030_));
 AO221x2_ASAP7_75t_R _13997_ (.A1(_05111_),
    .A2(_05120_),
    .B1(_06848_),
    .B2(_06849_),
    .C(_05145_),
    .Y(_07031_));
 OA211x2_ASAP7_75t_R _13998_ (.A1(_09615_),
    .A2(_07028_),
    .B(_07031_),
    .C(_03296_),
    .Y(_07032_));
 OR3x1_ASAP7_75t_R _13999_ (.A(_07027_),
    .B(_07030_),
    .C(_07032_),
    .Y(_07033_));
 OA21x2_ASAP7_75t_R _14000_ (.A1(_07023_),
    .A2(_07026_),
    .B(_07033_),
    .Y(_07034_));
 AND2x2_ASAP7_75t_R _14001_ (.A(_06881_),
    .B(_07034_),
    .Y(_07035_));
 BUFx4f_ASAP7_75t_R _14002_ (.A(_06576_),
    .Y(_07036_));
 BUFx4f_ASAP7_75t_R _14003_ (.A(_07036_),
    .Y(_07037_));
 OA211x2_ASAP7_75t_R _14004_ (.A1(_09580_),
    .A2(_06888_),
    .B(_06874_),
    .C(_06851_),
    .Y(_07038_));
 AO211x2_ASAP7_75t_R _14005_ (.A1(_06848_),
    .A2(_06849_),
    .B(_04239_),
    .C(_04265_),
    .Y(_07039_));
 OA211x2_ASAP7_75t_R _14006_ (.A1(_09575_),
    .A2(_06888_),
    .B(_07039_),
    .C(_06840_),
    .Y(_07040_));
 OR3x2_ASAP7_75t_R _14007_ (.A(_06868_),
    .B(_07038_),
    .C(_07040_),
    .Y(_07041_));
 BUFx4f_ASAP7_75t_R _14008_ (.A(_06838_),
    .Y(_07042_));
 BUFx4f_ASAP7_75t_R _14009_ (.A(_07042_),
    .Y(_07043_));
 BUFx4f_ASAP7_75t_R _14010_ (.A(_06888_),
    .Y(_07044_));
 OR3x1_ASAP7_75t_R _14011_ (.A(_06856_),
    .B(_03864_),
    .C(_03890_),
    .Y(_07045_));
 OA21x2_ASAP7_75t_R _14012_ (.A1(_07029_),
    .A2(_09565_),
    .B(_07045_),
    .Y(_07046_));
 AND2x2_ASAP7_75t_R _14013_ (.A(_07044_),
    .B(_07046_),
    .Y(_07047_));
 BUFx4f_ASAP7_75t_R _14014_ (.A(_07029_),
    .Y(_07048_));
 AND3x4_ASAP7_75t_R _14015_ (.A(_03024_),
    .B(net22),
    .C(_06832_),
    .Y(_07049_));
 AND2x2_ASAP7_75t_R _14016_ (.A(_03555_),
    .B(_06770_),
    .Y(_07050_));
 OA21x2_ASAP7_75t_R _14017_ (.A1(_07048_),
    .A2(_07049_),
    .B(_07050_),
    .Y(_07051_));
 OR3x1_ASAP7_75t_R _14018_ (.A(_07043_),
    .B(_07047_),
    .C(_07051_),
    .Y(_07052_));
 AND3x1_ASAP7_75t_R _14019_ (.A(_07037_),
    .B(_07041_),
    .C(_07052_),
    .Y(_07053_));
 BUFx4f_ASAP7_75t_R _14020_ (.A(_06833_),
    .Y(_07054_));
 OAI21x1_ASAP7_75t_R _14021_ (.A1(_07035_),
    .A2(_07053_),
    .B(_07054_),
    .Y(_07055_));
 BUFx4f_ASAP7_75t_R _14022_ (.A(_06892_),
    .Y(_07056_));
 AND2x2_ASAP7_75t_R _14023_ (.A(_07022_),
    .B(_07044_),
    .Y(_07057_));
 OR3x1_ASAP7_75t_R _14024_ (.A(_06840_),
    .B(_06797_),
    .C(_06821_),
    .Y(_07058_));
 AND2x2_ASAP7_75t_R _14025_ (.A(_06824_),
    .B(_07058_),
    .Y(_07059_));
 AND2x2_ASAP7_75t_R _14026_ (.A(_07057_),
    .B(_07059_),
    .Y(_07060_));
 BUFx4f_ASAP7_75t_R _14027_ (.A(_06862_),
    .Y(_07061_));
 BUFx4f_ASAP7_75t_R _14028_ (.A(_07061_),
    .Y(_07062_));
 BUFx4f_ASAP7_75t_R _14029_ (.A(_06861_),
    .Y(_07063_));
 OR3x1_ASAP7_75t_R _14030_ (.A(_03295_),
    .B(_06392_),
    .C(_06417_),
    .Y(_07064_));
 OA21x2_ASAP7_75t_R _14031_ (.A1(_07063_),
    .A2(_09685_),
    .B(_07064_),
    .Y(_07065_));
 BUFx3_ASAP7_75t_R _14032_ (.A(_06869_),
    .Y(_07066_));
 AO211x2_ASAP7_75t_R _14033_ (.A1(_06713_),
    .A2(_06118_),
    .B(_06145_),
    .C(_06861_),
    .Y(_07067_));
 OA211x2_ASAP7_75t_R _14034_ (.A1(_06902_),
    .A2(_09680_),
    .B(_07066_),
    .C(_07067_),
    .Y(_07068_));
 AO21x1_ASAP7_75t_R _14035_ (.A1(_07062_),
    .A2(_07065_),
    .B(_07068_),
    .Y(_07069_));
 NOR3x2_ASAP7_75t_R _14036_ (.B(_06486_),
    .C(_06498_),
    .Y(_07070_),
    .A(_03426_));
 OA21x2_ASAP7_75t_R _14037_ (.A1(_06507_),
    .A2(_06514_),
    .B(_06527_),
    .Y(_07071_));
 OR3x1_ASAP7_75t_R _14038_ (.A(_06897_),
    .B(_07070_),
    .C(_07071_),
    .Y(_07072_));
 OA211x2_ASAP7_75t_R _14039_ (.A1(_03296_),
    .A2(_09700_),
    .B(_07066_),
    .C(_07072_),
    .Y(_07073_));
 OA211x2_ASAP7_75t_R _14040_ (.A1(_06883_),
    .A2(_09705_),
    .B(_07061_),
    .C(_07058_),
    .Y(_07074_));
 OR3x1_ASAP7_75t_R _14041_ (.A(_07027_),
    .B(_07073_),
    .C(_07074_),
    .Y(_07075_));
 BUFx4f_ASAP7_75t_R _14042_ (.A(_06832_),
    .Y(_07076_));
 OA211x2_ASAP7_75t_R _14043_ (.A1(_07043_),
    .A2(_07069_),
    .B(_07075_),
    .C(_07076_),
    .Y(_07077_));
 AOI21x1_ASAP7_75t_R _14044_ (.A1(_07056_),
    .A2(_07060_),
    .B(_07077_),
    .Y(_07078_));
 OR4x2_ASAP7_75t_R _14045_ (.A(_05333_),
    .B(_05357_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07079_));
 OA211x2_ASAP7_75t_R _14046_ (.A1(_09645_),
    .A2(_07066_),
    .B(_07079_),
    .C(_03296_),
    .Y(_07080_));
 AO31x2_ASAP7_75t_R _14047_ (.A1(_07048_),
    .A2(_06906_),
    .A3(_06907_),
    .B(_07080_),
    .Y(_07081_));
 OA211x2_ASAP7_75t_R _14048_ (.A1(_09660_),
    .A2(_07061_),
    .B(_06915_),
    .C(_07029_),
    .Y(_07082_));
 OR4x2_ASAP7_75t_R _14049_ (.A(_06908_),
    .B(_06909_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07083_));
 OA211x2_ASAP7_75t_R _14050_ (.A1(_09665_),
    .A2(_07066_),
    .B(_07083_),
    .C(_03296_),
    .Y(_07084_));
 OR3x1_ASAP7_75t_R _14051_ (.A(_06674_),
    .B(_07082_),
    .C(_07084_),
    .Y(_07085_));
 OA21x2_ASAP7_75t_R _14052_ (.A1(_07043_),
    .A2(_07081_),
    .B(_07085_),
    .Y(_07086_));
 NAND2x1_ASAP7_75t_R _14053_ (.A(_06919_),
    .B(_07086_),
    .Y(_07087_));
 BUFx4f_ASAP7_75t_R _14054_ (.A(_06470_),
    .Y(_07088_));
 OA211x2_ASAP7_75t_R _14055_ (.A1(_06578_),
    .A2(_07078_),
    .B(_07087_),
    .C(_07088_),
    .Y(_07089_));
 AO21x1_ASAP7_75t_R _14056_ (.A1(_07021_),
    .A2(_07055_),
    .B(_07089_),
    .Y(_07090_));
 BUFx4f_ASAP7_75t_R _14057_ (.A(_06939_),
    .Y(_07091_));
 BUFx3_ASAP7_75t_R _14058_ (.A(_07012_),
    .Y(_07092_));
 BUFx4f_ASAP7_75t_R _14059_ (.A(_07001_),
    .Y(_07093_));
 INVx1_ASAP7_75t_R _14060_ (.A(_01215_),
    .Y(_07094_));
 AO32x1_ASAP7_75t_R _14061_ (.A1(_01216_),
    .A2(_07091_),
    .A3(_07092_),
    .B1(_07093_),
    .B2(_07094_),
    .Y(_07095_));
 INVx1_ASAP7_75t_R _14062_ (.A(_01065_),
    .Y(_07096_));
 BUFx3_ASAP7_75t_R _14063_ (.A(_07014_),
    .Y(_07097_));
 INVx1_ASAP7_75t_R _14064_ (.A(_01214_),
    .Y(_07098_));
 OR3x1_ASAP7_75t_R _14065_ (.A(_07098_),
    .B(_06934_),
    .C(_06938_),
    .Y(_07099_));
 OA211x2_ASAP7_75t_R _14066_ (.A1(_07096_),
    .A2(_07091_),
    .B(_07097_),
    .C(_07099_),
    .Y(_07100_));
 OAI21x1_ASAP7_75t_R _14067_ (.A1(_07095_),
    .A2(_07100_),
    .B(_07019_),
    .Y(_07101_));
 OAI21x1_ASAP7_75t_R _14068_ (.A1(_07019_),
    .A2(_07090_),
    .B(_07101_),
    .Y(net43));
 OR2x2_ASAP7_75t_R _14069_ (.A(_09610_),
    .B(_06862_),
    .Y(_07102_));
 OR2x2_ASAP7_75t_R _14070_ (.A(_09620_),
    .B(_06869_),
    .Y(_07103_));
 OA211x2_ASAP7_75t_R _14071_ (.A1(_09615_),
    .A2(_06862_),
    .B(_07031_),
    .C(_06851_),
    .Y(_07104_));
 AO31x2_ASAP7_75t_R _14072_ (.A1(_03296_),
    .A2(_07102_),
    .A3(_07103_),
    .B(_07104_),
    .Y(_07105_));
 OA211x2_ASAP7_75t_R _14073_ (.A1(_09595_),
    .A2(_06888_),
    .B(_07024_),
    .C(_06851_),
    .Y(_07106_));
 AO221x2_ASAP7_75t_R _14074_ (.A1(_04566_),
    .A2(_04581_),
    .B1(_06765_),
    .B2(_06767_),
    .C(_04608_),
    .Y(_07107_));
 OA211x2_ASAP7_75t_R _14075_ (.A1(_09590_),
    .A2(_06847_),
    .B(_07107_),
    .C(_06856_),
    .Y(_07108_));
 OR3x1_ASAP7_75t_R _14076_ (.A(_06838_),
    .B(_07106_),
    .C(_07108_),
    .Y(_07109_));
 OA21x2_ASAP7_75t_R _14077_ (.A1(_07027_),
    .A2(_07105_),
    .B(_07109_),
    .Y(_07110_));
 NAND2x1_ASAP7_75t_R _14078_ (.A(_06833_),
    .B(_07110_),
    .Y(_07111_));
 BUFx4f_ASAP7_75t_R _14079_ (.A(_06673_),
    .Y(_07112_));
 AND3x4_ASAP7_75t_R _14080_ (.A(_05358_),
    .B(_03714_),
    .C(_06827_),
    .Y(_07113_));
 AO221x1_ASAP7_75t_R _14081_ (.A1(_06713_),
    .A2(_03774_),
    .B1(_03746_),
    .B2(_05032_),
    .C(_03295_),
    .Y(_07114_));
 OA21x2_ASAP7_75t_R _14082_ (.A1(_06898_),
    .A2(_03554_),
    .B(_07114_),
    .Y(_07115_));
 AND4x1_ASAP7_75t_R _14083_ (.A(_07112_),
    .B(_07044_),
    .C(_07113_),
    .D(_07115_),
    .Y(_07116_));
 AO21x1_ASAP7_75t_R _14084_ (.A1(_07029_),
    .A2(_07028_),
    .B(_03555_),
    .Y(_07117_));
 BUFx3_ASAP7_75t_R _14085_ (.A(_03295_),
    .Y(_07118_));
 OR3x1_ASAP7_75t_R _14086_ (.A(_07118_),
    .B(_09565_),
    .C(_06894_),
    .Y(_07119_));
 AND4x1_ASAP7_75t_R _14087_ (.A(_06868_),
    .B(_07049_),
    .C(_07117_),
    .D(_07119_),
    .Y(_07120_));
 OA211x2_ASAP7_75t_R _14088_ (.A1(_09575_),
    .A2(_06896_),
    .B(_07039_),
    .C(_06861_),
    .Y(_07121_));
 OR4x2_ASAP7_75t_R _14089_ (.A(_03864_),
    .B(_03890_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07122_));
 OA211x2_ASAP7_75t_R _14090_ (.A1(_09580_),
    .A2(_06894_),
    .B(_07122_),
    .C(_07118_),
    .Y(_07123_));
 OA211x2_ASAP7_75t_R _14091_ (.A1(_07121_),
    .A2(_07123_),
    .B(_07022_),
    .C(_06832_),
    .Y(_07124_));
 OR3x1_ASAP7_75t_R _14092_ (.A(_07116_),
    .B(_07120_),
    .C(_07124_),
    .Y(_07125_));
 NOR2x1_ASAP7_75t_R _14093_ (.A(_06882_),
    .B(_07125_),
    .Y(_07126_));
 AO21x1_ASAP7_75t_R _14094_ (.A1(_06882_),
    .A2(_07111_),
    .B(_07126_),
    .Y(_07127_));
 NAND2x2_ASAP7_75t_R _14095_ (.A(_09652_),
    .B(_06769_),
    .Y(_07128_));
 OR2x2_ASAP7_75t_R _14096_ (.A(_09660_),
    .B(_06869_),
    .Y(_07129_));
 OA211x2_ASAP7_75t_R _14097_ (.A1(_09665_),
    .A2(_07066_),
    .B(_07083_),
    .C(_06883_),
    .Y(_07130_));
 AO31x2_ASAP7_75t_R _14098_ (.A1(_03297_),
    .A2(_07128_),
    .A3(_07129_),
    .B(_07130_),
    .Y(_07131_));
 NAND2x1_ASAP7_75t_R _14099_ (.A(_07043_),
    .B(_07131_),
    .Y(_07132_));
 OR4x2_ASAP7_75t_R _14100_ (.A(_06853_),
    .B(_06854_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07133_));
 OA31x2_ASAP7_75t_R _14101_ (.A1(_05442_),
    .A2(_05465_),
    .A3(_06769_),
    .B1(_07133_),
    .Y(_07134_));
 OA211x2_ASAP7_75t_R _14102_ (.A1(_09645_),
    .A2(_07066_),
    .B(_07079_),
    .C(_07029_),
    .Y(_07135_));
 AO21x1_ASAP7_75t_R _14103_ (.A1(_03297_),
    .A2(_07134_),
    .B(_07135_),
    .Y(_07136_));
 NAND2x1_ASAP7_75t_R _14104_ (.A(_06675_),
    .B(_07136_),
    .Y(_07137_));
 AO21x1_ASAP7_75t_R _14105_ (.A1(_07132_),
    .A2(_07137_),
    .B(_07056_),
    .Y(_07138_));
 OR3x1_ASAP7_75t_R _14106_ (.A(_03296_),
    .B(_07070_),
    .C(_07071_),
    .Y(_07139_));
 OA211x2_ASAP7_75t_R _14107_ (.A1(_07048_),
    .A2(_09690_),
    .B(_06770_),
    .C(_07139_),
    .Y(_07140_));
 AO21x1_ASAP7_75t_R _14108_ (.A1(_07062_),
    .A2(_06885_),
    .B(_07140_),
    .Y(_07141_));
 OR4x1_ASAP7_75t_R _14109_ (.A(_03427_),
    .B(_03496_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07142_));
 OA211x2_ASAP7_75t_R _14110_ (.A1(_09705_),
    .A2(_06769_),
    .B(_07142_),
    .C(_06851_),
    .Y(_07143_));
 OR3x1_ASAP7_75t_R _14111_ (.A(_07076_),
    .B(_06886_),
    .C(_07143_),
    .Y(_07144_));
 OA211x2_ASAP7_75t_R _14112_ (.A1(_06893_),
    .A2(_07141_),
    .B(_07144_),
    .C(_06891_),
    .Y(_07145_));
 OR4x2_ASAP7_75t_R _14113_ (.A(_06030_),
    .B(_06050_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07146_));
 OA211x2_ASAP7_75t_R _14114_ (.A1(_09680_),
    .A2(_06770_),
    .B(_07146_),
    .C(_06902_),
    .Y(_07147_));
 AO221x1_ASAP7_75t_R _14115_ (.A1(_06713_),
    .A2(_06301_),
    .B1(_06765_),
    .B2(_06767_),
    .C(_06321_),
    .Y(_07148_));
 OA211x2_ASAP7_75t_R _14116_ (.A1(_09675_),
    .A2(_07044_),
    .B(_07148_),
    .C(_07063_),
    .Y(_07149_));
 BUFx4f_ASAP7_75t_R _14117_ (.A(_07112_),
    .Y(_07150_));
 AND2x2_ASAP7_75t_R _14118_ (.A(_07150_),
    .B(_07076_),
    .Y(_07151_));
 OA21x2_ASAP7_75t_R _14119_ (.A1(_07147_),
    .A2(_07149_),
    .B(_07151_),
    .Y(_07152_));
 OAI21x1_ASAP7_75t_R _14120_ (.A1(_07145_),
    .A2(_07152_),
    .B(_06882_),
    .Y(_07153_));
 OA211x2_ASAP7_75t_R _14121_ (.A1(_06882_),
    .A2(_07138_),
    .B(_07153_),
    .C(_07088_),
    .Y(_07154_));
 AOI21x1_ASAP7_75t_R _14122_ (.A1(_07021_),
    .A2(_07127_),
    .B(_07154_),
    .Y(_07155_));
 BUFx4f_ASAP7_75t_R _14123_ (.A(_07004_),
    .Y(_07156_));
 AO21x1_ASAP7_75t_R _14124_ (.A1(_01158_),
    .A2(_07156_),
    .B(_07005_),
    .Y(_07157_));
 OAI21x1_ASAP7_75t_R _14125_ (.A1(_01158_),
    .A2(_07009_),
    .B(net164),
    .Y(_07158_));
 OA21x2_ASAP7_75t_R _14126_ (.A1(net163),
    .A2(_07157_),
    .B(_07158_),
    .Y(_07159_));
 BUFx3_ASAP7_75t_R _14127_ (.A(_07012_),
    .Y(_07160_));
 BUFx3_ASAP7_75t_R _14128_ (.A(_07014_),
    .Y(_07161_));
 INVx1_ASAP7_75t_R _14129_ (.A(_01212_),
    .Y(_07162_));
 AO22x1_ASAP7_75t_R _14130_ (.A1(_01213_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07162_),
    .Y(_07163_));
 AND2x2_ASAP7_75t_R _14131_ (.A(_07091_),
    .B(_07163_),
    .Y(_07164_));
 OR3x1_ASAP7_75t_R _14132_ (.A(_06831_),
    .B(_07159_),
    .C(_07164_),
    .Y(_07165_));
 OA21x2_ASAP7_75t_R _14133_ (.A1(_07019_),
    .A2(_07155_),
    .B(_07165_),
    .Y(net54));
 AO22x1_ASAP7_75t_R _14134_ (.A1(_01211_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_06949_),
    .Y(_07166_));
 INVx1_ASAP7_75t_R _14135_ (.A(net163),
    .Y(_07167_));
 AOI21x1_ASAP7_75t_R _14136_ (.A1(_03259_),
    .A2(_06897_),
    .B(_01215_),
    .Y(_07168_));
 AO21x1_ASAP7_75t_R _14137_ (.A1(_06824_),
    .A2(_07168_),
    .B(_07098_),
    .Y(_07169_));
 AO21x1_ASAP7_75t_R _14138_ (.A1(_07167_),
    .A2(_07169_),
    .B(_07162_),
    .Y(_07170_));
 OR3x1_ASAP7_75t_R _14139_ (.A(_03257_),
    .B(_06941_),
    .C(_07000_),
    .Y(_07171_));
 BUFx6f_ASAP7_75t_R _14140_ (.A(_07171_),
    .Y(_07172_));
 OAI21x1_ASAP7_75t_R _14141_ (.A1(_07009_),
    .A2(_07170_),
    .B(_07172_),
    .Y(_07173_));
 AND3x1_ASAP7_75t_R _14142_ (.A(_00998_),
    .B(_07156_),
    .C(_07170_),
    .Y(_07174_));
 AO221x1_ASAP7_75t_R _14143_ (.A1(_07091_),
    .A2(_07166_),
    .B1(_07173_),
    .B2(_06947_),
    .C(_07174_),
    .Y(_07175_));
 OA211x2_ASAP7_75t_R _14144_ (.A1(_09605_),
    .A2(_06862_),
    .B(_06844_),
    .C(_03295_),
    .Y(_07176_));
 AO31x2_ASAP7_75t_R _14145_ (.A1(_06883_),
    .A2(_07102_),
    .A3(_07103_),
    .B(_07176_),
    .Y(_07177_));
 OA211x2_ASAP7_75t_R _14146_ (.A1(_09590_),
    .A2(_06862_),
    .B(_07107_),
    .C(_06897_),
    .Y(_07178_));
 OA211x2_ASAP7_75t_R _14147_ (.A1(_09595_),
    .A2(_06769_),
    .B(_06872_),
    .C(_06856_),
    .Y(_07179_));
 OR3x1_ASAP7_75t_R _14148_ (.A(_06838_),
    .B(_07178_),
    .C(_07179_),
    .Y(_07180_));
 OA21x2_ASAP7_75t_R _14149_ (.A1(_07112_),
    .A2(_07177_),
    .B(_07180_),
    .Y(_07181_));
 AND2x2_ASAP7_75t_R _14150_ (.A(_06880_),
    .B(_07076_),
    .Y(_07182_));
 OA211x2_ASAP7_75t_R _14151_ (.A1(_09580_),
    .A2(_06869_),
    .B(_07122_),
    .C(_06897_),
    .Y(_07183_));
 AO31x2_ASAP7_75t_R _14152_ (.A1(_03296_),
    .A2(_06863_),
    .A3(_06864_),
    .B(_07183_),
    .Y(_07184_));
 AO21x1_ASAP7_75t_R _14153_ (.A1(_07063_),
    .A2(_07061_),
    .B(_07049_),
    .Y(_07185_));
 AO21x1_ASAP7_75t_R _14154_ (.A1(_03555_),
    .A2(_07185_),
    .B(_06839_),
    .Y(_07186_));
 OA211x2_ASAP7_75t_R _14155_ (.A1(_07150_),
    .A2(_07184_),
    .B(_07186_),
    .C(_06919_),
    .Y(_07187_));
 AO21x1_ASAP7_75t_R _14156_ (.A1(_07181_),
    .A2(_07182_),
    .B(_07187_),
    .Y(_07188_));
 OR2x2_ASAP7_75t_R _14157_ (.A(_07088_),
    .B(_07188_),
    .Y(_07189_));
 BUFx4f_ASAP7_75t_R _14158_ (.A(_06836_),
    .Y(_07190_));
 OA21x2_ASAP7_75t_R _14159_ (.A1(_09680_),
    .A2(_06770_),
    .B(_07146_),
    .Y(_07191_));
 NAND2x1_ASAP7_75t_R _14160_ (.A(_09667_),
    .B(_07066_),
    .Y(_07192_));
 AND3x1_ASAP7_75t_R _14161_ (.A(_06902_),
    .B(_07192_),
    .C(_06913_),
    .Y(_07193_));
 AO21x1_ASAP7_75t_R _14162_ (.A1(_07048_),
    .A2(_07191_),
    .B(_07193_),
    .Y(_07194_));
 OR4x1_ASAP7_75t_R _14163_ (.A(_06870_),
    .B(_06871_),
    .C(_06797_),
    .D(_06821_),
    .Y(_07195_));
 OA21x2_ASAP7_75t_R _14164_ (.A1(_09700_),
    .A2(_06894_),
    .B(_07195_),
    .Y(_07196_));
 OA211x2_ASAP7_75t_R _14165_ (.A1(_09705_),
    .A2(_06769_),
    .B(_07142_),
    .C(_06840_),
    .Y(_07197_));
 AO21x2_ASAP7_75t_R _14166_ (.A1(_07063_),
    .A2(_07196_),
    .B(_07197_),
    .Y(_07198_));
 OA211x2_ASAP7_75t_R _14167_ (.A1(_07118_),
    .A2(_09700_),
    .B(_06896_),
    .C(_07072_),
    .Y(_07199_));
 OA211x2_ASAP7_75t_R _14168_ (.A1(_06898_),
    .A2(_09685_),
    .B(_06894_),
    .C(_07064_),
    .Y(_07200_));
 OR3x1_ASAP7_75t_R _14169_ (.A(_06892_),
    .B(_07199_),
    .C(_07200_),
    .Y(_07201_));
 OA211x2_ASAP7_75t_R _14170_ (.A1(_07076_),
    .A2(_07198_),
    .B(_07201_),
    .C(_06860_),
    .Y(_07202_));
 AO21x1_ASAP7_75t_R _14171_ (.A1(_07151_),
    .A2(_07194_),
    .B(_07202_),
    .Y(_07203_));
 OA211x2_ASAP7_75t_R _14172_ (.A1(_09645_),
    .A2(_06862_),
    .B(_06910_),
    .C(_06856_),
    .Y(_07204_));
 AO31x2_ASAP7_75t_R _14173_ (.A1(_06883_),
    .A2(_07128_),
    .A3(_07129_),
    .B(_07204_),
    .Y(_07205_));
 OA211x2_ASAP7_75t_R _14174_ (.A1(_09625_),
    .A2(_06847_),
    .B(_06850_),
    .C(_06856_),
    .Y(_07206_));
 AO211x2_ASAP7_75t_R _14175_ (.A1(_06883_),
    .A2(_07134_),
    .B(_07206_),
    .C(_06838_),
    .Y(_07207_));
 OA21x2_ASAP7_75t_R _14176_ (.A1(_07112_),
    .A2(_07205_),
    .B(_07207_),
    .Y(_07208_));
 AO221x1_ASAP7_75t_R _14177_ (.A1(_07190_),
    .A2(_07203_),
    .B1(_07208_),
    .B2(_06919_),
    .C(_06921_),
    .Y(_07209_));
 AO21x1_ASAP7_75t_R _14178_ (.A1(_07189_),
    .A2(_07209_),
    .B(_06925_),
    .Y(_07210_));
 OA21x2_ASAP7_75t_R _14179_ (.A1(_06831_),
    .A2(_07175_),
    .B(_07210_),
    .Y(net57));
 AO21x1_ASAP7_75t_R _14180_ (.A1(_09705_),
    .A2(_06894_),
    .B(_06900_),
    .Y(_07211_));
 OA211x2_ASAP7_75t_R _14181_ (.A1(_09700_),
    .A2(_06769_),
    .B(_07195_),
    .C(_06840_),
    .Y(_07212_));
 AO21x1_ASAP7_75t_R _14182_ (.A1(_07063_),
    .A2(_07211_),
    .B(_07212_),
    .Y(_07213_));
 AND2x2_ASAP7_75t_R _14183_ (.A(_06868_),
    .B(_06889_),
    .Y(_07214_));
 AO21x1_ASAP7_75t_R _14184_ (.A1(_07042_),
    .A2(_07213_),
    .B(_07214_),
    .Y(_07215_));
 NAND2x1_ASAP7_75t_R _14185_ (.A(_06839_),
    .B(_06903_),
    .Y(_07216_));
 OR3x1_ASAP7_75t_R _14186_ (.A(_07022_),
    .B(_06914_),
    .C(_06916_),
    .Y(_07217_));
 AO21x1_ASAP7_75t_R _14187_ (.A1(_07216_),
    .A2(_07217_),
    .B(_06892_),
    .Y(_07218_));
 OA21x2_ASAP7_75t_R _14188_ (.A1(_06833_),
    .A2(_07215_),
    .B(_07218_),
    .Y(_07219_));
 OR3x1_ASAP7_75t_R _14189_ (.A(_07022_),
    .B(_06852_),
    .C(_06857_),
    .Y(_07220_));
 OA21x2_ASAP7_75t_R _14190_ (.A1(_06674_),
    .A2(_06912_),
    .B(_07220_),
    .Y(_07221_));
 AO22x1_ASAP7_75t_R _14191_ (.A1(_06881_),
    .A2(_07219_),
    .B1(_07221_),
    .B2(_06919_),
    .Y(_07222_));
 NAND2x1_ASAP7_75t_R _14192_ (.A(_06471_),
    .B(_06830_),
    .Y(_07223_));
 OA21x2_ASAP7_75t_R _14193_ (.A1(_06950_),
    .A2(_07008_),
    .B(_07172_),
    .Y(_07224_));
 NOR2x1_ASAP7_75t_R _14194_ (.A(_00965_),
    .B(_07224_),
    .Y(_07225_));
 AO22x1_ASAP7_75t_R _14195_ (.A1(_01209_),
    .A2(_06999_),
    .B1(_07013_),
    .B2(_06951_),
    .Y(_07226_));
 AO32x1_ASAP7_75t_R _14196_ (.A1(_00965_),
    .A2(_06950_),
    .A3(_07004_),
    .B1(_07226_),
    .B2(_06939_),
    .Y(_07227_));
 OR3x1_ASAP7_75t_R _14197_ (.A(_06829_),
    .B(_07225_),
    .C(_07227_),
    .Y(_07228_));
 OR3x1_ASAP7_75t_R _14198_ (.A(_06837_),
    .B(_06873_),
    .C(_06875_),
    .Y(_07229_));
 OA21x2_ASAP7_75t_R _14199_ (.A1(_06673_),
    .A2(_06846_),
    .B(_07229_),
    .Y(_07230_));
 AND2x2_ASAP7_75t_R _14200_ (.A(_06576_),
    .B(_06837_),
    .Y(_07231_));
 AO22x1_ASAP7_75t_R _14201_ (.A1(_06835_),
    .A2(_07230_),
    .B1(_07231_),
    .B2(_06867_),
    .Y(_07232_));
 OA21x2_ASAP7_75t_R _14202_ (.A1(_03554_),
    .A2(_06837_),
    .B(_06575_),
    .Y(_07233_));
 OA21x2_ASAP7_75t_R _14203_ (.A1(_06673_),
    .A2(_06867_),
    .B(_07233_),
    .Y(_07234_));
 AO21x1_ASAP7_75t_R _14204_ (.A1(_06835_),
    .A2(_07230_),
    .B(_07234_),
    .Y(_07235_));
 BUFx3_ASAP7_75t_R _14205_ (.A(_07049_),
    .Y(_07236_));
 AO32x1_ASAP7_75t_R _14206_ (.A1(_03714_),
    .A2(_07076_),
    .A3(_07232_),
    .B1(_07235_),
    .B2(_07236_),
    .Y(_07237_));
 OR3x1_ASAP7_75t_R _14207_ (.A(_06470_),
    .B(_06924_),
    .C(_07237_),
    .Y(_07238_));
 OA211x2_ASAP7_75t_R _14208_ (.A1(_07222_),
    .A2(_07223_),
    .B(_07228_),
    .C(_07238_),
    .Y(_07239_));
 BUFx12f_ASAP7_75t_R _14209_ (.A(_07239_),
    .Y(net58));
 BUFx4f_ASAP7_75t_R _14210_ (.A(_07004_),
    .Y(_07240_));
 AND3x1_ASAP7_75t_R _14211_ (.A(_01214_),
    .B(_01212_),
    .C(_01210_),
    .Y(_07241_));
 INVx1_ASAP7_75t_R _14212_ (.A(_07241_),
    .Y(_07242_));
 AOI21x1_ASAP7_75t_R _14213_ (.A1(_06824_),
    .A2(_07168_),
    .B(_07242_),
    .Y(_07243_));
 AO21x1_ASAP7_75t_R _14214_ (.A1(net164),
    .A2(_01212_),
    .B(_00998_),
    .Y(_07244_));
 AND2x2_ASAP7_75t_R _14215_ (.A(_01210_),
    .B(_07244_),
    .Y(_07245_));
 OA31x2_ASAP7_75t_R _14216_ (.A1(_00965_),
    .A2(_07243_),
    .A3(_07245_),
    .B1(_01208_),
    .Y(_07246_));
 XNOR2x1_ASAP7_75t_R _14217_ (.B(_07246_),
    .Y(_07247_),
    .A(_06945_));
 AO22x1_ASAP7_75t_R _14218_ (.A1(_01207_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_06953_),
    .Y(_07248_));
 BUFx4f_ASAP7_75t_R _14219_ (.A(_06940_),
    .Y(_07249_));
 AO222x2_ASAP7_75t_R _14220_ (.A1(_06945_),
    .A2(_07093_),
    .B1(_07240_),
    .B2(_07247_),
    .C1(_07248_),
    .C2(_07249_),
    .Y(_07250_));
 AND2x2_ASAP7_75t_R _14221_ (.A(_09700_),
    .B(_07066_),
    .Y(_07251_));
 AO21x1_ASAP7_75t_R _14222_ (.A1(_09690_),
    .A2(_07028_),
    .B(_03296_),
    .Y(_07252_));
 AO211x2_ASAP7_75t_R _14223_ (.A1(_09705_),
    .A2(_06894_),
    .B(_06900_),
    .C(_06898_),
    .Y(_07253_));
 OA211x2_ASAP7_75t_R _14224_ (.A1(_07251_),
    .A2(_07252_),
    .B(_07022_),
    .C(_07253_),
    .Y(_07254_));
 AND3x1_ASAP7_75t_R _14225_ (.A(_07112_),
    .B(_07044_),
    .C(_07059_),
    .Y(_07255_));
 OA21x2_ASAP7_75t_R _14226_ (.A1(_07254_),
    .A2(_07255_),
    .B(_06892_),
    .Y(_07256_));
 OR3x1_ASAP7_75t_R _14227_ (.A(_07042_),
    .B(_07082_),
    .C(_07084_),
    .Y(_07257_));
 OA211x2_ASAP7_75t_R _14228_ (.A1(_07150_),
    .A2(_07069_),
    .B(_07257_),
    .C(_06833_),
    .Y(_07258_));
 OA21x2_ASAP7_75t_R _14229_ (.A1(_07256_),
    .A2(_07258_),
    .B(_07190_),
    .Y(_07259_));
 OR3x1_ASAP7_75t_R _14230_ (.A(_07042_),
    .B(_07030_),
    .C(_07032_),
    .Y(_07260_));
 OA211x2_ASAP7_75t_R _14231_ (.A1(_07150_),
    .A2(_07081_),
    .B(_07260_),
    .C(_07076_),
    .Y(_07261_));
 AND2x2_ASAP7_75t_R _14232_ (.A(_07037_),
    .B(_07261_),
    .Y(_07262_));
 OR3x1_ASAP7_75t_R _14233_ (.A(_06921_),
    .B(_07259_),
    .C(_07262_),
    .Y(_07263_));
 OR3x1_ASAP7_75t_R _14234_ (.A(_06838_),
    .B(_07038_),
    .C(_07040_),
    .Y(_07264_));
 OA21x2_ASAP7_75t_R _14235_ (.A1(_07027_),
    .A2(_07026_),
    .B(_07264_),
    .Y(_07265_));
 OA211x2_ASAP7_75t_R _14236_ (.A1(_03555_),
    .A2(_07061_),
    .B(_06865_),
    .C(_06883_),
    .Y(_07266_));
 AND3x1_ASAP7_75t_R _14237_ (.A(_06902_),
    .B(_09565_),
    .C(_07044_),
    .Y(_07267_));
 OA21x2_ASAP7_75t_R _14238_ (.A1(_07266_),
    .A2(_07267_),
    .B(_06860_),
    .Y(_07268_));
 AND3x1_ASAP7_75t_R _14239_ (.A(_03714_),
    .B(_07036_),
    .C(_07268_),
    .Y(_07269_));
 AO21x1_ASAP7_75t_R _14240_ (.A1(_06881_),
    .A2(_07265_),
    .B(_07269_),
    .Y(_07270_));
 BUFx4f_ASAP7_75t_R _14241_ (.A(_06576_),
    .Y(_07271_));
 OA21x2_ASAP7_75t_R _14242_ (.A1(_06868_),
    .A2(_06770_),
    .B(_03555_),
    .Y(_07272_));
 AO21x1_ASAP7_75t_R _14243_ (.A1(_07046_),
    .A2(_07057_),
    .B(_07272_),
    .Y(_07273_));
 AND2x2_ASAP7_75t_R _14244_ (.A(_07271_),
    .B(_07273_),
    .Y(_07274_));
 AO221x1_ASAP7_75t_R _14245_ (.A1(_07054_),
    .A2(_07270_),
    .B1(_07274_),
    .B2(_07236_),
    .C(_07088_),
    .Y(_07275_));
 AO21x1_ASAP7_75t_R _14246_ (.A1(_07263_),
    .A2(_07275_),
    .B(_07019_),
    .Y(_07276_));
 OA21x2_ASAP7_75t_R _14247_ (.A1(_06831_),
    .A2(_07250_),
    .B(_07276_),
    .Y(net59));
 INVx1_ASAP7_75t_R _14248_ (.A(_01205_),
    .Y(_07277_));
 AO22x1_ASAP7_75t_R _14249_ (.A1(_01206_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07277_),
    .Y(_07278_));
 AO21x1_ASAP7_75t_R _14250_ (.A1(_06954_),
    .A2(_07156_),
    .B(_07005_),
    .Y(_07279_));
 BUFx6f_ASAP7_75t_R _14251_ (.A(_07008_),
    .Y(_07280_));
 OAI21x1_ASAP7_75t_R _14252_ (.A1(_06954_),
    .A2(_07280_),
    .B(_00898_),
    .Y(_07281_));
 OA21x2_ASAP7_75t_R _14253_ (.A1(_00898_),
    .A2(_07279_),
    .B(_07281_),
    .Y(_07282_));
 AOI21x1_ASAP7_75t_R _14254_ (.A1(_07249_),
    .A2(_07278_),
    .B(_07282_),
    .Y(_07283_));
 OR3x1_ASAP7_75t_R _14255_ (.A(_06674_),
    .B(_07147_),
    .C(_07149_),
    .Y(_07284_));
 OA21x2_ASAP7_75t_R _14256_ (.A1(_07043_),
    .A2(_07131_),
    .B(_07284_),
    .Y(_07285_));
 OR4x1_ASAP7_75t_R _14257_ (.A(_07070_),
    .B(_07071_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07286_));
 AND3x1_ASAP7_75t_R _14258_ (.A(_06861_),
    .B(_07148_),
    .C(_07286_),
    .Y(_07287_));
 AO211x2_ASAP7_75t_R _14259_ (.A1(_06848_),
    .A2(_06849_),
    .B(_06392_),
    .C(_06417_),
    .Y(_07288_));
 OA211x2_ASAP7_75t_R _14260_ (.A1(_09700_),
    .A2(_06847_),
    .B(_07288_),
    .C(_06856_),
    .Y(_07289_));
 OR3x1_ASAP7_75t_R _14261_ (.A(_06673_),
    .B(_07287_),
    .C(_07289_),
    .Y(_07290_));
 OR3x1_ASAP7_75t_R _14262_ (.A(_06838_),
    .B(_06886_),
    .C(_07143_),
    .Y(_07291_));
 AND2x2_ASAP7_75t_R _14263_ (.A(_07290_),
    .B(_07291_),
    .Y(_07292_));
 AND2x4_ASAP7_75t_R _14264_ (.A(_06469_),
    .B(_06892_),
    .Y(_07293_));
 INVx1_ASAP7_75t_R _14265_ (.A(_07293_),
    .Y(_07294_));
 OAI22x1_ASAP7_75t_R _14266_ (.A1(_07056_),
    .A2(_07285_),
    .B1(_07292_),
    .B2(_07294_),
    .Y(_07295_));
 NOR2x1_ASAP7_75t_R _14267_ (.A(_07150_),
    .B(_07136_),
    .Y(_07296_));
 NOR2x1_ASAP7_75t_R _14268_ (.A(_07023_),
    .B(_07105_),
    .Y(_07297_));
 OR4x1_ASAP7_75t_R _14269_ (.A(_06836_),
    .B(_06893_),
    .C(_07296_),
    .D(_07297_),
    .Y(_07298_));
 OA21x2_ASAP7_75t_R _14270_ (.A1(_06578_),
    .A2(_07295_),
    .B(_07298_),
    .Y(_07299_));
 OR3x2_ASAP7_75t_R _14271_ (.A(_07112_),
    .B(_07106_),
    .C(_07108_),
    .Y(_07300_));
 OR3x2_ASAP7_75t_R _14272_ (.A(_07022_),
    .B(_07121_),
    .C(_07123_),
    .Y(_07301_));
 AND3x1_ASAP7_75t_R _14273_ (.A(_06880_),
    .B(_07300_),
    .C(_07301_),
    .Y(_07302_));
 AND3x1_ASAP7_75t_R _14274_ (.A(_07036_),
    .B(_07057_),
    .C(_07115_),
    .Y(_07303_));
 OA21x2_ASAP7_75t_R _14275_ (.A1(_07302_),
    .A2(_07303_),
    .B(_07113_),
    .Y(_07304_));
 AO21x1_ASAP7_75t_R _14276_ (.A1(_07057_),
    .A2(_07115_),
    .B(_07272_),
    .Y(_07305_));
 AND2x2_ASAP7_75t_R _14277_ (.A(_07036_),
    .B(_07305_),
    .Y(_07306_));
 OA21x2_ASAP7_75t_R _14278_ (.A1(_07302_),
    .A2(_07306_),
    .B(_07236_),
    .Y(_07307_));
 OAI21x1_ASAP7_75t_R _14279_ (.A1(_07304_),
    .A2(_07307_),
    .B(_06921_),
    .Y(_07308_));
 OA211x2_ASAP7_75t_R _14280_ (.A1(_07021_),
    .A2(_07299_),
    .B(_07308_),
    .C(_06830_),
    .Y(_07309_));
 AOI21x1_ASAP7_75t_R _14281_ (.A1(_07019_),
    .A2(_07283_),
    .B(_07309_),
    .Y(net60));
 AO21x1_ASAP7_75t_R _14282_ (.A1(_07063_),
    .A2(_07134_),
    .B(_07206_),
    .Y(_07310_));
 OR2x2_ASAP7_75t_R _14283_ (.A(_07027_),
    .B(_07310_),
    .Y(_07311_));
 OR2x2_ASAP7_75t_R _14284_ (.A(_06839_),
    .B(_07177_),
    .Y(_07312_));
 OR4x1_ASAP7_75t_R _14285_ (.A(_06392_),
    .B(_06417_),
    .C(_06870_),
    .D(_06871_),
    .Y(_07313_));
 OA211x2_ASAP7_75t_R _14286_ (.A1(_09680_),
    .A2(_06869_),
    .B(_07313_),
    .C(_06897_),
    .Y(_07314_));
 AND3x1_ASAP7_75t_R _14287_ (.A(_03295_),
    .B(_07148_),
    .C(_07286_),
    .Y(_07315_));
 OR3x1_ASAP7_75t_R _14288_ (.A(_07027_),
    .B(_07314_),
    .C(_07315_),
    .Y(_07316_));
 OA21x2_ASAP7_75t_R _14289_ (.A1(_07023_),
    .A2(_07198_),
    .B(_07316_),
    .Y(_07317_));
 OR2x2_ASAP7_75t_R _14290_ (.A(_06839_),
    .B(_07205_),
    .Y(_07318_));
 OA211x2_ASAP7_75t_R _14291_ (.A1(_07150_),
    .A2(_07194_),
    .B(_07318_),
    .C(_06833_),
    .Y(_07319_));
 AO21x1_ASAP7_75t_R _14292_ (.A1(_07056_),
    .A2(_07317_),
    .B(_07319_),
    .Y(_07320_));
 AO32x1_ASAP7_75t_R _14293_ (.A1(_06919_),
    .A2(_07311_),
    .A3(_07312_),
    .B1(_07320_),
    .B2(_06882_),
    .Y(_07321_));
 OR3x1_ASAP7_75t_R _14294_ (.A(_06868_),
    .B(_07178_),
    .C(_07179_),
    .Y(_07322_));
 OA21x2_ASAP7_75t_R _14295_ (.A1(_06860_),
    .A2(_07184_),
    .B(_07322_),
    .Y(_07323_));
 AND3x2_ASAP7_75t_R _14296_ (.A(_07029_),
    .B(_06837_),
    .C(_06896_),
    .Y(_07324_));
 OA211x2_ASAP7_75t_R _14297_ (.A1(_07236_),
    .A2(_07324_),
    .B(_09561_),
    .C(_07271_),
    .Y(_07325_));
 AO21x1_ASAP7_75t_R _14298_ (.A1(_07190_),
    .A2(_07323_),
    .B(_07325_),
    .Y(_07326_));
 AND2x2_ASAP7_75t_R _14299_ (.A(_06921_),
    .B(_07054_),
    .Y(_07327_));
 AO221x2_ASAP7_75t_R _14300_ (.A1(_06472_),
    .A2(_07321_),
    .B1(_07326_),
    .B2(_07327_),
    .C(_07019_),
    .Y(_07328_));
 OA21x2_ASAP7_75t_R _14301_ (.A1(_00932_),
    .A2(_07246_),
    .B(_00931_),
    .Y(_07329_));
 OA21x2_ASAP7_75t_R _14302_ (.A1(_00898_),
    .A2(_07329_),
    .B(_01205_),
    .Y(_07330_));
 AOI211x1_ASAP7_75t_R _14303_ (.A1(_07240_),
    .A2(_07330_),
    .B(_00865_),
    .C(_07093_),
    .Y(_07331_));
 OA21x2_ASAP7_75t_R _14304_ (.A1(_07280_),
    .A2(_07330_),
    .B(_00865_),
    .Y(_07332_));
 INVx1_ASAP7_75t_R _14305_ (.A(_00864_),
    .Y(_07333_));
 AO22x1_ASAP7_75t_R _14306_ (.A1(_01204_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07333_),
    .Y(_07334_));
 AOI21x1_ASAP7_75t_R _14307_ (.A1(_07091_),
    .A2(_07334_),
    .B(_06830_),
    .Y(_07335_));
 OAI21x1_ASAP7_75t_R _14308_ (.A1(_07331_),
    .A2(_07332_),
    .B(_07335_),
    .Y(_07336_));
 AND2x6_ASAP7_75t_R _14309_ (.A(_07328_),
    .B(_07336_),
    .Y(net61));
 OR2x2_ASAP7_75t_R _14310_ (.A(_07042_),
    .B(_07213_),
    .Y(_07337_));
 OA211x2_ASAP7_75t_R _14311_ (.A1(_09685_),
    .A2(_06896_),
    .B(_06913_),
    .C(_06898_),
    .Y(_07338_));
 OA211x2_ASAP7_75t_R _14312_ (.A1(_09680_),
    .A2(_06894_),
    .B(_07313_),
    .C(_07118_),
    .Y(_07339_));
 OR3x1_ASAP7_75t_R _14313_ (.A(_06674_),
    .B(_07338_),
    .C(_07339_),
    .Y(_07340_));
 AO32x1_ASAP7_75t_R _14314_ (.A1(_06836_),
    .A2(_07337_),
    .A3(_07340_),
    .B1(_06889_),
    .B2(_07231_),
    .Y(_07341_));
 AND2x2_ASAP7_75t_R _14315_ (.A(_06880_),
    .B(_06918_),
    .Y(_07342_));
 AND2x2_ASAP7_75t_R _14316_ (.A(_07036_),
    .B(_06859_),
    .Y(_07343_));
 OR3x1_ASAP7_75t_R _14317_ (.A(_07056_),
    .B(_07342_),
    .C(_07343_),
    .Y(_07344_));
 OA21x2_ASAP7_75t_R _14318_ (.A1(_07054_),
    .A2(_07341_),
    .B(_07344_),
    .Y(_07345_));
 OA21x2_ASAP7_75t_R _14319_ (.A1(_06860_),
    .A2(_06867_),
    .B(_06876_),
    .Y(_07346_));
 OR2x2_ASAP7_75t_R _14320_ (.A(_03555_),
    .B(_06834_),
    .Y(_07347_));
 AND2x4_ASAP7_75t_R _14321_ (.A(_06834_),
    .B(_07113_),
    .Y(_07348_));
 AO21x1_ASAP7_75t_R _14322_ (.A1(_07236_),
    .A2(_07347_),
    .B(_07348_),
    .Y(_07349_));
 OA21x2_ASAP7_75t_R _14323_ (.A1(_06577_),
    .A2(_07346_),
    .B(_07349_),
    .Y(_07350_));
 OR3x1_ASAP7_75t_R _14324_ (.A(_07088_),
    .B(_06924_),
    .C(_07350_),
    .Y(_07351_));
 OAI21x1_ASAP7_75t_R _14325_ (.A1(_00865_),
    .A2(_06955_),
    .B(_00864_),
    .Y(_07352_));
 OR3x1_ASAP7_75t_R _14326_ (.A(_06939_),
    .B(_07002_),
    .C(_07352_),
    .Y(_07353_));
 AOI21x1_ASAP7_75t_R _14327_ (.A1(_07172_),
    .A2(_07353_),
    .B(_00831_),
    .Y(_07354_));
 INVx1_ASAP7_75t_R _14328_ (.A(_01202_),
    .Y(_07355_));
 AO22x1_ASAP7_75t_R _14329_ (.A1(_01203_),
    .A2(_06999_),
    .B1(_07013_),
    .B2(_07355_),
    .Y(_07356_));
 AO32x1_ASAP7_75t_R _14330_ (.A1(_00831_),
    .A2(_07004_),
    .A3(_07352_),
    .B1(_07356_),
    .B2(_06939_),
    .Y(_07357_));
 OR3x1_ASAP7_75t_R _14331_ (.A(_06830_),
    .B(_07354_),
    .C(_07357_),
    .Y(_07358_));
 OA211x2_ASAP7_75t_R _14332_ (.A1(_07223_),
    .A2(_07345_),
    .B(_07351_),
    .C(_07358_),
    .Y(_07359_));
 BUFx12_ASAP7_75t_R _14333_ (.A(_07359_),
    .Y(net62));
 INVx1_ASAP7_75t_R _14334_ (.A(_00798_),
    .Y(_07360_));
 OR4x1_ASAP7_75t_R _14335_ (.A(_00831_),
    .B(_00865_),
    .C(_00898_),
    .D(_00932_),
    .Y(_07361_));
 OR3x1_ASAP7_75t_R _14336_ (.A(_00965_),
    .B(_07245_),
    .C(_07361_),
    .Y(_07362_));
 OR2x2_ASAP7_75t_R _14337_ (.A(_00898_),
    .B(_00931_),
    .Y(_07363_));
 AO21x1_ASAP7_75t_R _14338_ (.A1(_01205_),
    .A2(_07363_),
    .B(_00865_),
    .Y(_07364_));
 AO21x1_ASAP7_75t_R _14339_ (.A1(_00864_),
    .A2(_07364_),
    .B(_00831_),
    .Y(_07365_));
 OA211x2_ASAP7_75t_R _14340_ (.A1(_01208_),
    .A2(_07361_),
    .B(_07365_),
    .C(_01202_),
    .Y(_07366_));
 OA21x2_ASAP7_75t_R _14341_ (.A1(_07243_),
    .A2(_07362_),
    .B(_07366_),
    .Y(_07367_));
 AO21x1_ASAP7_75t_R _14342_ (.A1(_07240_),
    .A2(_07367_),
    .B(_07093_),
    .Y(_07368_));
 INVx1_ASAP7_75t_R _14343_ (.A(_00797_),
    .Y(_07369_));
 AO22x1_ASAP7_75t_R _14344_ (.A1(_01201_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07369_),
    .Y(_07370_));
 NOR2x1_ASAP7_75t_R _14345_ (.A(_07009_),
    .B(_07367_),
    .Y(_07371_));
 AO221x1_ASAP7_75t_R _14346_ (.A1(_06940_),
    .A2(_07370_),
    .B1(_07371_),
    .B2(_00798_),
    .C(_06830_),
    .Y(_07372_));
 AO21x2_ASAP7_75t_R _14347_ (.A1(_07360_),
    .A2(_07368_),
    .B(_07372_),
    .Y(_07373_));
 BUFx4f_ASAP7_75t_R _14348_ (.A(_06893_),
    .Y(_07374_));
 AND2x2_ASAP7_75t_R _14349_ (.A(_07271_),
    .B(_07034_),
    .Y(_07375_));
 AO21x1_ASAP7_75t_R _14350_ (.A1(_07190_),
    .A2(_07086_),
    .B(_07375_),
    .Y(_07376_));
 OA21x2_ASAP7_75t_R _14351_ (.A1(_09685_),
    .A2(_07061_),
    .B(_06913_),
    .Y(_07377_));
 OA211x2_ASAP7_75t_R _14352_ (.A1(_09680_),
    .A2(_07028_),
    .B(_06915_),
    .C(_06898_),
    .Y(_07378_));
 AO21x1_ASAP7_75t_R _14353_ (.A1(_06902_),
    .A2(_07377_),
    .B(_07378_),
    .Y(_07379_));
 OA211x2_ASAP7_75t_R _14354_ (.A1(_07251_),
    .A2(_07252_),
    .B(_07027_),
    .C(_07253_),
    .Y(_07380_));
 AOI21x1_ASAP7_75t_R _14355_ (.A1(_06891_),
    .A2(_07379_),
    .B(_07380_),
    .Y(_07381_));
 NAND2x1_ASAP7_75t_R _14356_ (.A(_06577_),
    .B(_07060_),
    .Y(_07382_));
 OA21x2_ASAP7_75t_R _14357_ (.A1(_07271_),
    .A2(_07381_),
    .B(_07382_),
    .Y(_07383_));
 NAND2x1_ASAP7_75t_R _14358_ (.A(_07374_),
    .B(_07383_),
    .Y(_07384_));
 OA211x2_ASAP7_75t_R _14359_ (.A1(_07374_),
    .A2(_07376_),
    .B(_07384_),
    .C(_07088_),
    .Y(_07385_));
 AO221x1_ASAP7_75t_R _14360_ (.A1(_07062_),
    .A2(_07046_),
    .B1(_07050_),
    .B2(_07048_),
    .C(_06860_),
    .Y(_07386_));
 OA31x2_ASAP7_75t_R _14361_ (.A1(_07023_),
    .A2(_07047_),
    .A3(_07050_),
    .B1(_07041_),
    .Y(_07387_));
 AO32x1_ASAP7_75t_R _14362_ (.A1(_07041_),
    .A2(_07113_),
    .A3(_07386_),
    .B1(_07387_),
    .B2(_07236_),
    .Y(_07388_));
 AND3x1_ASAP7_75t_R _14363_ (.A(_09561_),
    .B(_07036_),
    .C(_07236_),
    .Y(_07389_));
 AO21x1_ASAP7_75t_R _14364_ (.A1(_06882_),
    .A2(_07388_),
    .B(_07389_),
    .Y(_07390_));
 AND2x2_ASAP7_75t_R _14365_ (.A(_07021_),
    .B(_07390_),
    .Y(_07391_));
 OR3x2_ASAP7_75t_R _14366_ (.A(_07019_),
    .B(_07385_),
    .C(_07391_),
    .Y(_07392_));
 AND2x6_ASAP7_75t_R _14367_ (.A(_07373_),
    .B(_07392_),
    .Y(net63));
 INVx1_ASAP7_75t_R _14368_ (.A(_06956_),
    .Y(_07393_));
 OAI21x1_ASAP7_75t_R _14369_ (.A1(_06955_),
    .A2(_06957_),
    .B(_06960_),
    .Y(_07394_));
 OAI21x1_ASAP7_75t_R _14370_ (.A1(_07394_),
    .A2(_07280_),
    .B(_07172_),
    .Y(_07395_));
 INVx1_ASAP7_75t_R _14371_ (.A(_01199_),
    .Y(_07396_));
 AO22x1_ASAP7_75t_R _14372_ (.A1(_01200_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07396_),
    .Y(_07397_));
 AO32x1_ASAP7_75t_R _14373_ (.A1(_06956_),
    .A2(_07394_),
    .A3(_07156_),
    .B1(_07397_),
    .B2(_06940_),
    .Y(_07398_));
 AO21x1_ASAP7_75t_R _14374_ (.A1(_07393_),
    .A2(_07395_),
    .B(_07398_),
    .Y(_07399_));
 AO21x1_ASAP7_75t_R _14375_ (.A1(_06881_),
    .A2(_07125_),
    .B(_07389_),
    .Y(_07400_));
 NAND2x1_ASAP7_75t_R _14376_ (.A(_07021_),
    .B(_07400_),
    .Y(_07401_));
 NAND2x1_ASAP7_75t_R _14377_ (.A(_09667_),
    .B(_06888_),
    .Y(_07402_));
 OR2x2_ASAP7_75t_R _14378_ (.A(_09675_),
    .B(_06841_),
    .Y(_07403_));
 OA211x2_ASAP7_75t_R _14379_ (.A1(_09680_),
    .A2(_06847_),
    .B(_06915_),
    .C(_06856_),
    .Y(_07404_));
 AO31x2_ASAP7_75t_R _14380_ (.A1(_06883_),
    .A2(_07402_),
    .A3(_07403_),
    .B(_07404_),
    .Y(_07405_));
 OR3x1_ASAP7_75t_R _14381_ (.A(_06838_),
    .B(_07287_),
    .C(_07289_),
    .Y(_07406_));
 OA211x2_ASAP7_75t_R _14382_ (.A1(_07150_),
    .A2(_07405_),
    .B(_07406_),
    .C(_06892_),
    .Y(_07407_));
 NOR2x1_ASAP7_75t_R _14383_ (.A(_07037_),
    .B(_07407_),
    .Y(_07408_));
 OA211x2_ASAP7_75t_R _14384_ (.A1(_06886_),
    .A2(_07143_),
    .B(_07023_),
    .C(_06892_),
    .Y(_07409_));
 NOR2x1_ASAP7_75t_R _14385_ (.A(_07190_),
    .B(_07409_),
    .Y(_07410_));
 AO221x1_ASAP7_75t_R _14386_ (.A1(_07138_),
    .A2(_07408_),
    .B1(_07410_),
    .B2(_07111_),
    .C(_06921_),
    .Y(_07411_));
 AOI21x1_ASAP7_75t_R _14387_ (.A1(_07401_),
    .A2(_07411_),
    .B(_06925_),
    .Y(_07412_));
 AO21x2_ASAP7_75t_R _14388_ (.A1(_07019_),
    .A2(_07399_),
    .B(_07412_),
    .Y(net33));
 AND2x2_ASAP7_75t_R _14389_ (.A(_06576_),
    .B(_07181_),
    .Y(_07413_));
 AND2x2_ASAP7_75t_R _14390_ (.A(_06880_),
    .B(_07208_),
    .Y(_07414_));
 OA211x2_ASAP7_75t_R _14391_ (.A1(_09660_),
    .A2(_06869_),
    .B(_07146_),
    .C(_06897_),
    .Y(_07415_));
 AO31x2_ASAP7_75t_R _14392_ (.A1(_07118_),
    .A2(_07402_),
    .A3(_07403_),
    .B(_07415_),
    .Y(_07416_));
 OR3x1_ASAP7_75t_R _14393_ (.A(_06837_),
    .B(_07314_),
    .C(_07315_),
    .Y(_07417_));
 OA21x2_ASAP7_75t_R _14394_ (.A1(_06868_),
    .A2(_07416_),
    .B(_07417_),
    .Y(_07418_));
 AO221x1_ASAP7_75t_R _14395_ (.A1(_07198_),
    .A2(_07231_),
    .B1(_07418_),
    .B2(_06880_),
    .C(_07076_),
    .Y(_07419_));
 OA31x2_ASAP7_75t_R _14396_ (.A1(_06893_),
    .A2(_07413_),
    .A3(_07414_),
    .B1(_07419_),
    .Y(_07420_));
 AND4x1_ASAP7_75t_R _14397_ (.A(_07063_),
    .B(_03555_),
    .C(_06868_),
    .D(_07044_),
    .Y(_07421_));
 AO21x1_ASAP7_75t_R _14398_ (.A1(_07023_),
    .A2(_07184_),
    .B(_07421_),
    .Y(_07422_));
 NAND2x2_ASAP7_75t_R _14399_ (.A(_06835_),
    .B(_06839_),
    .Y(_07423_));
 AND3x1_ASAP7_75t_R _14400_ (.A(_06835_),
    .B(_06839_),
    .C(_07184_),
    .Y(_07424_));
 AO21x1_ASAP7_75t_R _14401_ (.A1(_09561_),
    .A2(_07423_),
    .B(_07424_),
    .Y(_07425_));
 AO221x1_ASAP7_75t_R _14402_ (.A1(_07348_),
    .A2(_07422_),
    .B1(_07425_),
    .B2(_07236_),
    .C(_06470_),
    .Y(_07426_));
 OA21x2_ASAP7_75t_R _14403_ (.A1(_06921_),
    .A2(_07420_),
    .B(_07426_),
    .Y(_07427_));
 AND2x2_ASAP7_75t_R _14404_ (.A(_01199_),
    .B(_06960_),
    .Y(_07428_));
 OA211x2_ASAP7_75t_R _14405_ (.A1(_06957_),
    .A2(_07330_),
    .B(_07428_),
    .C(_07004_),
    .Y(_07429_));
 AND3x1_ASAP7_75t_R _14406_ (.A(_06956_),
    .B(_01199_),
    .C(_07004_),
    .Y(_07430_));
 INVx1_ASAP7_75t_R _14407_ (.A(_01197_),
    .Y(_07431_));
 AO22x1_ASAP7_75t_R _14408_ (.A1(_01198_),
    .A2(_06999_),
    .B1(_07013_),
    .B2(_07431_),
    .Y(_07432_));
 AND2x2_ASAP7_75t_R _14409_ (.A(_06939_),
    .B(_07432_),
    .Y(_07433_));
 OR4x1_ASAP7_75t_R _14410_ (.A(_00731_),
    .B(_06829_),
    .C(_07001_),
    .D(_07433_),
    .Y(_07434_));
 OR3x1_ASAP7_75t_R _14411_ (.A(_07429_),
    .B(_07430_),
    .C(_07434_),
    .Y(_07435_));
 OAI21x1_ASAP7_75t_R _14412_ (.A1(_06957_),
    .A2(_07330_),
    .B(_07428_),
    .Y(_07436_));
 AOI21x1_ASAP7_75t_R _14413_ (.A1(_06956_),
    .A2(_01199_),
    .B(_07008_),
    .Y(_07437_));
 INVx1_ASAP7_75t_R _14414_ (.A(_00731_),
    .Y(_07438_));
 OR3x1_ASAP7_75t_R _14415_ (.A(_07438_),
    .B(_06829_),
    .C(_07433_),
    .Y(_07439_));
 AO21x1_ASAP7_75t_R _14416_ (.A1(_07436_),
    .A2(_07437_),
    .B(_07439_),
    .Y(_07440_));
 OA211x2_ASAP7_75t_R _14417_ (.A1(_06925_),
    .A2(_07427_),
    .B(_07435_),
    .C(_07440_),
    .Y(_07441_));
 BUFx10_ASAP7_75t_R _14418_ (.A(_07441_),
    .Y(net34));
 OA211x2_ASAP7_75t_R _14419_ (.A1(_09665_),
    .A2(_06896_),
    .B(_06910_),
    .C(_06898_),
    .Y(_07442_));
 OA211x2_ASAP7_75t_R _14420_ (.A1(_09660_),
    .A2(_06894_),
    .B(_07146_),
    .C(_07118_),
    .Y(_07443_));
 OA21x2_ASAP7_75t_R _14421_ (.A1(_07442_),
    .A2(_07443_),
    .B(_07022_),
    .Y(_07444_));
 OA21x2_ASAP7_75t_R _14422_ (.A1(_07338_),
    .A2(_07339_),
    .B(_07112_),
    .Y(_07445_));
 OR3x1_ASAP7_75t_R _14423_ (.A(_06576_),
    .B(_07444_),
    .C(_07445_),
    .Y(_07446_));
 OA211x2_ASAP7_75t_R _14424_ (.A1(_06881_),
    .A2(_07215_),
    .B(_07446_),
    .C(_06893_),
    .Y(_07447_));
 OR2x2_ASAP7_75t_R _14425_ (.A(_06577_),
    .B(_07221_),
    .Y(_07448_));
 OA211x2_ASAP7_75t_R _14426_ (.A1(_06882_),
    .A2(_07230_),
    .B(_07448_),
    .C(_07054_),
    .Y(_07449_));
 OA21x2_ASAP7_75t_R _14427_ (.A1(_07447_),
    .A2(_07449_),
    .B(_06472_),
    .Y(_07450_));
 AND2x2_ASAP7_75t_R _14428_ (.A(_03555_),
    .B(_07049_),
    .Y(_07451_));
 BUFx4f_ASAP7_75t_R _14429_ (.A(_07451_),
    .Y(_07452_));
 AND3x1_ASAP7_75t_R _14430_ (.A(_07190_),
    .B(_06891_),
    .C(_06867_),
    .Y(_07453_));
 AO21x1_ASAP7_75t_R _14431_ (.A1(_07452_),
    .A2(_07423_),
    .B(_07453_),
    .Y(_07454_));
 AO21x1_ASAP7_75t_R _14432_ (.A1(_07327_),
    .A2(_07454_),
    .B(_07019_),
    .Y(_07455_));
 BUFx4f_ASAP7_75t_R _14433_ (.A(_06830_),
    .Y(_07456_));
 OA21x2_ASAP7_75t_R _14434_ (.A1(_06955_),
    .A2(_06958_),
    .B(_06962_),
    .Y(_07457_));
 NAND2x1_ASAP7_75t_R _14435_ (.A(_01197_),
    .B(_07457_),
    .Y(_07458_));
 OA21x2_ASAP7_75t_R _14436_ (.A1(_07458_),
    .A2(_07009_),
    .B(_07172_),
    .Y(_07459_));
 NOR2x1_ASAP7_75t_R _14437_ (.A(_00698_),
    .B(_07459_),
    .Y(_07460_));
 BUFx3_ASAP7_75t_R _14438_ (.A(_07004_),
    .Y(_07461_));
 INVx1_ASAP7_75t_R _14439_ (.A(_01195_),
    .Y(_07462_));
 AO22x1_ASAP7_75t_R _14440_ (.A1(_01196_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07462_),
    .Y(_07463_));
 AO32x1_ASAP7_75t_R _14441_ (.A1(_00698_),
    .A2(_07458_),
    .A3(_07461_),
    .B1(_07463_),
    .B2(_06940_),
    .Y(_07464_));
 OR3x1_ASAP7_75t_R _14442_ (.A(_07456_),
    .B(_07460_),
    .C(_07464_),
    .Y(_07465_));
 OA21x2_ASAP7_75t_R _14443_ (.A1(_07450_),
    .A2(_07455_),
    .B(_07465_),
    .Y(net35));
 INVx1_ASAP7_75t_R _14444_ (.A(_00665_),
    .Y(_07466_));
 OR4x1_ASAP7_75t_R _14445_ (.A(_00698_),
    .B(_00731_),
    .C(_06956_),
    .D(_00798_),
    .Y(_07467_));
 OA21x2_ASAP7_75t_R _14446_ (.A1(_06956_),
    .A2(_00797_),
    .B(_01199_),
    .Y(_07468_));
 OA21x2_ASAP7_75t_R _14447_ (.A1(_00731_),
    .A2(_07468_),
    .B(_01197_),
    .Y(_07469_));
 OA21x2_ASAP7_75t_R _14448_ (.A1(_00698_),
    .A2(_07469_),
    .B(_01195_),
    .Y(_07470_));
 OA21x2_ASAP7_75t_R _14449_ (.A1(_07367_),
    .A2(_07467_),
    .B(_07470_),
    .Y(_07471_));
 AO21x1_ASAP7_75t_R _14450_ (.A1(_07240_),
    .A2(_07471_),
    .B(_07093_),
    .Y(_07472_));
 INVx1_ASAP7_75t_R _14451_ (.A(_07471_),
    .Y(_07473_));
 INVx1_ASAP7_75t_R _14452_ (.A(_01193_),
    .Y(_07474_));
 AO22x1_ASAP7_75t_R _14453_ (.A1(_01194_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07474_),
    .Y(_07475_));
 AO32x1_ASAP7_75t_R _14454_ (.A1(_00665_),
    .A2(_07461_),
    .A3(_07473_),
    .B1(_07475_),
    .B2(_06940_),
    .Y(_07476_));
 AO21x1_ASAP7_75t_R _14455_ (.A1(_07466_),
    .A2(_07472_),
    .B(_07476_),
    .Y(_07477_));
 AND2x2_ASAP7_75t_R _14456_ (.A(_07076_),
    .B(_07265_),
    .Y(_07478_));
 NOR2x1_ASAP7_75t_R _14457_ (.A(_07256_),
    .B(_07478_),
    .Y(_07479_));
 OA21x2_ASAP7_75t_R _14458_ (.A1(_09660_),
    .A2(_07044_),
    .B(_06907_),
    .Y(_07480_));
 AO21x1_ASAP7_75t_R _14459_ (.A1(_07192_),
    .A2(_06910_),
    .B(_07048_),
    .Y(_07481_));
 OAI21x1_ASAP7_75t_R _14460_ (.A1(_03297_),
    .A2(_07480_),
    .B(_07481_),
    .Y(_07482_));
 NOR2x1_ASAP7_75t_R _14461_ (.A(_07023_),
    .B(_07379_),
    .Y(_07483_));
 AOI21x1_ASAP7_75t_R _14462_ (.A1(_06891_),
    .A2(_07482_),
    .B(_07483_),
    .Y(_07484_));
 AOI211x1_ASAP7_75t_R _14463_ (.A1(_07374_),
    .A2(_07484_),
    .B(_07261_),
    .C(_07037_),
    .Y(_07485_));
 AOI21x1_ASAP7_75t_R _14464_ (.A1(_06578_),
    .A2(_07479_),
    .B(_07485_),
    .Y(_07486_));
 OR3x2_ASAP7_75t_R _14465_ (.A(_06576_),
    .B(_07027_),
    .C(_06770_),
    .Y(_07487_));
 AND4x1_ASAP7_75t_R _14466_ (.A(_06835_),
    .B(_07042_),
    .C(_07062_),
    .D(_07046_),
    .Y(_07488_));
 AO21x1_ASAP7_75t_R _14467_ (.A1(_09561_),
    .A2(_07487_),
    .B(_07488_),
    .Y(_07489_));
 AO221x1_ASAP7_75t_R _14468_ (.A1(_07268_),
    .A2(_07348_),
    .B1(_07489_),
    .B2(_07236_),
    .C(_06471_),
    .Y(_07490_));
 OA211x2_ASAP7_75t_R _14469_ (.A1(_07021_),
    .A2(_07486_),
    .B(_07490_),
    .C(_07456_),
    .Y(_07491_));
 AO21x2_ASAP7_75t_R _14470_ (.A1(_07019_),
    .A2(_07477_),
    .B(_07491_),
    .Y(net36));
 INVx1_ASAP7_75t_R _14471_ (.A(_00632_),
    .Y(_07492_));
 INVx1_ASAP7_75t_R _14472_ (.A(_00698_),
    .Y(_07493_));
 AOI21x1_ASAP7_75t_R _14473_ (.A1(_07493_),
    .A2(_07458_),
    .B(_07462_),
    .Y(_07494_));
 OAI21x1_ASAP7_75t_R _14474_ (.A1(_00665_),
    .A2(_07494_),
    .B(_01193_),
    .Y(_07495_));
 OAI21x1_ASAP7_75t_R _14475_ (.A1(_07280_),
    .A2(_07495_),
    .B(_07172_),
    .Y(_07496_));
 INVx1_ASAP7_75t_R _14476_ (.A(_01191_),
    .Y(_07497_));
 AO22x1_ASAP7_75t_R _14477_ (.A1(_01192_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07497_),
    .Y(_07498_));
 AO32x1_ASAP7_75t_R _14478_ (.A1(_00632_),
    .A2(_07461_),
    .A3(_07495_),
    .B1(_07498_),
    .B2(_07091_),
    .Y(_07499_));
 AOI21x1_ASAP7_75t_R _14479_ (.A1(_07492_),
    .A2(_07496_),
    .B(_07499_),
    .Y(_07500_));
 AND5x1_ASAP7_75t_R _14480_ (.A(_06882_),
    .B(_06891_),
    .C(_07062_),
    .D(_07054_),
    .E(_07115_),
    .Y(_07501_));
 AO21x1_ASAP7_75t_R _14481_ (.A1(_07452_),
    .A2(_07487_),
    .B(_06472_),
    .Y(_07502_));
 OAI21x1_ASAP7_75t_R _14482_ (.A1(_07501_),
    .A2(_07502_),
    .B(_06831_),
    .Y(_07503_));
 OA211x2_ASAP7_75t_R _14483_ (.A1(_05841_),
    .A2(_05850_),
    .B(_06848_),
    .C(_06849_),
    .Y(_07504_));
 OR2x2_ASAP7_75t_R _14484_ (.A(_05861_),
    .B(_05870_),
    .Y(_07505_));
 AOI221x1_ASAP7_75t_R _14485_ (.A1(_09652_),
    .A2(_06888_),
    .B1(_07504_),
    .B2(_07505_),
    .C(_06861_),
    .Y(_07506_));
 OA211x2_ASAP7_75t_R _14486_ (.A1(_09645_),
    .A2(_06769_),
    .B(_07083_),
    .C(_06897_),
    .Y(_07507_));
 OR3x1_ASAP7_75t_R _14487_ (.A(_06673_),
    .B(_07506_),
    .C(_07507_),
    .Y(_07508_));
 OA211x2_ASAP7_75t_R _14488_ (.A1(_07042_),
    .A2(_07405_),
    .B(_07508_),
    .C(_06835_),
    .Y(_07509_));
 AOI21x1_ASAP7_75t_R _14489_ (.A1(_07036_),
    .A2(_07292_),
    .B(_07509_),
    .Y(_07510_));
 OR3x1_ASAP7_75t_R _14490_ (.A(_07271_),
    .B(_07296_),
    .C(_07297_),
    .Y(_07511_));
 NAND3x1_ASAP7_75t_R _14491_ (.A(_07037_),
    .B(_07300_),
    .C(_07301_),
    .Y(_07512_));
 AO21x1_ASAP7_75t_R _14492_ (.A1(_07511_),
    .A2(_07512_),
    .B(_07374_),
    .Y(_07513_));
 OA211x2_ASAP7_75t_R _14493_ (.A1(_07054_),
    .A2(_07510_),
    .B(_07513_),
    .C(_06472_),
    .Y(_07514_));
 OAI22x1_ASAP7_75t_R _14494_ (.A1(_06831_),
    .A2(_07500_),
    .B1(_07503_),
    .B2(_07514_),
    .Y(net37));
 INVx1_ASAP7_75t_R _14495_ (.A(_00598_),
    .Y(_07515_));
 AO22x1_ASAP7_75t_R _14496_ (.A1(_01190_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07515_),
    .Y(_07516_));
 AO21x1_ASAP7_75t_R _14497_ (.A1(_07249_),
    .A2(_07516_),
    .B(_07456_),
    .Y(_07517_));
 OA21x2_ASAP7_75t_R _14498_ (.A1(_00665_),
    .A2(_07471_),
    .B(_01193_),
    .Y(_07518_));
 OA211x2_ASAP7_75t_R _14499_ (.A1(_00632_),
    .A2(_07518_),
    .B(_07156_),
    .C(_01191_),
    .Y(_07519_));
 INVx1_ASAP7_75t_R _14500_ (.A(_00599_),
    .Y(_07520_));
 OA21x2_ASAP7_75t_R _14501_ (.A1(_07093_),
    .A2(_07519_),
    .B(_07520_),
    .Y(_07521_));
 OAI21x1_ASAP7_75t_R _14502_ (.A1(_00632_),
    .A2(_07518_),
    .B(_01191_),
    .Y(_07522_));
 AND3x1_ASAP7_75t_R _14503_ (.A(_00599_),
    .B(_07240_),
    .C(_07522_),
    .Y(_07523_));
 AND3x1_ASAP7_75t_R _14504_ (.A(_06836_),
    .B(_07311_),
    .C(_07312_),
    .Y(_07524_));
 AND2x2_ASAP7_75t_R _14505_ (.A(_07036_),
    .B(_07323_),
    .Y(_07525_));
 AO21x1_ASAP7_75t_R _14506_ (.A1(_07324_),
    .A2(_07348_),
    .B(_07049_),
    .Y(_07526_));
 AND2x2_ASAP7_75t_R _14507_ (.A(_09561_),
    .B(_07526_),
    .Y(_07527_));
 AO21x1_ASAP7_75t_R _14508_ (.A1(_06470_),
    .A2(_06833_),
    .B(_07527_),
    .Y(_07528_));
 OA21x2_ASAP7_75t_R _14509_ (.A1(_07524_),
    .A2(_07525_),
    .B(_07528_),
    .Y(_07529_));
 AO32x1_ASAP7_75t_R _14510_ (.A1(_07271_),
    .A2(_07293_),
    .A3(_07317_),
    .B1(_07527_),
    .B2(_07020_),
    .Y(_07530_));
 OR3x1_ASAP7_75t_R _14511_ (.A(_05442_),
    .B(_05465_),
    .C(_06869_),
    .Y(_07531_));
 AND3x1_ASAP7_75t_R _14512_ (.A(_07029_),
    .B(_07128_),
    .C(_07531_),
    .Y(_07532_));
 OA211x2_ASAP7_75t_R _14513_ (.A1(_09645_),
    .A2(_07066_),
    .B(_07083_),
    .C(_07118_),
    .Y(_07533_));
 OR3x2_ASAP7_75t_R _14514_ (.A(_06674_),
    .B(_07532_),
    .C(_07533_),
    .Y(_07534_));
 OR2x2_ASAP7_75t_R _14515_ (.A(_06860_),
    .B(_07416_),
    .Y(_07535_));
 AND3x1_ASAP7_75t_R _14516_ (.A(_06470_),
    .B(_06880_),
    .C(_06893_),
    .Y(_07536_));
 AND3x1_ASAP7_75t_R _14517_ (.A(_07534_),
    .B(_07535_),
    .C(_07536_),
    .Y(_07537_));
 OR4x2_ASAP7_75t_R _14518_ (.A(_06924_),
    .B(_07529_),
    .C(_07530_),
    .D(_07537_),
    .Y(_07538_));
 OA31x2_ASAP7_75t_R _14519_ (.A1(_07517_),
    .A2(_07521_),
    .A3(_07523_),
    .B1(_07538_),
    .Y(net38));
 INVx1_ASAP7_75t_R _14520_ (.A(_01188_),
    .Y(_07539_));
 AO22x1_ASAP7_75t_R _14521_ (.A1(_01189_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07539_),
    .Y(_07540_));
 AND2x2_ASAP7_75t_R _14522_ (.A(_07091_),
    .B(_07540_),
    .Y(_07541_));
 OR2x2_ASAP7_75t_R _14523_ (.A(_06966_),
    .B(_06969_),
    .Y(_07542_));
 AO21x1_ASAP7_75t_R _14524_ (.A1(_07542_),
    .A2(_07156_),
    .B(_07005_),
    .Y(_07543_));
 OAI21x1_ASAP7_75t_R _14525_ (.A1(_07542_),
    .A2(_07009_),
    .B(_00565_),
    .Y(_07544_));
 OA21x2_ASAP7_75t_R _14526_ (.A1(_00565_),
    .A2(_07543_),
    .B(_07544_),
    .Y(_07545_));
 OA211x2_ASAP7_75t_R _14527_ (.A1(_09645_),
    .A2(_07061_),
    .B(_06850_),
    .C(_07029_),
    .Y(_07546_));
 AO31x2_ASAP7_75t_R _14528_ (.A1(_03297_),
    .A2(_07128_),
    .A3(_07531_),
    .B(_07546_),
    .Y(_07547_));
 OR3x1_ASAP7_75t_R _14529_ (.A(_07042_),
    .B(_07442_),
    .C(_07443_),
    .Y(_07548_));
 OA211x2_ASAP7_75t_R _14530_ (.A1(_07150_),
    .A2(_07547_),
    .B(_07548_),
    .C(_06836_),
    .Y(_07549_));
 AND3x1_ASAP7_75t_R _14531_ (.A(_06577_),
    .B(_07337_),
    .C(_07340_),
    .Y(_07550_));
 OA21x2_ASAP7_75t_R _14532_ (.A1(_07549_),
    .A2(_07550_),
    .B(_07056_),
    .Y(_07551_));
 OA21x2_ASAP7_75t_R _14533_ (.A1(_06879_),
    .A2(_07551_),
    .B(_06472_),
    .Y(_07552_));
 OA21x2_ASAP7_75t_R _14534_ (.A1(_07021_),
    .A2(_06878_),
    .B(_07452_),
    .Y(_07553_));
 AND3x4_ASAP7_75t_R _14535_ (.A(_06920_),
    .B(_06835_),
    .C(_06892_),
    .Y(_07554_));
 AND2x2_ASAP7_75t_R _14536_ (.A(_06891_),
    .B(_07554_),
    .Y(_07555_));
 AO21x1_ASAP7_75t_R _14537_ (.A1(_06889_),
    .A2(_07555_),
    .B(_06925_),
    .Y(_07556_));
 OA33x2_ASAP7_75t_R _14538_ (.A1(_06831_),
    .A2(_07541_),
    .A3(_07545_),
    .B1(_07552_),
    .B2(_07553_),
    .B3(_07556_),
    .Y(net39));
 AO21x1_ASAP7_75t_R _14539_ (.A1(_06578_),
    .A2(_07387_),
    .B(_07035_),
    .Y(_07557_));
 OA31x2_ASAP7_75t_R _14540_ (.A1(_05442_),
    .A2(_05465_),
    .A3(_06888_),
    .B1(_06855_),
    .Y(_07558_));
 OA211x2_ASAP7_75t_R _14541_ (.A1(_09645_),
    .A2(_07028_),
    .B(_06850_),
    .C(_07118_),
    .Y(_07559_));
 AOI211x1_ASAP7_75t_R _14542_ (.A1(_07048_),
    .A2(_07558_),
    .B(_07559_),
    .C(_06675_),
    .Y(_07560_));
 AOI21x1_ASAP7_75t_R _14543_ (.A1(_06675_),
    .A2(_07482_),
    .B(_07560_),
    .Y(_07561_));
 NAND2x1_ASAP7_75t_R _14544_ (.A(_07037_),
    .B(_07381_),
    .Y(_07562_));
 OA211x2_ASAP7_75t_R _14545_ (.A1(_06578_),
    .A2(_07561_),
    .B(_07562_),
    .C(_07293_),
    .Y(_07563_));
 AO21x1_ASAP7_75t_R _14546_ (.A1(_07452_),
    .A2(_07557_),
    .B(_07563_),
    .Y(_07564_));
 OA21x2_ASAP7_75t_R _14547_ (.A1(_03555_),
    .A2(_06469_),
    .B(_07049_),
    .Y(_07565_));
 AO21x2_ASAP7_75t_R _14548_ (.A1(_06920_),
    .A2(_07565_),
    .B(_06924_),
    .Y(_07566_));
 AOI21x1_ASAP7_75t_R _14549_ (.A1(_07060_),
    .A2(_07554_),
    .B(_07566_),
    .Y(_07567_));
 OAI21x1_ASAP7_75t_R _14550_ (.A1(_07021_),
    .A2(_07055_),
    .B(_07567_),
    .Y(_07568_));
 INVx1_ASAP7_75t_R _14551_ (.A(_01186_),
    .Y(_07569_));
 AO22x1_ASAP7_75t_R _14552_ (.A1(_01187_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07569_),
    .Y(_07570_));
 AO21x1_ASAP7_75t_R _14553_ (.A1(_07249_),
    .A2(_07570_),
    .B(_07456_),
    .Y(_07571_));
 OR3x1_ASAP7_75t_R _14554_ (.A(_00565_),
    .B(_06967_),
    .C(_07467_),
    .Y(_07572_));
 OR2x2_ASAP7_75t_R _14555_ (.A(_06967_),
    .B(_07470_),
    .Y(_07573_));
 AO21x1_ASAP7_75t_R _14556_ (.A1(_06964_),
    .A2(_07573_),
    .B(_00565_),
    .Y(_07574_));
 OA211x2_ASAP7_75t_R _14557_ (.A1(_07367_),
    .A2(_07572_),
    .B(_07574_),
    .C(_01188_),
    .Y(_07575_));
 AO21x1_ASAP7_75t_R _14558_ (.A1(_07461_),
    .A2(_07575_),
    .B(_07005_),
    .Y(_07576_));
 OAI21x1_ASAP7_75t_R _14559_ (.A1(_07280_),
    .A2(_07575_),
    .B(_00532_),
    .Y(_07577_));
 OA21x2_ASAP7_75t_R _14560_ (.A1(_00532_),
    .A2(_07576_),
    .B(_07577_),
    .Y(_07578_));
 OAI22x1_ASAP7_75t_R _14561_ (.A1(_07564_),
    .A2(_07568_),
    .B1(_07571_),
    .B2(_07578_),
    .Y(_07579_));
 INVx8_ASAP7_75t_R _14562_ (.A(_07579_),
    .Y(net40));
 INVx1_ASAP7_75t_R _14563_ (.A(_00499_),
    .Y(_07580_));
 OA21x2_ASAP7_75t_R _14564_ (.A1(_00565_),
    .A2(_07542_),
    .B(_01188_),
    .Y(_07581_));
 OA21x2_ASAP7_75t_R _14565_ (.A1(_00532_),
    .A2(_07581_),
    .B(_01186_),
    .Y(_07582_));
 AO21x1_ASAP7_75t_R _14566_ (.A1(_07461_),
    .A2(_07582_),
    .B(_07093_),
    .Y(_07583_));
 INVx1_ASAP7_75t_R _14567_ (.A(_07582_),
    .Y(_07584_));
 INVx1_ASAP7_75t_R _14568_ (.A(_01184_),
    .Y(_07585_));
 AO22x1_ASAP7_75t_R _14569_ (.A1(_01185_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07585_),
    .Y(_07586_));
 AO32x1_ASAP7_75t_R _14570_ (.A1(_00499_),
    .A2(_07461_),
    .A3(_07584_),
    .B1(_07586_),
    .B2(_06940_),
    .Y(_07587_));
 AO21x1_ASAP7_75t_R _14571_ (.A1(_07580_),
    .A2(_07583_),
    .B(_07587_),
    .Y(_07588_));
 AND3x1_ASAP7_75t_R _14572_ (.A(_06898_),
    .B(_07031_),
    .C(_07079_),
    .Y(_07589_));
 AO21x1_ASAP7_75t_R _14573_ (.A1(_06902_),
    .A2(_07558_),
    .B(_07589_),
    .Y(_07590_));
 OA21x2_ASAP7_75t_R _14574_ (.A1(_07506_),
    .A2(_07507_),
    .B(_06868_),
    .Y(_07591_));
 AO21x1_ASAP7_75t_R _14575_ (.A1(_07042_),
    .A2(_07590_),
    .B(_07591_),
    .Y(_07592_));
 AO221x1_ASAP7_75t_R _14576_ (.A1(_07110_),
    .A2(_07113_),
    .B1(_07592_),
    .B2(_06893_),
    .C(_06920_),
    .Y(_07593_));
 OA211x2_ASAP7_75t_R _14577_ (.A1(_06471_),
    .A2(_07409_),
    .B(_07593_),
    .C(_06881_),
    .Y(_07594_));
 AND3x1_ASAP7_75t_R _14578_ (.A(_06674_),
    .B(_07062_),
    .C(_07115_),
    .Y(_07595_));
 OA21x2_ASAP7_75t_R _14579_ (.A1(_07121_),
    .A2(_07123_),
    .B(_07022_),
    .Y(_07596_));
 OA21x2_ASAP7_75t_R _14580_ (.A1(_07595_),
    .A2(_07596_),
    .B(_07113_),
    .Y(_07597_));
 OA211x2_ASAP7_75t_R _14581_ (.A1(_07597_),
    .A2(_07407_),
    .B(_06471_),
    .C(_07037_),
    .Y(_07598_));
 AND3x1_ASAP7_75t_R _14582_ (.A(_07112_),
    .B(_07117_),
    .C(_07119_),
    .Y(_07599_));
 OR3x1_ASAP7_75t_R _14583_ (.A(_06880_),
    .B(_07599_),
    .C(_07596_),
    .Y(_07600_));
 OA21x2_ASAP7_75t_R _14584_ (.A1(_06577_),
    .A2(_07110_),
    .B(_07600_),
    .Y(_07601_));
 OA21x2_ASAP7_75t_R _14585_ (.A1(_07020_),
    .A2(_07601_),
    .B(_07565_),
    .Y(_07602_));
 OR4x1_ASAP7_75t_R _14586_ (.A(_06925_),
    .B(_07594_),
    .C(_07598_),
    .D(_07602_),
    .Y(_07603_));
 OA21x2_ASAP7_75t_R _14587_ (.A1(_06831_),
    .A2(_07588_),
    .B(_07603_),
    .Y(net41));
 INVx1_ASAP7_75t_R _14588_ (.A(_01182_),
    .Y(_07604_));
 AO22x1_ASAP7_75t_R _14589_ (.A1(_01183_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07604_),
    .Y(_07605_));
 AO21x1_ASAP7_75t_R _14590_ (.A1(_07249_),
    .A2(_07605_),
    .B(_07456_),
    .Y(_07606_));
 OA21x2_ASAP7_75t_R _14591_ (.A1(_06944_),
    .A2(_07575_),
    .B(_06971_),
    .Y(_07607_));
 AO21x1_ASAP7_75t_R _14592_ (.A1(_07461_),
    .A2(_07607_),
    .B(_07005_),
    .Y(_07608_));
 OAI21x1_ASAP7_75t_R _14593_ (.A1(_07280_),
    .A2(_07607_),
    .B(_00466_),
    .Y(_07609_));
 OA21x2_ASAP7_75t_R _14594_ (.A1(_00466_),
    .A2(_07608_),
    .B(_07609_),
    .Y(_07610_));
 AND3x1_ASAP7_75t_R _14595_ (.A(_07029_),
    .B(_07133_),
    .C(_07103_),
    .Y(_07611_));
 AND3x1_ASAP7_75t_R _14596_ (.A(_03296_),
    .B(_07031_),
    .C(_07079_),
    .Y(_07612_));
 OR3x1_ASAP7_75t_R _14597_ (.A(_07027_),
    .B(_07611_),
    .C(_07612_),
    .Y(_07613_));
 OR3x1_ASAP7_75t_R _14598_ (.A(_06839_),
    .B(_07532_),
    .C(_07533_),
    .Y(_07614_));
 AND3x1_ASAP7_75t_R _14599_ (.A(_06881_),
    .B(_07613_),
    .C(_07614_),
    .Y(_07615_));
 AO21x1_ASAP7_75t_R _14600_ (.A1(_06578_),
    .A2(_07418_),
    .B(_07615_),
    .Y(_07616_));
 AO221x1_ASAP7_75t_R _14601_ (.A1(_07088_),
    .A2(_07188_),
    .B1(_07198_),
    .B2(_07555_),
    .C(_07566_),
    .Y(_07617_));
 AO21x1_ASAP7_75t_R _14602_ (.A1(_07293_),
    .A2(_07616_),
    .B(_07617_),
    .Y(_07618_));
 OA21x2_ASAP7_75t_R _14603_ (.A1(_07606_),
    .A2(_07610_),
    .B(_07618_),
    .Y(net42));
 AND2x2_ASAP7_75t_R _14604_ (.A(_06970_),
    .B(_06972_),
    .Y(_07619_));
 OAI21x1_ASAP7_75t_R _14605_ (.A1(_00466_),
    .A2(_07619_),
    .B(_01182_),
    .Y(_07620_));
 OA21x2_ASAP7_75t_R _14606_ (.A1(_07620_),
    .A2(_07280_),
    .B(_07172_),
    .Y(_07621_));
 NOR2x1_ASAP7_75t_R _14607_ (.A(_00433_),
    .B(_07621_),
    .Y(_07622_));
 INVx1_ASAP7_75t_R _14608_ (.A(_01180_),
    .Y(_07623_));
 AO22x1_ASAP7_75t_R _14609_ (.A1(_01181_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07623_),
    .Y(_07624_));
 AND2x2_ASAP7_75t_R _14610_ (.A(_07620_),
    .B(_07156_),
    .Y(_07625_));
 AO221x1_ASAP7_75t_R _14611_ (.A1(_07091_),
    .A2(_07624_),
    .B1(_07625_),
    .B2(_00433_),
    .C(_06830_),
    .Y(_07626_));
 OA211x2_ASAP7_75t_R _14612_ (.A1(_09625_),
    .A2(_07028_),
    .B(_06844_),
    .C(_06898_),
    .Y(_07627_));
 OA211x2_ASAP7_75t_R _14613_ (.A1(_09620_),
    .A2(_07066_),
    .B(_07133_),
    .C(_07118_),
    .Y(_07628_));
 OR3x1_ASAP7_75t_R _14614_ (.A(_07027_),
    .B(_07627_),
    .C(_07628_),
    .Y(_07629_));
 OA211x2_ASAP7_75t_R _14615_ (.A1(_07043_),
    .A2(_07547_),
    .B(_07629_),
    .C(_06880_),
    .Y(_07630_));
 OA21x2_ASAP7_75t_R _14616_ (.A1(_07444_),
    .A2(_07445_),
    .B(_06577_),
    .Y(_07631_));
 OA21x2_ASAP7_75t_R _14617_ (.A1(_07630_),
    .A2(_07631_),
    .B(_07056_),
    .Y(_07632_));
 AO21x1_ASAP7_75t_R _14618_ (.A1(_07113_),
    .A2(_07232_),
    .B(_07632_),
    .Y(_07633_));
 AO221x1_ASAP7_75t_R _14619_ (.A1(_07215_),
    .A2(_07554_),
    .B1(_07565_),
    .B2(_07235_),
    .C(_07566_),
    .Y(_07634_));
 AO21x1_ASAP7_75t_R _14620_ (.A1(_06472_),
    .A2(_07633_),
    .B(_07634_),
    .Y(_07635_));
 OA21x2_ASAP7_75t_R _14621_ (.A1(_07622_),
    .A2(_07626_),
    .B(_07635_),
    .Y(net44));
 AO21x1_ASAP7_75t_R _14622_ (.A1(_07274_),
    .A2(_07565_),
    .B(_07566_),
    .Y(_07636_));
 OA21x2_ASAP7_75t_R _14623_ (.A1(_09620_),
    .A2(_07028_),
    .B(_06842_),
    .Y(_07637_));
 OA211x2_ASAP7_75t_R _14624_ (.A1(_09625_),
    .A2(_07028_),
    .B(_06844_),
    .C(_07118_),
    .Y(_07638_));
 AO21x1_ASAP7_75t_R _14625_ (.A1(_07063_),
    .A2(_07637_),
    .B(_07638_),
    .Y(_07639_));
 AO211x2_ASAP7_75t_R _14626_ (.A1(_07063_),
    .A2(_07558_),
    .B(_07559_),
    .C(_06839_),
    .Y(_07640_));
 OA21x2_ASAP7_75t_R _14627_ (.A1(_06674_),
    .A2(_07639_),
    .B(_07640_),
    .Y(_07641_));
 AO21x1_ASAP7_75t_R _14628_ (.A1(_07056_),
    .A2(_07641_),
    .B(_07478_),
    .Y(_07642_));
 AND2x2_ASAP7_75t_R _14629_ (.A(_07020_),
    .B(_07256_),
    .Y(_07643_));
 AO221x1_ASAP7_75t_R _14630_ (.A1(_07265_),
    .A2(_07452_),
    .B1(_07642_),
    .B2(_07088_),
    .C(_07643_),
    .Y(_07644_));
 AND2x2_ASAP7_75t_R _14631_ (.A(_06470_),
    .B(_07113_),
    .Y(_07645_));
 AO221x1_ASAP7_75t_R _14632_ (.A1(_07293_),
    .A2(_07484_),
    .B1(_07645_),
    .B2(_07268_),
    .C(_06882_),
    .Y(_07646_));
 OA21x2_ASAP7_75t_R _14633_ (.A1(_06578_),
    .A2(_07644_),
    .B(_07646_),
    .Y(_07647_));
 INVx1_ASAP7_75t_R _14634_ (.A(_01178_),
    .Y(_07648_));
 AO22x1_ASAP7_75t_R _14635_ (.A1(_01179_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07648_),
    .Y(_07649_));
 AO21x1_ASAP7_75t_R _14636_ (.A1(_07249_),
    .A2(_07649_),
    .B(_07456_),
    .Y(_07650_));
 AND3x1_ASAP7_75t_R _14637_ (.A(_01188_),
    .B(_06977_),
    .C(_06971_),
    .Y(_07651_));
 OA211x2_ASAP7_75t_R _14638_ (.A1(_07367_),
    .A2(_07572_),
    .B(_07651_),
    .C(_07574_),
    .Y(_07652_));
 AND3x1_ASAP7_75t_R _14639_ (.A(_06977_),
    .B(_06971_),
    .C(_06944_),
    .Y(_07653_));
 AO21x2_ASAP7_75t_R _14640_ (.A1(_06977_),
    .A2(_06973_),
    .B(_07653_),
    .Y(_07654_));
 OR2x2_ASAP7_75t_R _14641_ (.A(_07652_),
    .B(_07654_),
    .Y(_07655_));
 NAND2x1_ASAP7_75t_R _14642_ (.A(_00400_),
    .B(_07240_),
    .Y(_07656_));
 AOI21x1_ASAP7_75t_R _14643_ (.A1(_07240_),
    .A2(_07655_),
    .B(_07093_),
    .Y(_07657_));
 OAI22x1_ASAP7_75t_R _14644_ (.A1(_07655_),
    .A2(_07656_),
    .B1(_07657_),
    .B2(_00400_),
    .Y(_07658_));
 OA22x2_ASAP7_75t_R _14645_ (.A1(_07636_),
    .A2(_07647_),
    .B1(_07650_),
    .B2(_07658_),
    .Y(net45));
 OA211x2_ASAP7_75t_R _14646_ (.A1(_09615_),
    .A2(_06896_),
    .B(_07024_),
    .C(_06898_),
    .Y(_07659_));
 AO21x1_ASAP7_75t_R _14647_ (.A1(_06902_),
    .A2(_07637_),
    .B(_07659_),
    .Y(_07660_));
 AO211x2_ASAP7_75t_R _14648_ (.A1(_06902_),
    .A2(_07558_),
    .B(_07589_),
    .C(_07022_),
    .Y(_07661_));
 OA21x2_ASAP7_75t_R _14649_ (.A1(_06674_),
    .A2(_07660_),
    .B(_07661_),
    .Y(_07662_));
 AND2x2_ASAP7_75t_R _14650_ (.A(_06881_),
    .B(_07662_),
    .Y(_07663_));
 OA211x2_ASAP7_75t_R _14651_ (.A1(_06891_),
    .A2(_07405_),
    .B(_07508_),
    .C(_06577_),
    .Y(_07664_));
 OA21x2_ASAP7_75t_R _14652_ (.A1(_07663_),
    .A2(_07664_),
    .B(_07374_),
    .Y(_07665_));
 OA21x2_ASAP7_75t_R _14653_ (.A1(_07304_),
    .A2(_07665_),
    .B(_06472_),
    .Y(_07666_));
 OR3x1_ASAP7_75t_R _14654_ (.A(_07020_),
    .B(_07302_),
    .C(_07306_),
    .Y(_07667_));
 AO221x1_ASAP7_75t_R _14655_ (.A1(_07292_),
    .A2(_07554_),
    .B1(_07565_),
    .B2(_07667_),
    .C(_06925_),
    .Y(_07668_));
 OR3x1_ASAP7_75t_R _14656_ (.A(_00400_),
    .B(_07619_),
    .C(_06973_),
    .Y(_07669_));
 NAND2x1_ASAP7_75t_R _14657_ (.A(_06978_),
    .B(_07669_),
    .Y(_07670_));
 OA21x2_ASAP7_75t_R _14658_ (.A1(_07670_),
    .A2(_07009_),
    .B(_07172_),
    .Y(_07671_));
 NOR2x1_ASAP7_75t_R _14659_ (.A(_00367_),
    .B(_07671_),
    .Y(_07672_));
 AND3x1_ASAP7_75t_R _14660_ (.A(_00367_),
    .B(_07670_),
    .C(_07156_),
    .Y(_07673_));
 INVx1_ASAP7_75t_R _14661_ (.A(_01176_),
    .Y(_07674_));
 AO22x1_ASAP7_75t_R _14662_ (.A1(_01177_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07674_),
    .Y(_07675_));
 AO21x1_ASAP7_75t_R _14663_ (.A1(_06940_),
    .A2(_07675_),
    .B(_06830_),
    .Y(_07676_));
 OR3x2_ASAP7_75t_R _14664_ (.A(_07672_),
    .B(_07673_),
    .C(_07676_),
    .Y(_07677_));
 OA21x2_ASAP7_75t_R _14665_ (.A1(_07666_),
    .A2(_07668_),
    .B(_07677_),
    .Y(net46));
 OA211x2_ASAP7_75t_R _14666_ (.A1(_09610_),
    .A2(_06862_),
    .B(_07107_),
    .C(_06897_),
    .Y(_07678_));
 OA211x2_ASAP7_75t_R _14667_ (.A1(_09615_),
    .A2(_06862_),
    .B(_07024_),
    .C(_03295_),
    .Y(_07679_));
 OR3x1_ASAP7_75t_R _14668_ (.A(_07150_),
    .B(_07678_),
    .C(_07679_),
    .Y(_07680_));
 OR3x1_ASAP7_75t_R _14669_ (.A(_07023_),
    .B(_07611_),
    .C(_07612_),
    .Y(_07681_));
 AND3x1_ASAP7_75t_R _14670_ (.A(_06881_),
    .B(_07680_),
    .C(_07681_),
    .Y(_07682_));
 AND3x1_ASAP7_75t_R _14671_ (.A(_07271_),
    .B(_07534_),
    .C(_07535_),
    .Y(_07683_));
 OA21x2_ASAP7_75t_R _14672_ (.A1(_07682_),
    .A2(_07683_),
    .B(_07088_),
    .Y(_07684_));
 AND3x1_ASAP7_75t_R _14673_ (.A(_07020_),
    .B(_07190_),
    .C(_07317_),
    .Y(_07685_));
 OA21x2_ASAP7_75t_R _14674_ (.A1(_07684_),
    .A2(_07685_),
    .B(_07374_),
    .Y(_07686_));
 AO21x1_ASAP7_75t_R _14675_ (.A1(_07088_),
    .A2(_07054_),
    .B(_07452_),
    .Y(_07687_));
 AO21x1_ASAP7_75t_R _14676_ (.A1(_07326_),
    .A2(_07687_),
    .B(_07566_),
    .Y(_07688_));
 INVx1_ASAP7_75t_R _14677_ (.A(_00333_),
    .Y(_07689_));
 AO22x1_ASAP7_75t_R _14678_ (.A1(_01175_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07689_),
    .Y(_07690_));
 AO21x1_ASAP7_75t_R _14679_ (.A1(_07249_),
    .A2(_07690_),
    .B(_07456_),
    .Y(_07691_));
 OA21x2_ASAP7_75t_R _14680_ (.A1(_00367_),
    .A2(_01178_),
    .B(_01176_),
    .Y(_07692_));
 OA31x2_ASAP7_75t_R _14681_ (.A1(_06974_),
    .A2(_07652_),
    .A3(_07654_),
    .B1(_07692_),
    .Y(_07693_));
 AO21x1_ASAP7_75t_R _14682_ (.A1(_07461_),
    .A2(_07693_),
    .B(_07005_),
    .Y(_07694_));
 OAI21x1_ASAP7_75t_R _14683_ (.A1(_07280_),
    .A2(_07693_),
    .B(_00334_),
    .Y(_07695_));
 OA21x2_ASAP7_75t_R _14684_ (.A1(_00334_),
    .A2(_07694_),
    .B(_07695_),
    .Y(_07696_));
 OA22x2_ASAP7_75t_R _14685_ (.A1(_07686_),
    .A2(_07688_),
    .B1(_07691_),
    .B2(_07696_),
    .Y(net47));
 AO21x1_ASAP7_75t_R _14686_ (.A1(_06976_),
    .A2(_06979_),
    .B(_00334_),
    .Y(_07697_));
 NAND2x1_ASAP7_75t_R _14687_ (.A(_00333_),
    .B(_07697_),
    .Y(_07698_));
 OA21x2_ASAP7_75t_R _14688_ (.A1(_07698_),
    .A2(_07009_),
    .B(_07172_),
    .Y(_07699_));
 INVx1_ASAP7_75t_R _14689_ (.A(_01173_),
    .Y(_07700_));
 AO22x1_ASAP7_75t_R _14690_ (.A1(_01174_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07700_),
    .Y(_07701_));
 AND4x1_ASAP7_75t_R _14691_ (.A(_00300_),
    .B(_07698_),
    .C(_07172_),
    .D(_07156_),
    .Y(_07702_));
 AOI21x1_ASAP7_75t_R _14692_ (.A1(_07091_),
    .A2(_07701_),
    .B(_07702_),
    .Y(_07703_));
 OA21x2_ASAP7_75t_R _14693_ (.A1(_00300_),
    .A2(_07699_),
    .B(_07703_),
    .Y(_07704_));
 OA211x2_ASAP7_75t_R _14694_ (.A1(_06675_),
    .A2(_07547_),
    .B(_07548_),
    .C(_07036_),
    .Y(_07705_));
 INVx1_ASAP7_75t_R _14695_ (.A(_07705_),
    .Y(_07706_));
 NOR3x1_ASAP7_75t_R _14696_ (.A(_07043_),
    .B(_07627_),
    .C(_07628_),
    .Y(_07707_));
 NAND2x1_ASAP7_75t_R _14697_ (.A(_07102_),
    .B(_07107_),
    .Y(_07708_));
 OR2x2_ASAP7_75t_R _14698_ (.A(_09605_),
    .B(_06896_),
    .Y(_07709_));
 OR2x2_ASAP7_75t_R _14699_ (.A(_09595_),
    .B(_06769_),
    .Y(_07710_));
 NAND3x1_ASAP7_75t_R _14700_ (.A(_07063_),
    .B(_07709_),
    .C(_07710_),
    .Y(_07711_));
 OA211x2_ASAP7_75t_R _14701_ (.A1(_07048_),
    .A2(_07708_),
    .B(_07711_),
    .C(_06860_),
    .Y(_07712_));
 OR3x1_ASAP7_75t_R _14702_ (.A(_07271_),
    .B(_07707_),
    .C(_07712_),
    .Y(_07713_));
 AO21x1_ASAP7_75t_R _14703_ (.A1(_07706_),
    .A2(_07713_),
    .B(_07054_),
    .Y(_07714_));
 NOR2x1_ASAP7_75t_R _14704_ (.A(_06921_),
    .B(_07350_),
    .Y(_07715_));
 AOI21x1_ASAP7_75t_R _14705_ (.A1(_07374_),
    .A2(_07341_),
    .B(_07452_),
    .Y(_07716_));
 AO221x1_ASAP7_75t_R _14706_ (.A1(_07714_),
    .A2(_07715_),
    .B1(_07716_),
    .B2(_07021_),
    .C(_06925_),
    .Y(_07717_));
 OAI21x1_ASAP7_75t_R _14707_ (.A1(_06831_),
    .A2(_07704_),
    .B(_07717_),
    .Y(net48));
 INVx1_ASAP7_75t_R _14708_ (.A(_01171_),
    .Y(_07718_));
 AO22x1_ASAP7_75t_R _14709_ (.A1(_01172_),
    .A2(_07160_),
    .B1(_07161_),
    .B2(_07718_),
    .Y(_07719_));
 OR2x2_ASAP7_75t_R _14710_ (.A(_00300_),
    .B(_00334_),
    .Y(_07720_));
 OA21x2_ASAP7_75t_R _14711_ (.A1(_00300_),
    .A2(_00333_),
    .B(_01173_),
    .Y(_07721_));
 OA21x2_ASAP7_75t_R _14712_ (.A1(_07692_),
    .A2(_07720_),
    .B(_07721_),
    .Y(_07722_));
 OR2x2_ASAP7_75t_R _14713_ (.A(_06974_),
    .B(_07720_),
    .Y(_07723_));
 AND2x2_ASAP7_75t_R _14714_ (.A(_07722_),
    .B(_07723_),
    .Y(_07724_));
 AO21x1_ASAP7_75t_R _14715_ (.A1(_07156_),
    .A2(_07724_),
    .B(_07005_),
    .Y(_07725_));
 INVx1_ASAP7_75t_R _14716_ (.A(_00267_),
    .Y(_07726_));
 AO221x1_ASAP7_75t_R _14717_ (.A1(_07091_),
    .A2(_07719_),
    .B1(_07725_),
    .B2(_07726_),
    .C(_07456_),
    .Y(_07727_));
 OR3x1_ASAP7_75t_R _14718_ (.A(_07652_),
    .B(_07654_),
    .C(_07723_),
    .Y(_07728_));
 AOI21x1_ASAP7_75t_R _14719_ (.A1(_07722_),
    .A2(_07728_),
    .B(_07726_),
    .Y(_07729_));
 AND3x1_ASAP7_75t_R _14720_ (.A(_07726_),
    .B(_07655_),
    .C(_07722_),
    .Y(_07730_));
 OA21x2_ASAP7_75t_R _14721_ (.A1(_07729_),
    .A2(_07730_),
    .B(_07240_),
    .Y(_07731_));
 OA211x2_ASAP7_75t_R _14722_ (.A1(_07037_),
    .A2(_07387_),
    .B(_07565_),
    .C(_07347_),
    .Y(_07732_));
 AND4x1_ASAP7_75t_R _14723_ (.A(_06471_),
    .B(_07041_),
    .C(_07348_),
    .D(_07386_),
    .Y(_07733_));
 OR3x1_ASAP7_75t_R _14724_ (.A(_07566_),
    .B(_07732_),
    .C(_07733_),
    .Y(_07734_));
 OA21x2_ASAP7_75t_R _14725_ (.A1(_09600_),
    .A2(_07062_),
    .B(_06874_),
    .Y(_07735_));
 AND3x1_ASAP7_75t_R _14726_ (.A(_03297_),
    .B(_07709_),
    .C(_07710_),
    .Y(_07736_));
 AO21x1_ASAP7_75t_R _14727_ (.A1(_07048_),
    .A2(_07735_),
    .B(_07736_),
    .Y(_07737_));
 OR2x2_ASAP7_75t_R _14728_ (.A(_07043_),
    .B(_07639_),
    .Y(_07738_));
 OA211x2_ASAP7_75t_R _14729_ (.A1(_06675_),
    .A2(_07737_),
    .B(_07738_),
    .C(_07190_),
    .Y(_07739_));
 AOI21x1_ASAP7_75t_R _14730_ (.A1(_06578_),
    .A2(_07561_),
    .B(_07739_),
    .Y(_07740_));
 AO21x1_ASAP7_75t_R _14731_ (.A1(_06921_),
    .A2(_07383_),
    .B(_07054_),
    .Y(_07741_));
 AOI21x1_ASAP7_75t_R _14732_ (.A1(_06472_),
    .A2(_07740_),
    .B(_07741_),
    .Y(_07742_));
 OAI22x1_ASAP7_75t_R _14733_ (.A1(_07727_),
    .A2(_07731_),
    .B1(_07734_),
    .B2(_07742_),
    .Y(_07743_));
 CKINVDCx8_ASAP7_75t_R _14734_ (.A(_07743_),
    .Y(net49));
 OR3x1_ASAP7_75t_R _14735_ (.A(_06823_),
    .B(_04338_),
    .C(_04359_),
    .Y(_07744_));
 OA21x2_ASAP7_75t_R _14736_ (.A1(_06840_),
    .A2(_09585_),
    .B(_07744_),
    .Y(_07745_));
 AO221x1_ASAP7_75t_R _14737_ (.A1(_04439_),
    .A2(_04457_),
    .B1(_04483_),
    .B2(_06713_),
    .C(_03294_),
    .Y(_07746_));
 OA211x2_ASAP7_75t_R _14738_ (.A1(_06851_),
    .A2(_09600_),
    .B(_06869_),
    .C(_07746_),
    .Y(_07747_));
 AO21x1_ASAP7_75t_R _14739_ (.A1(_07028_),
    .A2(_07745_),
    .B(_07747_),
    .Y(_07748_));
 OR2x2_ASAP7_75t_R _14740_ (.A(_07112_),
    .B(_07748_),
    .Y(_07749_));
 OA211x2_ASAP7_75t_R _14741_ (.A1(_07023_),
    .A2(_07660_),
    .B(_07749_),
    .C(_06880_),
    .Y(_07750_));
 AO21x1_ASAP7_75t_R _14742_ (.A1(_07037_),
    .A2(_07592_),
    .B(_07750_),
    .Y(_07751_));
 AO21x1_ASAP7_75t_R _14743_ (.A1(_07374_),
    .A2(_07751_),
    .B(_07400_),
    .Y(_07752_));
 INVx1_ASAP7_75t_R _14744_ (.A(_00234_),
    .Y(_07753_));
 AO21x1_ASAP7_75t_R _14745_ (.A1(_01173_),
    .A2(_06981_),
    .B(_00267_),
    .Y(_07754_));
 AND2x2_ASAP7_75t_R _14746_ (.A(_01171_),
    .B(_07754_),
    .Y(_07755_));
 XNOR2x1_ASAP7_75t_R _14747_ (.B(_07755_),
    .Y(_07756_),
    .A(_07753_));
 INVx1_ASAP7_75t_R _14748_ (.A(_00233_),
    .Y(_07757_));
 AO22x1_ASAP7_75t_R _14749_ (.A1(_01170_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07757_),
    .Y(_07758_));
 AO221x1_ASAP7_75t_R _14750_ (.A1(_07753_),
    .A2(_07001_),
    .B1(_07758_),
    .B2(_06939_),
    .C(_06829_),
    .Y(_07759_));
 AO21x1_ASAP7_75t_R _14751_ (.A1(_07461_),
    .A2(_07756_),
    .B(_07759_),
    .Y(_07760_));
 OA211x2_ASAP7_75t_R _14752_ (.A1(_06674_),
    .A2(_07405_),
    .B(_07406_),
    .C(_06835_),
    .Y(_07761_));
 OA211x2_ASAP7_75t_R _14753_ (.A1(_06886_),
    .A2(_07143_),
    .B(_06576_),
    .C(_07042_),
    .Y(_07762_));
 OA21x2_ASAP7_75t_R _14754_ (.A1(_07761_),
    .A2(_07762_),
    .B(_06893_),
    .Y(_07763_));
 OR4x1_ASAP7_75t_R _14755_ (.A(_06471_),
    .B(_06924_),
    .C(_07451_),
    .D(_07763_),
    .Y(_07764_));
 OA211x2_ASAP7_75t_R _14756_ (.A1(_07223_),
    .A2(_07752_),
    .B(_07760_),
    .C(_07764_),
    .Y(_07765_));
 BUFx12_ASAP7_75t_R _14757_ (.A(_07765_),
    .Y(net50));
 OR3x1_ASAP7_75t_R _14758_ (.A(_00234_),
    .B(_00267_),
    .C(_07720_),
    .Y(_07766_));
 OA21x2_ASAP7_75t_R _14759_ (.A1(_00267_),
    .A2(_07721_),
    .B(_01171_),
    .Y(_07767_));
 OA21x2_ASAP7_75t_R _14760_ (.A1(_00234_),
    .A2(_07767_),
    .B(_00233_),
    .Y(_07768_));
 OA211x2_ASAP7_75t_R _14761_ (.A1(_07693_),
    .A2(_07766_),
    .B(_07768_),
    .C(_07004_),
    .Y(_07769_));
 INVx1_ASAP7_75t_R _14762_ (.A(_00200_),
    .Y(_07770_));
 AO22x1_ASAP7_75t_R _14763_ (.A1(_01169_),
    .A2(_06999_),
    .B1(_07013_),
    .B2(_07770_),
    .Y(_07771_));
 AO21x1_ASAP7_75t_R _14764_ (.A1(_06939_),
    .A2(_07771_),
    .B(_06829_),
    .Y(_07772_));
 OR4x1_ASAP7_75t_R _14765_ (.A(_01168_),
    .B(_07005_),
    .C(_07769_),
    .D(_07772_),
    .Y(_07773_));
 AO22x1_ASAP7_75t_R _14766_ (.A1(_07198_),
    .A2(_07231_),
    .B1(_07418_),
    .B2(_06836_),
    .Y(_07774_));
 AND3x1_ASAP7_75t_R _14767_ (.A(_07020_),
    .B(_07056_),
    .C(_07774_),
    .Y(_07775_));
 OAI21x1_ASAP7_75t_R _14768_ (.A1(_06920_),
    .A2(_07423_),
    .B(_09563_),
    .Y(_07776_));
 OR3x1_ASAP7_75t_R _14769_ (.A(_06920_),
    .B(_07184_),
    .C(_07423_),
    .Y(_07777_));
 AND3x1_ASAP7_75t_R _14770_ (.A(_07236_),
    .B(_07776_),
    .C(_07777_),
    .Y(_07778_));
 OR3x1_ASAP7_75t_R _14771_ (.A(_06897_),
    .B(_04239_),
    .C(_04265_),
    .Y(_07779_));
 OA21x2_ASAP7_75t_R _14772_ (.A1(_06840_),
    .A2(_09580_),
    .B(_07779_),
    .Y(_07780_));
 OR3x1_ASAP7_75t_R _14773_ (.A(_03295_),
    .B(_04338_),
    .C(_04359_),
    .Y(_07781_));
 OA211x2_ASAP7_75t_R _14774_ (.A1(_06861_),
    .A2(_09595_),
    .B(_06769_),
    .C(_07781_),
    .Y(_07782_));
 AO21x1_ASAP7_75t_R _14775_ (.A1(_07061_),
    .A2(_07780_),
    .B(_07782_),
    .Y(_07783_));
 OR3x1_ASAP7_75t_R _14776_ (.A(_06838_),
    .B(_07678_),
    .C(_07679_),
    .Y(_07784_));
 OA211x2_ASAP7_75t_R _14777_ (.A1(_07112_),
    .A2(_07783_),
    .B(_07784_),
    .C(_06834_),
    .Y(_07785_));
 AO31x2_ASAP7_75t_R _14778_ (.A1(_07036_),
    .A2(_07613_),
    .A3(_07614_),
    .B(_07785_),
    .Y(_07786_));
 AO32x1_ASAP7_75t_R _14779_ (.A1(_06470_),
    .A2(_07348_),
    .A3(_07422_),
    .B1(_07786_),
    .B2(_07293_),
    .Y(_07787_));
 OR4x1_ASAP7_75t_R _14780_ (.A(_06924_),
    .B(_07775_),
    .C(_07778_),
    .D(_07787_),
    .Y(_07788_));
 OR4x1_ASAP7_75t_R _14781_ (.A(_06974_),
    .B(_07009_),
    .C(_07655_),
    .D(_07766_),
    .Y(_07789_));
 OA21x2_ASAP7_75t_R _14782_ (.A1(_07692_),
    .A2(_07766_),
    .B(_07768_),
    .Y(_07790_));
 INVx1_ASAP7_75t_R _14783_ (.A(_07772_),
    .Y(_07791_));
 OA211x2_ASAP7_75t_R _14784_ (.A1(_07009_),
    .A2(_07790_),
    .B(_07791_),
    .C(_01168_),
    .Y(_07792_));
 NAND2x1_ASAP7_75t_R _14785_ (.A(_07789_),
    .B(_07792_),
    .Y(_07793_));
 AND3x4_ASAP7_75t_R _14786_ (.A(_07773_),
    .B(_07788_),
    .C(_07793_),
    .Y(net51));
 OA21x2_ASAP7_75t_R _14787_ (.A1(_06981_),
    .A2(_06983_),
    .B(_06987_),
    .Y(_07794_));
 AO21x1_ASAP7_75t_R _14788_ (.A1(_07240_),
    .A2(_07794_),
    .B(_07093_),
    .Y(_07795_));
 OAI21x1_ASAP7_75t_R _14789_ (.A1(_07280_),
    .A2(_07794_),
    .B(_06982_),
    .Y(_07796_));
 OA21x2_ASAP7_75t_R _14790_ (.A1(_06982_),
    .A2(_07795_),
    .B(_07796_),
    .Y(_07797_));
 INVx1_ASAP7_75t_R _14791_ (.A(_00166_),
    .Y(_07798_));
 AO22x1_ASAP7_75t_R _14792_ (.A1(_01167_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07798_),
    .Y(_07799_));
 AO21x1_ASAP7_75t_R _14793_ (.A1(_07249_),
    .A2(_07799_),
    .B(_07456_),
    .Y(_07800_));
 AND2x2_ASAP7_75t_R _14794_ (.A(_06851_),
    .B(_09577_),
    .Y(_07801_));
 AND2x2_ASAP7_75t_R _14795_ (.A(_06856_),
    .B(_09582_),
    .Y(_07802_));
 OAI21x1_ASAP7_75t_R _14796_ (.A1(_07801_),
    .A2(_07802_),
    .B(_07062_),
    .Y(_07803_));
 OA21x2_ASAP7_75t_R _14797_ (.A1(_07062_),
    .A2(_07745_),
    .B(_07803_),
    .Y(_07804_));
 OA21x2_ASAP7_75t_R _14798_ (.A1(_07048_),
    .A2(_07708_),
    .B(_07711_),
    .Y(_07805_));
 NAND2x1_ASAP7_75t_R _14799_ (.A(_07150_),
    .B(_07805_),
    .Y(_07806_));
 OA211x2_ASAP7_75t_R _14800_ (.A1(_06675_),
    .A2(_07804_),
    .B(_07806_),
    .C(_06836_),
    .Y(_07807_));
 OA211x2_ASAP7_75t_R _14801_ (.A1(_06891_),
    .A2(_07547_),
    .B(_07629_),
    .C(_06577_),
    .Y(_07808_));
 OA211x2_ASAP7_75t_R _14802_ (.A1(_07807_),
    .A2(_07808_),
    .B(_06471_),
    .C(_07374_),
    .Y(_07809_));
 OA21x2_ASAP7_75t_R _14803_ (.A1(_07452_),
    .A2(_07447_),
    .B(_06921_),
    .Y(_07810_));
 AND4x1_ASAP7_75t_R _14804_ (.A(_06470_),
    .B(_06836_),
    .C(_06891_),
    .D(_06833_),
    .Y(_07811_));
 OA22x2_ASAP7_75t_R _14805_ (.A1(_06867_),
    .A2(_07423_),
    .B1(_07811_),
    .B2(_07452_),
    .Y(_07812_));
 OR4x1_ASAP7_75t_R _14806_ (.A(_06925_),
    .B(_07809_),
    .C(_07810_),
    .D(_07812_),
    .Y(_07813_));
 OA21x2_ASAP7_75t_R _14807_ (.A1(_07797_),
    .A2(_07800_),
    .B(_07813_),
    .Y(net52));
 INVx1_ASAP7_75t_R _14808_ (.A(_00133_),
    .Y(_07814_));
 AO22x1_ASAP7_75t_R _14809_ (.A1(_01166_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07814_),
    .Y(_07815_));
 AO21x1_ASAP7_75t_R _14810_ (.A1(_07249_),
    .A2(_07815_),
    .B(_07456_),
    .Y(_07816_));
 OR3x1_ASAP7_75t_R _14811_ (.A(_06982_),
    .B(_06983_),
    .C(_07723_),
    .Y(_07817_));
 OA21x2_ASAP7_75t_R _14812_ (.A1(_01168_),
    .A2(_07790_),
    .B(_00200_),
    .Y(_07818_));
 OA21x2_ASAP7_75t_R _14813_ (.A1(_06982_),
    .A2(_07818_),
    .B(_00166_),
    .Y(_07819_));
 OA31x2_ASAP7_75t_R _14814_ (.A1(_07652_),
    .A2(_07654_),
    .A3(_07817_),
    .B1(_07819_),
    .Y(_07820_));
 AO21x1_ASAP7_75t_R _14815_ (.A1(_07461_),
    .A2(_07820_),
    .B(_07005_),
    .Y(_07821_));
 OAI21x1_ASAP7_75t_R _14816_ (.A1(_07280_),
    .A2(_07820_),
    .B(_01165_),
    .Y(_07822_));
 OA21x2_ASAP7_75t_R _14817_ (.A1(_01165_),
    .A2(_07821_),
    .B(_07822_),
    .Y(_07823_));
 AND3x1_ASAP7_75t_R _14818_ (.A(_07020_),
    .B(_07271_),
    .C(_06893_),
    .Y(_07824_));
 OA21x2_ASAP7_75t_R _14819_ (.A1(_07254_),
    .A2(_07255_),
    .B(_07824_),
    .Y(_07825_));
 AND3x1_ASAP7_75t_R _14820_ (.A(_06471_),
    .B(_07268_),
    .C(_07348_),
    .Y(_07826_));
 OA211x2_ASAP7_75t_R _14821_ (.A1(_06883_),
    .A2(_09575_),
    .B(_07061_),
    .C(_07045_),
    .Y(_07827_));
 AO21x1_ASAP7_75t_R _14822_ (.A1(_06770_),
    .A2(_07780_),
    .B(_07827_),
    .Y(_07828_));
 AND2x2_ASAP7_75t_R _14823_ (.A(_07023_),
    .B(_07828_),
    .Y(_07829_));
 AO21x1_ASAP7_75t_R _14824_ (.A1(_06675_),
    .A2(_07737_),
    .B(_07829_),
    .Y(_07830_));
 AND3x1_ASAP7_75t_R _14825_ (.A(_07271_),
    .B(_07293_),
    .C(_07641_),
    .Y(_07831_));
 AO21x1_ASAP7_75t_R _14826_ (.A1(_07536_),
    .A2(_07830_),
    .B(_07831_),
    .Y(_07832_));
 AO221x1_ASAP7_75t_R _14827_ (.A1(_07484_),
    .A2(_07554_),
    .B1(_07565_),
    .B2(_07489_),
    .C(_07566_),
    .Y(_07833_));
 OR4x1_ASAP7_75t_R _14828_ (.A(_07825_),
    .B(_07826_),
    .C(_07832_),
    .D(_07833_),
    .Y(_07834_));
 OA21x2_ASAP7_75t_R _14829_ (.A1(_07816_),
    .A2(_07823_),
    .B(_07834_),
    .Y(net53));
 AND5x1_ASAP7_75t_R _14830_ (.A(_06470_),
    .B(_06836_),
    .C(_07043_),
    .D(_07062_),
    .E(_07076_),
    .Y(_07835_));
 OA22x2_ASAP7_75t_R _14831_ (.A1(_07115_),
    .A2(_07487_),
    .B1(_07835_),
    .B2(_07452_),
    .Y(_07836_));
 NOR3x1_ASAP7_75t_R _14832_ (.A(_07061_),
    .B(_07801_),
    .C(_07802_),
    .Y(_07837_));
 OA211x2_ASAP7_75t_R _14833_ (.A1(_06861_),
    .A2(_09570_),
    .B(_06896_),
    .C(_07114_),
    .Y(_07838_));
 OR3x1_ASAP7_75t_R _14834_ (.A(_06868_),
    .B(_07837_),
    .C(_07838_),
    .Y(_07839_));
 OA211x2_ASAP7_75t_R _14835_ (.A1(_06860_),
    .A2(_07748_),
    .B(_07839_),
    .C(_06835_),
    .Y(_07840_));
 AO21x1_ASAP7_75t_R _14836_ (.A1(_06577_),
    .A2(_07662_),
    .B(_07840_),
    .Y(_07841_));
 NAND2x1_ASAP7_75t_R _14837_ (.A(_07020_),
    .B(_07510_),
    .Y(_07842_));
 OA211x2_ASAP7_75t_R _14838_ (.A1(_07020_),
    .A2(_07841_),
    .B(_07842_),
    .C(_07056_),
    .Y(_07843_));
 INVx1_ASAP7_75t_R _14839_ (.A(_00099_),
    .Y(_07844_));
 AO22x1_ASAP7_75t_R _14840_ (.A1(_01164_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07844_),
    .Y(_07845_));
 AO21x1_ASAP7_75t_R _14841_ (.A1(_06940_),
    .A2(_07845_),
    .B(_06830_),
    .Y(_07846_));
 INVx1_ASAP7_75t_R _14842_ (.A(_00100_),
    .Y(_07847_));
 AND5x1_ASAP7_75t_R _14843_ (.A(_07847_),
    .B(_00166_),
    .C(_00133_),
    .D(_07004_),
    .E(_07794_),
    .Y(_07848_));
 OA21x2_ASAP7_75t_R _14844_ (.A1(_06982_),
    .A2(_07794_),
    .B(_00166_),
    .Y(_07849_));
 OA21x2_ASAP7_75t_R _14845_ (.A1(_01165_),
    .A2(_07849_),
    .B(_00133_),
    .Y(_07850_));
 NOR2x1_ASAP7_75t_R _14846_ (.A(_07008_),
    .B(_07850_),
    .Y(_07851_));
 AO21x1_ASAP7_75t_R _14847_ (.A1(_00166_),
    .A2(_06982_),
    .B(_01165_),
    .Y(_07852_));
 AND3x1_ASAP7_75t_R _14848_ (.A(_00133_),
    .B(_07003_),
    .C(_07852_),
    .Y(_07853_));
 OR3x1_ASAP7_75t_R _14849_ (.A(_00100_),
    .B(_07001_),
    .C(_07853_),
    .Y(_07854_));
 OA21x2_ASAP7_75t_R _14850_ (.A1(_07847_),
    .A2(_07851_),
    .B(_07854_),
    .Y(_07855_));
 OA33x2_ASAP7_75t_R _14851_ (.A1(_07566_),
    .A2(_07836_),
    .A3(_07843_),
    .B1(_07846_),
    .B2(_07848_),
    .B3(_07855_),
    .Y(net55));
 INVx1_ASAP7_75t_R _14852_ (.A(_01162_),
    .Y(_07856_));
 OA21x2_ASAP7_75t_R _14853_ (.A1(_06982_),
    .A2(_00200_),
    .B(_00166_),
    .Y(_07857_));
 OA21x2_ASAP7_75t_R _14854_ (.A1(_00234_),
    .A2(_01171_),
    .B(_00233_),
    .Y(_07858_));
 OR3x1_ASAP7_75t_R _14855_ (.A(_06982_),
    .B(_01168_),
    .C(_07858_),
    .Y(_07859_));
 AO21x1_ASAP7_75t_R _14856_ (.A1(_07857_),
    .A2(_07859_),
    .B(_01165_),
    .Y(_07860_));
 AO21x1_ASAP7_75t_R _14857_ (.A1(_00133_),
    .A2(_07860_),
    .B(_00100_),
    .Y(_07861_));
 OA211x2_ASAP7_75t_R _14858_ (.A1(_06984_),
    .A2(_07722_),
    .B(_07861_),
    .C(_00099_),
    .Y(_07862_));
 OA21x2_ASAP7_75t_R _14859_ (.A1(_06984_),
    .A2(_07728_),
    .B(_07862_),
    .Y(_07863_));
 XNOR2x1_ASAP7_75t_R _14860_ (.B(_07863_),
    .Y(_07864_),
    .A(_07856_));
 INVx1_ASAP7_75t_R _14861_ (.A(_01161_),
    .Y(_07865_));
 AO22x1_ASAP7_75t_R _14862_ (.A1(_01163_),
    .A2(_07092_),
    .B1(_07097_),
    .B2(_07865_),
    .Y(_07866_));
 AO222x2_ASAP7_75t_R _14863_ (.A1(_07856_),
    .A2(_07093_),
    .B1(_07240_),
    .B2(_07864_),
    .C1(_07866_),
    .C2(_07249_),
    .Y(_07867_));
 AO33x2_ASAP7_75t_R _14864_ (.A1(_03025_),
    .A2(net22),
    .A3(_06833_),
    .B1(_07324_),
    .B2(_07348_),
    .B3(_06471_),
    .Y(_07868_));
 AO21x1_ASAP7_75t_R _14865_ (.A1(_09561_),
    .A2(_07868_),
    .B(_06925_),
    .Y(_07869_));
 AND3x1_ASAP7_75t_R _14866_ (.A(_07190_),
    .B(_07534_),
    .C(_07535_),
    .Y(_07870_));
 AND2x2_ASAP7_75t_R _14867_ (.A(_07037_),
    .B(_07317_),
    .Y(_07871_));
 OA211x2_ASAP7_75t_R _14868_ (.A1(_07870_),
    .A2(_07871_),
    .B(_07021_),
    .C(_07374_),
    .Y(_07872_));
 OA21x2_ASAP7_75t_R _14869_ (.A1(_09561_),
    .A2(_06770_),
    .B(_07122_),
    .Y(_07873_));
 NAND2x1_ASAP7_75t_R _14870_ (.A(_09565_),
    .B(_07044_),
    .Y(_07874_));
 OA211x2_ASAP7_75t_R _14871_ (.A1(_09577_),
    .A2(_07044_),
    .B(_07874_),
    .C(_03297_),
    .Y(_07875_));
 INVx1_ASAP7_75t_R _14872_ (.A(_07875_),
    .Y(_07876_));
 OA211x2_ASAP7_75t_R _14873_ (.A1(_03297_),
    .A2(_07873_),
    .B(_07876_),
    .C(_07043_),
    .Y(_07877_));
 AO21x1_ASAP7_75t_R _14874_ (.A1(_06675_),
    .A2(_07783_),
    .B(_07877_),
    .Y(_07878_));
 AO21x1_ASAP7_75t_R _14875_ (.A1(_07680_),
    .A2(_07681_),
    .B(_07190_),
    .Y(_07879_));
 OA211x2_ASAP7_75t_R _14876_ (.A1(_06578_),
    .A2(_07878_),
    .B(_07879_),
    .C(_07293_),
    .Y(_07880_));
 OR3x1_ASAP7_75t_R _14877_ (.A(_07869_),
    .B(_07872_),
    .C(_07880_),
    .Y(_07881_));
 OA21x2_ASAP7_75t_R _14878_ (.A1(_06831_),
    .A2(_07867_),
    .B(_07881_),
    .Y(net56));
 CKINVDCx20_ASAP7_75t_R _14879_ (.A(net31),
    .Y(_01219_));
 BUFx3_ASAP7_75t_R _14880_ (.A(_05092_),
    .Y(_07882_));
 AO21x1_ASAP7_75t_R _14881_ (.A1(_03024_),
    .A2(net26),
    .B(_03238_),
    .Y(_07883_));
 OR3x4_ASAP7_75t_R _14882_ (.A(_03284_),
    .B(_03288_),
    .C(_07883_),
    .Y(_07884_));
 BUFx3_ASAP7_75t_R _14883_ (.A(_07884_),
    .Y(_07885_));
 AND2x2_ASAP7_75t_R _14884_ (.A(_07882_),
    .B(_07885_),
    .Y(_07886_));
 BUFx4f_ASAP7_75t_R _14885_ (.A(_07886_),
    .Y(_07887_));
 NAND2x2_ASAP7_75t_R _14886_ (.A(_04984_),
    .B(_07884_),
    .Y(_07888_));
 BUFx4f_ASAP7_75t_R _14887_ (.A(_07888_),
    .Y(_07889_));
 OR3x1_ASAP7_75t_R _14888_ (.A(_03427_),
    .B(_03496_),
    .C(_07889_),
    .Y(_07890_));
 OA21x2_ASAP7_75t_R _14889_ (.A1(net65),
    .A2(_07887_),
    .B(_07890_),
    .Y(_09713_));
 OR3x1_ASAP7_75t_R _14890_ (.A(_06797_),
    .B(_06821_),
    .C(_07889_),
    .Y(_07891_));
 OA21x2_ASAP7_75t_R _14891_ (.A1(net76),
    .A2(_07887_),
    .B(_07891_),
    .Y(_09552_));
 BUFx3_ASAP7_75t_R _14892_ (.A(_07888_),
    .Y(_07892_));
 BUFx3_ASAP7_75t_R _14893_ (.A(_07882_),
    .Y(_07893_));
 BUFx3_ASAP7_75t_R _14894_ (.A(_07885_),
    .Y(_07894_));
 AO21x1_ASAP7_75t_R _14895_ (.A1(_07893_),
    .A2(_07894_),
    .B(net87),
    .Y(_07895_));
 OA21x2_ASAP7_75t_R _14896_ (.A1(_09705_),
    .A2(_07892_),
    .B(_07895_),
    .Y(_09715_));
 AO21x1_ASAP7_75t_R _14897_ (.A1(_07893_),
    .A2(_07894_),
    .B(net90),
    .Y(_07896_));
 OA21x2_ASAP7_75t_R _14898_ (.A1(_09700_),
    .A2(_07892_),
    .B(_07896_),
    .Y(_09721_));
 BUFx4f_ASAP7_75t_R _14899_ (.A(_07888_),
    .Y(_07897_));
 OR3x1_ASAP7_75t_R _14900_ (.A(_07070_),
    .B(_07071_),
    .C(_07897_),
    .Y(_07898_));
 OA21x2_ASAP7_75t_R _14901_ (.A1(net91),
    .A2(_07887_),
    .B(_07898_),
    .Y(_09723_));
 OR3x1_ASAP7_75t_R _14902_ (.A(_06392_),
    .B(_06417_),
    .C(_07897_),
    .Y(_07899_));
 OA21x2_ASAP7_75t_R _14903_ (.A1(net92),
    .A2(_07887_),
    .B(_07899_),
    .Y(_09725_));
 AO21x1_ASAP7_75t_R _14904_ (.A1(_07893_),
    .A2(_07894_),
    .B(net93),
    .Y(_07900_));
 OA21x2_ASAP7_75t_R _14905_ (.A1(_09685_),
    .A2(_07892_),
    .B(_07900_),
    .Y(_09727_));
 AO21x1_ASAP7_75t_R _14906_ (.A1(_07893_),
    .A2(_07894_),
    .B(net94),
    .Y(_07901_));
 OA21x2_ASAP7_75t_R _14907_ (.A1(_09680_),
    .A2(_07892_),
    .B(_07901_),
    .Y(_09729_));
 AO21x1_ASAP7_75t_R _14908_ (.A1(_07893_),
    .A2(_07894_),
    .B(net95),
    .Y(_07902_));
 OA21x2_ASAP7_75t_R _14909_ (.A1(_09675_),
    .A2(_07892_),
    .B(_07902_),
    .Y(_09731_));
 OR3x1_ASAP7_75t_R _14910_ (.A(_06030_),
    .B(_06050_),
    .C(_07897_),
    .Y(_07903_));
 OA21x2_ASAP7_75t_R _14911_ (.A1(net96),
    .A2(_07887_),
    .B(_07903_),
    .Y(_09733_));
 AO21x1_ASAP7_75t_R _14912_ (.A1(_07893_),
    .A2(_07894_),
    .B(net66),
    .Y(_07904_));
 OA21x2_ASAP7_75t_R _14913_ (.A1(_09665_),
    .A2(_07892_),
    .B(_07904_),
    .Y(_09735_));
 AO21x1_ASAP7_75t_R _14914_ (.A1(_07893_),
    .A2(_07894_),
    .B(net67),
    .Y(_07905_));
 OA21x2_ASAP7_75t_R _14915_ (.A1(_09660_),
    .A2(_07892_),
    .B(_07905_),
    .Y(_09737_));
 OR3x2_ASAP7_75t_R _14916_ (.A(_06908_),
    .B(_06909_),
    .C(_07897_),
    .Y(_07906_));
 OA21x2_ASAP7_75t_R _14917_ (.A1(net68),
    .A2(_07887_),
    .B(_07906_),
    .Y(_09739_));
 NAND2x1_ASAP7_75t_R _14918_ (.A(_09652_),
    .B(_07886_),
    .Y(_07907_));
 OA21x2_ASAP7_75t_R _14919_ (.A1(net69),
    .A2(_07887_),
    .B(_07907_),
    .Y(_09741_));
 AO21x1_ASAP7_75t_R _14920_ (.A1(_07893_),
    .A2(_07894_),
    .B(net70),
    .Y(_07908_));
 OA21x2_ASAP7_75t_R _14921_ (.A1(_09645_),
    .A2(_07892_),
    .B(_07908_),
    .Y(_09743_));
 OR3x1_ASAP7_75t_R _14922_ (.A(_05442_),
    .B(_05465_),
    .C(_07897_),
    .Y(_07909_));
 OA21x2_ASAP7_75t_R _14923_ (.A1(net71),
    .A2(_07887_),
    .B(_07909_),
    .Y(_09745_));
 OR3x1_ASAP7_75t_R _14924_ (.A(_05333_),
    .B(_05357_),
    .C(_07897_),
    .Y(_07910_));
 OA21x2_ASAP7_75t_R _14925_ (.A1(net72),
    .A2(_07887_),
    .B(_07910_),
    .Y(_09747_));
 OR3x1_ASAP7_75t_R _14926_ (.A(_06853_),
    .B(_06854_),
    .C(_07897_),
    .Y(_07911_));
 OA21x2_ASAP7_75t_R _14927_ (.A1(net73),
    .A2(_07887_),
    .B(_07911_),
    .Y(_09749_));
 AO21x1_ASAP7_75t_R _14928_ (.A1(_07893_),
    .A2(_07894_),
    .B(net74),
    .Y(_07912_));
 OA21x2_ASAP7_75t_R _14929_ (.A1(_09625_),
    .A2(_07892_),
    .B(_07912_),
    .Y(_09751_));
 AO21x1_ASAP7_75t_R _14930_ (.A1(_07893_),
    .A2(_07894_),
    .B(net75),
    .Y(_07913_));
 OA21x2_ASAP7_75t_R _14931_ (.A1(_09620_),
    .A2(_07892_),
    .B(_07913_),
    .Y(_09753_));
 AO21x1_ASAP7_75t_R _14932_ (.A1(_07882_),
    .A2(_07885_),
    .B(net77),
    .Y(_07914_));
 OA21x2_ASAP7_75t_R _14933_ (.A1(_09615_),
    .A2(_07889_),
    .B(_07914_),
    .Y(_09755_));
 AO21x1_ASAP7_75t_R _14934_ (.A1(_07882_),
    .A2(_07885_),
    .B(net78),
    .Y(_07915_));
 OA21x2_ASAP7_75t_R _14935_ (.A1(_09610_),
    .A2(_07889_),
    .B(_07915_),
    .Y(_09757_));
 AO21x1_ASAP7_75t_R _14936_ (.A1(_07882_),
    .A2(_07885_),
    .B(net79),
    .Y(_07916_));
 OA21x2_ASAP7_75t_R _14937_ (.A1(_09605_),
    .A2(_07889_),
    .B(_07916_),
    .Y(_09759_));
 AO21x1_ASAP7_75t_R _14938_ (.A1(_07882_),
    .A2(_07885_),
    .B(net80),
    .Y(_07917_));
 OA21x2_ASAP7_75t_R _14939_ (.A1(_09600_),
    .A2(_07889_),
    .B(_07917_),
    .Y(_09761_));
 AO21x1_ASAP7_75t_R _14940_ (.A1(_07882_),
    .A2(_07885_),
    .B(net81),
    .Y(_07918_));
 OA21x2_ASAP7_75t_R _14941_ (.A1(_09595_),
    .A2(_07889_),
    .B(_07918_),
    .Y(_09763_));
 OR3x2_ASAP7_75t_R _14942_ (.A(_04338_),
    .B(_04359_),
    .C(_07897_),
    .Y(_07919_));
 OA21x2_ASAP7_75t_R _14943_ (.A1(net82),
    .A2(_07886_),
    .B(_07919_),
    .Y(_09765_));
 OR3x1_ASAP7_75t_R _14944_ (.A(_04239_),
    .B(_04265_),
    .C(_07897_),
    .Y(_07920_));
 OA21x2_ASAP7_75t_R _14945_ (.A1(net83),
    .A2(_07886_),
    .B(_07920_),
    .Y(_09767_));
 AO21x1_ASAP7_75t_R _14946_ (.A1(_07882_),
    .A2(_07885_),
    .B(net84),
    .Y(_07921_));
 OA21x2_ASAP7_75t_R _14947_ (.A1(_09580_),
    .A2(_07889_),
    .B(_07921_),
    .Y(_09769_));
 AO21x1_ASAP7_75t_R _14948_ (.A1(_07882_),
    .A2(_07885_),
    .B(net85),
    .Y(_07922_));
 OA21x2_ASAP7_75t_R _14949_ (.A1(_09575_),
    .A2(_07889_),
    .B(_07922_),
    .Y(_09771_));
 OR3x1_ASAP7_75t_R _14950_ (.A(_03864_),
    .B(_03890_),
    .C(_07897_),
    .Y(_07923_));
 OA21x2_ASAP7_75t_R _14951_ (.A1(net86),
    .A2(_07886_),
    .B(_07923_),
    .Y(_09773_));
 AO21x1_ASAP7_75t_R _14952_ (.A1(_07882_),
    .A2(_07885_),
    .B(net88),
    .Y(_07924_));
 OA21x2_ASAP7_75t_R _14953_ (.A1(_09565_),
    .A2(_07889_),
    .B(_07924_),
    .Y(_09775_));
 NOR2x1_ASAP7_75t_R _14954_ (.A(_03281_),
    .B(_03292_),
    .Y(_09714_));
 NOR2x1_ASAP7_75t_R _14955_ (.A(_03779_),
    .B(_04878_),
    .Y(_09756_));
 NOR2x1_ASAP7_75t_R _14956_ (.A(_03779_),
    .B(_04765_),
    .Y(_09758_));
 NOR2x1_ASAP7_75t_R _14957_ (.A(_03779_),
    .B(_04658_),
    .Y(_09760_));
 NOR2x1_ASAP7_75t_R _14958_ (.A(_03779_),
    .B(_04546_),
    .Y(_09762_));
 NOR2x1_ASAP7_75t_R _14959_ (.A(_03779_),
    .B(_04424_),
    .Y(_09764_));
 INVx1_ASAP7_75t_R _14960_ (.A(_04162_),
    .Y(_09768_));
 OR3x1_ASAP7_75t_R _14961_ (.A(_03212_),
    .B(_05358_),
    .C(_06929_),
    .Y(_07925_));
 AO221x1_ASAP7_75t_R _14962_ (.A1(_04484_),
    .A2(_03774_),
    .B1(_03746_),
    .B2(_05032_),
    .C(_03706_),
    .Y(_07926_));
 AO32x1_ASAP7_75t_R _14963_ (.A1(_09570_),
    .A2(_03960_),
    .A3(_09575_),
    .B1(_09565_),
    .B2(_03706_),
    .Y(_07927_));
 AND2x2_ASAP7_75t_R _14964_ (.A(_03830_),
    .B(_07926_),
    .Y(_07928_));
 AO21x1_ASAP7_75t_R _14965_ (.A1(_03960_),
    .A2(_09575_),
    .B(_09570_),
    .Y(_07929_));
 XNOR2x1_ASAP7_75t_R _14966_ (.B(_03640_),
    .Y(_07930_),
    .A(_03554_));
 AOI221x1_ASAP7_75t_R _14967_ (.A1(_07926_),
    .A2(_07927_),
    .B1(_07928_),
    .B2(_07929_),
    .C(_07930_),
    .Y(_07931_));
 OR3x1_ASAP7_75t_R _14968_ (.A(_03864_),
    .B(_03890_),
    .C(_03960_),
    .Y(_07932_));
 OA21x2_ASAP7_75t_R _14969_ (.A1(_09575_),
    .A2(_07932_),
    .B(_07926_),
    .Y(_07933_));
 OR4x1_ASAP7_75t_R _14970_ (.A(_03781_),
    .B(_03829_),
    .C(_03864_),
    .D(_03890_),
    .Y(_07934_));
 OA31x2_ASAP7_75t_R _14971_ (.A1(_03830_),
    .A2(_03960_),
    .A3(_09575_),
    .B1(_07934_),
    .Y(_07935_));
 AOI22x1_ASAP7_75t_R _14972_ (.A1(_03706_),
    .A2(_09565_),
    .B1(_07933_),
    .B2(_07935_),
    .Y(_07936_));
 NOR2x1_ASAP7_75t_R _14973_ (.A(_03554_),
    .B(_03640_),
    .Y(_07937_));
 OA21x2_ASAP7_75t_R _14974_ (.A1(_03256_),
    .A2(_06942_),
    .B(_03640_),
    .Y(_07938_));
 AO32x2_ASAP7_75t_R _14975_ (.A1(_05775_),
    .A2(_05468_),
    .A3(_07937_),
    .B1(_07938_),
    .B2(_03554_),
    .Y(_07939_));
 AO21x2_ASAP7_75t_R _14976_ (.A1(_07931_),
    .A2(_07936_),
    .B(_07939_),
    .Y(_07940_));
 OR2x4_ASAP7_75t_R _14977_ (.A(_03127_),
    .B(_04210_),
    .Y(_07941_));
 NAND3x1_ASAP7_75t_R _14978_ (.A(_09580_),
    .B(_07941_),
    .C(_09585_),
    .Y(_07942_));
 OA211x2_ASAP7_75t_R _14979_ (.A1(_04239_),
    .A2(_04265_),
    .B(_04102_),
    .C(_07941_),
    .Y(_07943_));
 AOI21x1_ASAP7_75t_R _14980_ (.A1(_04102_),
    .A2(_09580_),
    .B(_07943_),
    .Y(_07944_));
 AND2x2_ASAP7_75t_R _14981_ (.A(_07942_),
    .B(_07944_),
    .Y(_07945_));
 NOR2x1_ASAP7_75t_R _14982_ (.A(_04163_),
    .B(_04312_),
    .Y(_07946_));
 AND2x2_ASAP7_75t_R _14983_ (.A(_07946_),
    .B(_09592_),
    .Y(_07947_));
 AOI22x1_ASAP7_75t_R _14984_ (.A1(_04313_),
    .A2(_09590_),
    .B1(_04421_),
    .B2(_09595_),
    .Y(_07948_));
 INVx1_ASAP7_75t_R _14985_ (.A(_04102_),
    .Y(_07949_));
 NOR3x1_ASAP7_75t_R _14986_ (.A(_07941_),
    .B(_04239_),
    .C(_04265_),
    .Y(_07950_));
 MAJx2_ASAP7_75t_R _14987_ (.A(_07949_),
    .B(_09582_),
    .C(_07950_),
    .Y(_07951_));
 OR3x1_ASAP7_75t_R _14988_ (.A(_07947_),
    .B(_07948_),
    .C(_07951_),
    .Y(_07952_));
 AND3x1_ASAP7_75t_R _14989_ (.A(_07931_),
    .B(_07945_),
    .C(_07952_),
    .Y(_07953_));
 NOR2x2_ASAP7_75t_R _14990_ (.A(_07940_),
    .B(_07953_),
    .Y(_07954_));
 AOI21x1_ASAP7_75t_R _14991_ (.A1(_07931_),
    .A2(_07936_),
    .B(_07939_),
    .Y(_07955_));
 AO21x1_ASAP7_75t_R _14992_ (.A1(_04656_),
    .A2(_09605_),
    .B(_09600_),
    .Y(_07956_));
 AO31x2_ASAP7_75t_R _14993_ (.A1(_09610_),
    .A2(_04877_),
    .A3(_09615_),
    .B(_04763_),
    .Y(_07957_));
 AO21x1_ASAP7_75t_R _14994_ (.A1(_04877_),
    .A2(_09615_),
    .B(_09610_),
    .Y(_07958_));
 AO32x1_ASAP7_75t_R _14995_ (.A1(_09600_),
    .A2(_04656_),
    .A3(_09605_),
    .B1(_04976_),
    .B2(_05033_),
    .Y(_07959_));
 AOI221x1_ASAP7_75t_R _14996_ (.A1(_04544_),
    .A2(_07956_),
    .B1(_07957_),
    .B2(_07958_),
    .C(_07959_),
    .Y(_07960_));
 AND2x2_ASAP7_75t_R _14997_ (.A(_05091_),
    .B(_09625_),
    .Y(_07961_));
 OAI21x1_ASAP7_75t_R _14998_ (.A1(_05278_),
    .A2(_05306_),
    .B(_03705_),
    .Y(_07962_));
 OA21x2_ASAP7_75t_R _14999_ (.A1(_05333_),
    .A2(_05357_),
    .B(_07962_),
    .Y(_07963_));
 MAJx2_ASAP7_75t_R _15000_ (.A(_05194_),
    .B(_09630_),
    .C(_07963_),
    .Y(_07964_));
 OA22x2_ASAP7_75t_R _15001_ (.A1(_04976_),
    .A2(_09620_),
    .B1(_05091_),
    .B2(_09625_),
    .Y(_07965_));
 OAI21x1_ASAP7_75t_R _15002_ (.A1(_07961_),
    .A2(_07964_),
    .B(_07965_),
    .Y(_07966_));
 OR2x2_ASAP7_75t_R _15003_ (.A(_04763_),
    .B(_09610_),
    .Y(_07967_));
 AO211x2_ASAP7_75t_R _15004_ (.A1(_04763_),
    .A2(_09610_),
    .B(_04877_),
    .C(_09615_),
    .Y(_07968_));
 AND2x2_ASAP7_75t_R _15005_ (.A(_04544_),
    .B(_09600_),
    .Y(_07969_));
 AOI221x1_ASAP7_75t_R _15006_ (.A1(_04656_),
    .A2(_09605_),
    .B1(_07967_),
    .B2(_07968_),
    .C(_07969_),
    .Y(_07970_));
 OR2x2_ASAP7_75t_R _15007_ (.A(_04656_),
    .B(_09605_),
    .Y(_07971_));
 OR2x2_ASAP7_75t_R _15008_ (.A(_04544_),
    .B(_09600_),
    .Y(_07972_));
 OAI21x1_ASAP7_75t_R _15009_ (.A1(_07969_),
    .A2(_07971_),
    .B(_07972_),
    .Y(_07973_));
 AOI211x1_ASAP7_75t_R _15010_ (.A1(_07960_),
    .A2(_07966_),
    .B(_07970_),
    .C(_07973_),
    .Y(_07974_));
 AOI221x1_ASAP7_75t_R _15011_ (.A1(_04439_),
    .A2(_04457_),
    .B1(_04483_),
    .B2(_06713_),
    .C(_04421_),
    .Y(_07975_));
 MAJx2_ASAP7_75t_R _15012_ (.A(_07946_),
    .B(_09592_),
    .C(_07975_),
    .Y(_07976_));
 AO31x2_ASAP7_75t_R _15013_ (.A1(_07942_),
    .A2(_07944_),
    .A3(_07976_),
    .B(_07951_),
    .Y(_07977_));
 NAND2x1_ASAP7_75t_R _15014_ (.A(_07931_),
    .B(_07977_),
    .Y(_07978_));
 AND3x2_ASAP7_75t_R _15015_ (.A(_07955_),
    .B(_07974_),
    .C(_07978_),
    .Y(_07979_));
 OR5x1_ASAP7_75t_R _15016_ (.A(_03213_),
    .B(_06927_),
    .C(_03217_),
    .D(_07954_),
    .E(_07979_),
    .Y(_07980_));
 NOR2x1_ASAP7_75t_R _15017_ (.A(_06191_),
    .B(_06236_),
    .Y(_07981_));
 AO21x1_ASAP7_75t_R _15018_ (.A1(_06499_),
    .A2(_06528_),
    .B(net125),
    .Y(_07982_));
 MAJx2_ASAP7_75t_R _15019_ (.A(net126),
    .B(_09692_),
    .C(_07982_),
    .Y(_07983_));
 MAJx2_ASAP7_75t_R _15020_ (.A(net127),
    .B(_09687_),
    .C(_07983_),
    .Y(_07984_));
 NAND2x2_ASAP7_75t_R _15021_ (.A(_06191_),
    .B(_06236_),
    .Y(_07985_));
 OA21x2_ASAP7_75t_R _15022_ (.A1(_07981_),
    .A2(_07984_),
    .B(_07985_),
    .Y(_07986_));
 AND2x2_ASAP7_75t_R _15023_ (.A(_06573_),
    .B(_06617_),
    .Y(_07987_));
 OR3x1_ASAP7_75t_R _15024_ (.A(_03176_),
    .B(_03427_),
    .C(_03496_),
    .Y(_07988_));
 MAJx2_ASAP7_75t_R _15025_ (.A(_06764_),
    .B(_09549_),
    .C(_07988_),
    .Y(_07989_));
 MAJx2_ASAP7_75t_R _15026_ (.A(_06670_),
    .B(_06714_),
    .C(_07989_),
    .Y(_07990_));
 OR2x2_ASAP7_75t_R _15027_ (.A(_06573_),
    .B(_09700_),
    .Y(_07991_));
 OAI21x1_ASAP7_75t_R _15028_ (.A1(_07987_),
    .A2(_07990_),
    .B(_07991_),
    .Y(_07992_));
 NAND2x1_ASAP7_75t_R _15029_ (.A(_06280_),
    .B(_09685_),
    .Y(_07993_));
 AND3x1_ASAP7_75t_R _15030_ (.A(net125),
    .B(_06499_),
    .C(_06528_),
    .Y(_07994_));
 MAJx2_ASAP7_75t_R _15031_ (.A(net126),
    .B(_09692_),
    .C(_07994_),
    .Y(_07995_));
 NOR2x1_ASAP7_75t_R _15032_ (.A(_06280_),
    .B(_09685_),
    .Y(_07996_));
 AO221x1_ASAP7_75t_R _15033_ (.A1(net128),
    .A2(_09682_),
    .B1(_07993_),
    .B2(_07995_),
    .C(_07996_),
    .Y(_07997_));
 AND2x2_ASAP7_75t_R _15034_ (.A(_05829_),
    .B(_05871_),
    .Y(_07998_));
 AO211x2_ASAP7_75t_R _15035_ (.A1(_04484_),
    .A2(_06118_),
    .B(_06145_),
    .C(_06094_),
    .Y(_07999_));
 MAJx2_ASAP7_75t_R _15036_ (.A(_06005_),
    .B(_09670_),
    .C(_07999_),
    .Y(_08000_));
 MAJx2_ASAP7_75t_R _15037_ (.A(_05917_),
    .B(_09665_),
    .C(_08000_),
    .Y(_08001_));
 OR2x2_ASAP7_75t_R _15038_ (.A(_05829_),
    .B(_09660_),
    .Y(_08002_));
 OAI21x1_ASAP7_75t_R _15039_ (.A1(_07998_),
    .A2(_08001_),
    .B(_08002_),
    .Y(_08003_));
 AO221x1_ASAP7_75t_R _15040_ (.A1(_07986_),
    .A2(_07992_),
    .B1(_07997_),
    .B2(_07985_),
    .C(_08003_),
    .Y(_08004_));
 AO21x1_ASAP7_75t_R _15041_ (.A1(_05743_),
    .A2(_05774_),
    .B(_05715_),
    .Y(_08005_));
 MAJx2_ASAP7_75t_R _15042_ (.A(_05610_),
    .B(_09652_),
    .C(_08005_),
    .Y(_08006_));
 MAJx2_ASAP7_75t_R _15043_ (.A(_05518_),
    .B(_09647_),
    .C(_08006_),
    .Y(_08007_));
 MAJx2_ASAP7_75t_R _15044_ (.A(_05417_),
    .B(_09642_),
    .C(_08007_),
    .Y(_08008_));
 OR2x2_ASAP7_75t_R _15045_ (.A(_05917_),
    .B(_09665_),
    .Y(_08009_));
 OA21x2_ASAP7_75t_R _15046_ (.A1(_07998_),
    .A2(_08009_),
    .B(_08002_),
    .Y(_08010_));
 OR2x2_ASAP7_75t_R _15047_ (.A(_06005_),
    .B(_09670_),
    .Y(_08011_));
 AO22x1_ASAP7_75t_R _15048_ (.A1(_06005_),
    .A2(_09670_),
    .B1(_06094_),
    .B2(_09675_),
    .Y(_08012_));
 AO221x1_ASAP7_75t_R _15049_ (.A1(_05917_),
    .A2(_09665_),
    .B1(_08011_),
    .B2(_08012_),
    .C(_07998_),
    .Y(_08013_));
 NAND2x1_ASAP7_75t_R _15050_ (.A(_08010_),
    .B(_08013_),
    .Y(_08014_));
 AND2x2_ASAP7_75t_R _15051_ (.A(_08008_),
    .B(_08014_),
    .Y(_08015_));
 AND3x1_ASAP7_75t_R _15052_ (.A(_05715_),
    .B(_05743_),
    .C(_05774_),
    .Y(_08016_));
 MAJx2_ASAP7_75t_R _15053_ (.A(_05610_),
    .B(_09652_),
    .C(_08016_),
    .Y(_08017_));
 MAJx2_ASAP7_75t_R _15054_ (.A(_05518_),
    .B(_09647_),
    .C(_08017_),
    .Y(_08018_));
 MAJx3_ASAP7_75t_R _15055_ (.A(_05417_),
    .B(_09642_),
    .C(_08018_),
    .Y(_08019_));
 AOI21x1_ASAP7_75t_R _15056_ (.A1(_08004_),
    .A2(_08015_),
    .B(_08019_),
    .Y(_08020_));
 AO21x2_ASAP7_75t_R _15057_ (.A1(_07925_),
    .A2(_07980_),
    .B(_08020_),
    .Y(_08021_));
 NOR2x2_ASAP7_75t_R _15058_ (.A(_07954_),
    .B(_07979_),
    .Y(_08022_));
 NAND2x1_ASAP7_75t_R _15059_ (.A(_07985_),
    .B(_07997_),
    .Y(_08023_));
 OA211x2_ASAP7_75t_R _15060_ (.A1(_06764_),
    .A2(_09549_),
    .B(_03176_),
    .C(_09555_),
    .Y(_08024_));
 OAI21x1_ASAP7_75t_R _15061_ (.A1(_06670_),
    .A2(_09705_),
    .B(_08024_),
    .Y(_08025_));
 OA211x2_ASAP7_75t_R _15062_ (.A1(_06670_),
    .A2(_06714_),
    .B(_06764_),
    .C(_09549_),
    .Y(_08026_));
 AOI211x1_ASAP7_75t_R _15063_ (.A1(_06670_),
    .A2(_06714_),
    .B(_07987_),
    .C(_08026_),
    .Y(_08027_));
 AOI22x1_ASAP7_75t_R _15064_ (.A1(net124),
    .A2(_09702_),
    .B1(_08025_),
    .B2(_08027_),
    .Y(_08028_));
 OAI21x1_ASAP7_75t_R _15065_ (.A1(_07981_),
    .A2(_07984_),
    .B(_07985_),
    .Y(_08029_));
 AO221x1_ASAP7_75t_R _15066_ (.A1(_08010_),
    .A2(_08013_),
    .B1(_08023_),
    .B2(_08028_),
    .C(_08029_),
    .Y(_08030_));
 NOR2x1_ASAP7_75t_R _15067_ (.A(_08019_),
    .B(_08003_),
    .Y(_08031_));
 AO211x2_ASAP7_75t_R _15068_ (.A1(_05338_),
    .A2(_05343_),
    .B(_05356_),
    .C(_03426_),
    .Y(_08032_));
 OA31x2_ASAP7_75t_R _15069_ (.A1(_04003_),
    .A2(_05320_),
    .A3(_05332_),
    .B1(_05307_),
    .Y(_08033_));
 NAND2x1_ASAP7_75t_R _15070_ (.A(_08032_),
    .B(_08033_),
    .Y(_08034_));
 OA222x2_ASAP7_75t_R _15071_ (.A1(_05091_),
    .A2(_09625_),
    .B1(_09630_),
    .B2(_08034_),
    .C1(_05193_),
    .C2(_04163_),
    .Y(_08035_));
 AOI22x1_ASAP7_75t_R _15072_ (.A1(_05224_),
    .A2(_05247_),
    .B1(_08032_),
    .B2(_08033_),
    .Y(_08036_));
 MAJx2_ASAP7_75t_R _15073_ (.A(_05091_),
    .B(_05146_),
    .C(_08036_),
    .Y(_08037_));
 OR2x2_ASAP7_75t_R _15074_ (.A(_04976_),
    .B(_09620_),
    .Y(_08038_));
 OAI21x1_ASAP7_75t_R _15075_ (.A1(_08035_),
    .A2(_08037_),
    .B(_08038_),
    .Y(_08039_));
 AO211x2_ASAP7_75t_R _15076_ (.A1(_07960_),
    .A2(_08039_),
    .B(_07970_),
    .C(_07973_),
    .Y(_08040_));
 OA211x2_ASAP7_75t_R _15077_ (.A1(_07939_),
    .A2(_07931_),
    .B(_07945_),
    .C(_07952_),
    .Y(_08041_));
 AND2x2_ASAP7_75t_R _15078_ (.A(_07931_),
    .B(_07977_),
    .Y(_08042_));
 AO211x2_ASAP7_75t_R _15079_ (.A1(_08040_),
    .A2(_08041_),
    .B(_07940_),
    .C(_08042_),
    .Y(_08043_));
 INVx1_ASAP7_75t_R _15080_ (.A(_08008_),
    .Y(_08044_));
 AOI211x1_ASAP7_75t_R _15081_ (.A1(_08030_),
    .A2(_08031_),
    .B(_08043_),
    .C(_08044_),
    .Y(_08045_));
 NAND2x1_ASAP7_75t_R _15082_ (.A(_06826_),
    .B(_06928_),
    .Y(_08046_));
 AO21x1_ASAP7_75t_R _15083_ (.A1(_08004_),
    .A2(_08015_),
    .B(_08019_),
    .Y(_08047_));
 AO211x2_ASAP7_75t_R _15084_ (.A1(_08022_),
    .A2(_08045_),
    .B(_08046_),
    .C(_08047_),
    .Y(_08048_));
 AND2x2_ASAP7_75t_R _15085_ (.A(_03024_),
    .B(_03217_),
    .Y(_08049_));
 OA21x2_ASAP7_75t_R _15086_ (.A1(_03212_),
    .A2(_05358_),
    .B(_03024_),
    .Y(_08050_));
 AO21x1_ASAP7_75t_R _15087_ (.A1(_08030_),
    .A2(_08031_),
    .B(_08044_),
    .Y(_08051_));
 OR3x1_ASAP7_75t_R _15088_ (.A(_07954_),
    .B(_07979_),
    .C(_08043_),
    .Y(_08052_));
 OR5x2_ASAP7_75t_R _15089_ (.A(_08049_),
    .B(_08047_),
    .C(_08050_),
    .D(_08051_),
    .E(_08052_),
    .Y(_08053_));
 AND3x2_ASAP7_75t_R _15090_ (.A(_08021_),
    .B(_08048_),
    .C(_08053_),
    .Y(_08054_));
 BUFx4f_ASAP7_75t_R _15091_ (.A(_08054_),
    .Y(_08055_));
 OR4x1_ASAP7_75t_R _15092_ (.A(_08019_),
    .B(_07940_),
    .C(_08042_),
    .D(_08040_),
    .Y(_08056_));
 AO21x2_ASAP7_75t_R _15093_ (.A1(_08004_),
    .A2(_08015_),
    .B(_08056_),
    .Y(_08057_));
 AND3x4_ASAP7_75t_R _15094_ (.A(_07000_),
    .B(_08022_),
    .C(_08057_),
    .Y(_08058_));
 AND3x1_ASAP7_75t_R _15095_ (.A(_03024_),
    .B(_05358_),
    .C(_03217_),
    .Y(_08059_));
 AOI21x1_ASAP7_75t_R _15096_ (.A1(_08022_),
    .A2(_08057_),
    .B(_08059_),
    .Y(_08060_));
 OR2x2_ASAP7_75t_R _15097_ (.A(_08058_),
    .B(_08060_),
    .Y(_08061_));
 BUFx4f_ASAP7_75t_R _15098_ (.A(_08061_),
    .Y(_08062_));
 BUFx4f_ASAP7_75t_R _15099_ (.A(_03256_),
    .Y(_08063_));
 AO21x2_ASAP7_75t_R _15100_ (.A1(_08055_),
    .A2(_08062_),
    .B(_08063_),
    .Y(_08064_));
 AND3x2_ASAP7_75t_R _15101_ (.A(_05775_),
    .B(_05468_),
    .C(_06930_),
    .Y(_08065_));
 AOI21x1_ASAP7_75t_R _15102_ (.A1(_08043_),
    .A2(_08065_),
    .B(_05467_),
    .Y(_08066_));
 BUFx4f_ASAP7_75t_R _15103_ (.A(_08066_),
    .Y(_08067_));
 BUFx4f_ASAP7_75t_R _15104_ (.A(_08067_),
    .Y(_08068_));
 NAND2x2_ASAP7_75t_R _15105_ (.A(_08064_),
    .B(_08068_),
    .Y(_08069_));
 BUFx4f_ASAP7_75t_R _15106_ (.A(_08069_),
    .Y(_08070_));
 BUFx3_ASAP7_75t_R _15107_ (.A(_08064_),
    .Y(_08071_));
 BUFx3_ASAP7_75t_R _15108_ (.A(_08068_),
    .Y(_08072_));
 INVx1_ASAP7_75t_R _15109_ (.A(_01067_),
    .Y(_08073_));
 AO21x1_ASAP7_75t_R _15110_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08073_),
    .Y(_08074_));
 OA21x2_ASAP7_75t_R _15111_ (.A1(net65),
    .A2(_08070_),
    .B(_08074_),
    .Y(_01220_));
 INVx1_ASAP7_75t_R _15112_ (.A(_01070_),
    .Y(_08075_));
 AO21x1_ASAP7_75t_R _15113_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08075_),
    .Y(_08076_));
 OA21x2_ASAP7_75t_R _15114_ (.A1(net76),
    .A2(_08070_),
    .B(_08076_),
    .Y(_01221_));
 INVx1_ASAP7_75t_R _15115_ (.A(_00732_),
    .Y(_01223_));
 INVx1_ASAP7_75t_R _15116_ (.A(_00699_),
    .Y(_01224_));
 INVx1_ASAP7_75t_R _15117_ (.A(_00633_),
    .Y(_01226_));
 INVx1_ASAP7_75t_R _15118_ (.A(_00600_),
    .Y(_01227_));
 INVx1_ASAP7_75t_R _15119_ (.A(_00566_),
    .Y(_01228_));
 INVx1_ASAP7_75t_R _15120_ (.A(_00467_),
    .Y(_01231_));
 INVx1_ASAP7_75t_R _15121_ (.A(_00434_),
    .Y(_01232_));
 INVx1_ASAP7_75t_R _15122_ (.A(_01032_),
    .Y(_01233_));
 INVx1_ASAP7_75t_R _15123_ (.A(_00401_),
    .Y(_01234_));
 INVx1_ASAP7_75t_R _15124_ (.A(_00368_),
    .Y(_01235_));
 INVx1_ASAP7_75t_R _15125_ (.A(_00335_),
    .Y(_01236_));
 INVx1_ASAP7_75t_R _15126_ (.A(_00301_),
    .Y(_01237_));
 INVx1_ASAP7_75t_R _15127_ (.A(_00201_),
    .Y(_01240_));
 INVx1_ASAP7_75t_R _15128_ (.A(_00168_),
    .Y(_01241_));
 INVx1_ASAP7_75t_R _15129_ (.A(_00134_),
    .Y(_01242_));
 INVx1_ASAP7_75t_R _15130_ (.A(_00101_),
    .Y(_01243_));
 INVx1_ASAP7_75t_R _15131_ (.A(_00999_),
    .Y(_01244_));
 INVx1_ASAP7_75t_R _15132_ (.A(_00067_),
    .Y(_01245_));
 INVx1_ASAP7_75t_R _15133_ (.A(_00966_),
    .Y(_01247_));
 INVx1_ASAP7_75t_R _15134_ (.A(_00899_),
    .Y(_01249_));
 INVx1_ASAP7_75t_R _15135_ (.A(_00866_),
    .Y(_01250_));
 INVx1_ASAP7_75t_R _15136_ (.A(_00832_),
    .Y(_01251_));
 INVx1_ASAP7_75t_R _15137_ (.A(_00799_),
    .Y(_01252_));
 INVx1_ASAP7_75t_R _15138_ (.A(_00765_),
    .Y(_01253_));
 NAND3x2_ASAP7_75t_R _15139_ (.B(_08048_),
    .C(_08053_),
    .Y(_08077_),
    .A(_08021_));
 BUFx3_ASAP7_75t_R _15140_ (.A(_08077_),
    .Y(_08078_));
 NOR2x2_ASAP7_75t_R _15141_ (.A(_08058_),
    .B(_08060_),
    .Y(_08079_));
 BUFx3_ASAP7_75t_R _15142_ (.A(_08079_),
    .Y(_08080_));
 AO21x2_ASAP7_75t_R _15143_ (.A1(_08043_),
    .A2(_08065_),
    .B(_05467_),
    .Y(_08081_));
 BUFx4f_ASAP7_75t_R _15144_ (.A(_08081_),
    .Y(_08082_));
 OR4x1_ASAP7_75t_R _15145_ (.A(_08073_),
    .B(_08078_),
    .C(_08080_),
    .D(_08082_),
    .Y(_08083_));
 BUFx4f_ASAP7_75t_R _15146_ (.A(_08077_),
    .Y(_08084_));
 AND2x2_ASAP7_75t_R _15147_ (.A(_01066_),
    .B(_05777_),
    .Y(_08085_));
 NAND2x1_ASAP7_75t_R _15148_ (.A(_08084_),
    .B(_08085_),
    .Y(_08086_));
 BUFx4f_ASAP7_75t_R _15149_ (.A(_08079_),
    .Y(_08087_));
 BUFx4f_ASAP7_75t_R _15150_ (.A(_08066_),
    .Y(_08088_));
 BUFx3_ASAP7_75t_R _15151_ (.A(_08088_),
    .Y(_08089_));
 AND3x1_ASAP7_75t_R _15152_ (.A(_01067_),
    .B(_08063_),
    .C(_08089_),
    .Y(_08090_));
 AOI221x1_ASAP7_75t_R _15153_ (.A1(_01066_),
    .A2(_08082_),
    .B1(_08085_),
    .B2(_08087_),
    .C(_08090_),
    .Y(_08091_));
 AND3x4_ASAP7_75t_R _15154_ (.A(_08083_),
    .B(_08086_),
    .C(_08091_),
    .Y(_08092_));
 BUFx4f_ASAP7_75t_R _15155_ (.A(_08092_),
    .Y(_08093_));
 AOI21x1_ASAP7_75t_R _15156_ (.A1(_03025_),
    .A2(net28),
    .B(_03278_),
    .Y(_08094_));
 INVx1_ASAP7_75t_R _15157_ (.A(_03269_),
    .Y(_08095_));
 OR3x4_ASAP7_75t_R _15158_ (.A(_06926_),
    .B(_03222_),
    .C(_08095_),
    .Y(_08096_));
 AND3x4_ASAP7_75t_R _15159_ (.A(_08094_),
    .B(_06715_),
    .C(_08096_),
    .Y(_08097_));
 BUFx16f_ASAP7_75t_R _15160_ (.A(_08097_),
    .Y(_08098_));
 INVx1_ASAP7_75t_R _15161_ (.A(net5),
    .Y(_08099_));
 AOI21x1_ASAP7_75t_R _15162_ (.A1(_03024_),
    .A2(net30),
    .B(_03238_),
    .Y(_08100_));
 AND4x2_ASAP7_75t_R _15163_ (.A(_03025_),
    .B(_08099_),
    .C(net2),
    .D(_08100_),
    .Y(_08101_));
 BUFx16f_ASAP7_75t_R _15164_ (.A(_08101_),
    .Y(_08102_));
 AND2x6_ASAP7_75t_R _15165_ (.A(_08098_),
    .B(_08102_),
    .Y(_08103_));
 INVx2_ASAP7_75t_R _15166_ (.A(_05467_),
    .Y(_08104_));
 NAND2x2_ASAP7_75t_R _15167_ (.A(_08104_),
    .B(_07884_),
    .Y(_08105_));
 BUFx16f_ASAP7_75t_R _15168_ (.A(_08105_),
    .Y(_08106_));
 NAND2x2_ASAP7_75t_R _15169_ (.A(_08103_),
    .B(_08106_),
    .Y(_08107_));
 BUFx4f_ASAP7_75t_R _15170_ (.A(_06935_),
    .Y(_08108_));
 AND3x1_ASAP7_75t_R _15171_ (.A(\readdata[0] ),
    .B(_03222_),
    .C(_03224_),
    .Y(_08109_));
 AO21x2_ASAP7_75t_R _15172_ (.A1(_08108_),
    .A2(net32),
    .B(_08109_),
    .Y(_08110_));
 BUFx6f_ASAP7_75t_R _15173_ (.A(_08110_),
    .Y(_08111_));
 AND2x4_ASAP7_75t_R _15174_ (.A(_08104_),
    .B(_07884_),
    .Y(_08112_));
 BUFx16f_ASAP7_75t_R _15175_ (.A(_08112_),
    .Y(_08113_));
 BUFx16f_ASAP7_75t_R _15176_ (.A(_08113_),
    .Y(_08114_));
 BUFx16f_ASAP7_75t_R _15177_ (.A(_08114_),
    .Y(_08115_));
 NAND2x2_ASAP7_75t_R _15178_ (.A(_08103_),
    .B(_08115_),
    .Y(_08116_));
 BUFx12f_ASAP7_75t_R _15179_ (.A(_08097_),
    .Y(_08117_));
 NAND2x2_ASAP7_75t_R _15180_ (.A(_08117_),
    .B(_08102_),
    .Y(_08118_));
 NAND2x1_ASAP7_75t_R _15181_ (.A(_00010_),
    .B(_08118_),
    .Y(_08119_));
 OA21x2_ASAP7_75t_R _15182_ (.A1(_08111_),
    .A2(_08116_),
    .B(_08119_),
    .Y(_08120_));
 OA21x2_ASAP7_75t_R _15183_ (.A1(_08093_),
    .A2(_08107_),
    .B(_08120_),
    .Y(_01254_));
 BUFx6f_ASAP7_75t_R _15184_ (.A(_08107_),
    .Y(_08121_));
 OR4x2_ASAP7_75t_R _15185_ (.A(_01081_),
    .B(_01084_),
    .C(_01087_),
    .D(_01090_),
    .Y(_08122_));
 OR3x4_ASAP7_75t_R _15186_ (.A(_01075_),
    .B(_01078_),
    .C(_01218_),
    .Y(_08123_));
 OR2x2_ASAP7_75t_R _15187_ (.A(_08122_),
    .B(_08123_),
    .Y(_08124_));
 BUFx4f_ASAP7_75t_R _15188_ (.A(_08124_),
    .Y(_08125_));
 XNOR2x1_ASAP7_75t_R _15189_ (.B(_08125_),
    .Y(_08126_),
    .A(net66));
 AND2x2_ASAP7_75t_R _15190_ (.A(_05777_),
    .B(_08126_),
    .Y(_08127_));
 AND2x2_ASAP7_75t_R _15191_ (.A(_08084_),
    .B(_08127_),
    .Y(_08128_));
 OA21x2_ASAP7_75t_R _15192_ (.A1(_01071_),
    .A2(_01159_),
    .B(_01074_),
    .Y(_08129_));
 OA21x2_ASAP7_75t_R _15193_ (.A1(_01073_),
    .A2(_08129_),
    .B(_01077_),
    .Y(_08130_));
 OA21x2_ASAP7_75t_R _15194_ (.A1(_01076_),
    .A2(_08130_),
    .B(_01080_),
    .Y(_08131_));
 OR2x2_ASAP7_75t_R _15195_ (.A(_01079_),
    .B(_01082_),
    .Y(_08132_));
 OA21x2_ASAP7_75t_R _15196_ (.A1(_01083_),
    .A2(_01082_),
    .B(_01086_),
    .Y(_08133_));
 OA21x2_ASAP7_75t_R _15197_ (.A1(_08131_),
    .A2(_08132_),
    .B(_08133_),
    .Y(_08134_));
 OA21x2_ASAP7_75t_R _15198_ (.A1(_01085_),
    .A2(_08134_),
    .B(_01089_),
    .Y(_08135_));
 OA21x2_ASAP7_75t_R _15199_ (.A1(_01088_),
    .A2(_08135_),
    .B(_01092_),
    .Y(_08136_));
 OA21x2_ASAP7_75t_R _15200_ (.A1(_01091_),
    .A2(_08136_),
    .B(_01095_),
    .Y(_08137_));
 XOR2x1_ASAP7_75t_R _15201_ (.A(_01094_),
    .Y(_08138_),
    .B(_08137_));
 AND4x1_ASAP7_75t_R _15202_ (.A(_08055_),
    .B(_08062_),
    .C(_08068_),
    .D(_08138_),
    .Y(_08139_));
 BUFx3_ASAP7_75t_R _15203_ (.A(_08088_),
    .Y(_08140_));
 AND3x1_ASAP7_75t_R _15204_ (.A(_08063_),
    .B(_08140_),
    .C(_08138_),
    .Y(_08141_));
 AO221x1_ASAP7_75t_R _15205_ (.A1(_08082_),
    .A2(_08126_),
    .B1(_08127_),
    .B2(_08087_),
    .C(_08141_),
    .Y(_08142_));
 OR3x4_ASAP7_75t_R _15206_ (.A(_08128_),
    .B(_08139_),
    .C(_08142_),
    .Y(_08143_));
 BUFx12_ASAP7_75t_R _15207_ (.A(_08118_),
    .Y(_08144_));
 BUFx6f_ASAP7_75t_R _15208_ (.A(_08098_),
    .Y(_08145_));
 BUFx6f_ASAP7_75t_R _15209_ (.A(_08102_),
    .Y(_08146_));
 AND3x2_ASAP7_75t_R _15210_ (.A(_08145_),
    .B(_08146_),
    .C(_08113_),
    .Y(_08147_));
 BUFx10_ASAP7_75t_R _15211_ (.A(_08147_),
    .Y(_08148_));
 AND2x4_ASAP7_75t_R _15212_ (.A(_03222_),
    .B(_03224_),
    .Y(_08149_));
 BUFx6f_ASAP7_75t_R _15213_ (.A(_08149_),
    .Y(_08150_));
 OR3x4_ASAP7_75t_R _15214_ (.A(_08049_),
    .B(_06935_),
    .C(_05468_),
    .Y(_08151_));
 AND5x2_ASAP7_75t_R _15215_ (.A(\readdata[7] ),
    .B(_03218_),
    .C(_08149_),
    .D(_06942_),
    .E(_07000_),
    .Y(_08152_));
 AO21x1_ASAP7_75t_R _15216_ (.A1(\readdata[10] ),
    .A2(_08151_),
    .B(_08152_),
    .Y(_08153_));
 OR2x2_ASAP7_75t_R _15217_ (.A(_06935_),
    .B(_08153_),
    .Y(_08154_));
 OAI21x1_ASAP7_75t_R _15218_ (.A1(_08150_),
    .A2(net33),
    .B(_08154_),
    .Y(_08155_));
 BUFx6f_ASAP7_75t_R _15219_ (.A(_08155_),
    .Y(_08156_));
 AOI22x1_ASAP7_75t_R _15220_ (.A1(_00742_),
    .A2(_08144_),
    .B1(_08148_),
    .B2(_08156_),
    .Y(_08157_));
 OA21x2_ASAP7_75t_R _15221_ (.A1(_08121_),
    .A2(_08143_),
    .B(_08157_),
    .Y(_01255_));
 OR3x2_ASAP7_75t_R _15222_ (.A(_09717_),
    .B(_09718_),
    .C(_01075_),
    .Y(_08158_));
 OR2x2_ASAP7_75t_R _15223_ (.A(_01078_),
    .B(_08158_),
    .Y(_08159_));
 OR3x1_ASAP7_75t_R _15224_ (.A(_01093_),
    .B(_08122_),
    .C(_08159_),
    .Y(_08160_));
 XNOR2x1_ASAP7_75t_R _15225_ (.B(_08160_),
    .Y(_08161_),
    .A(net67));
 AND2x2_ASAP7_75t_R _15226_ (.A(_05777_),
    .B(_08161_),
    .Y(_08162_));
 AND2x2_ASAP7_75t_R _15227_ (.A(_08084_),
    .B(_08162_),
    .Y(_08163_));
 OA21x2_ASAP7_75t_R _15228_ (.A1(_01069_),
    .A2(_09554_),
    .B(_01072_),
    .Y(_08164_));
 OA21x2_ASAP7_75t_R _15229_ (.A1(_01071_),
    .A2(_08164_),
    .B(_01074_),
    .Y(_08165_));
 OR2x2_ASAP7_75t_R _15230_ (.A(_01073_),
    .B(_01076_),
    .Y(_08166_));
 OA21x2_ASAP7_75t_R _15231_ (.A1(_01077_),
    .A2(_01076_),
    .B(_01080_),
    .Y(_08167_));
 OA21x2_ASAP7_75t_R _15232_ (.A1(_08165_),
    .A2(_08166_),
    .B(_08167_),
    .Y(_08168_));
 OA21x2_ASAP7_75t_R _15233_ (.A1(_08132_),
    .A2(_08168_),
    .B(_08133_),
    .Y(_08169_));
 OA21x2_ASAP7_75t_R _15234_ (.A1(_01085_),
    .A2(_08169_),
    .B(_01089_),
    .Y(_08170_));
 OA21x2_ASAP7_75t_R _15235_ (.A1(_01088_),
    .A2(_08170_),
    .B(_01092_),
    .Y(_08171_));
 OA21x2_ASAP7_75t_R _15236_ (.A1(_01091_),
    .A2(_08171_),
    .B(_01095_),
    .Y(_08172_));
 OA21x2_ASAP7_75t_R _15237_ (.A1(_01094_),
    .A2(_08172_),
    .B(_01098_),
    .Y(_08173_));
 XOR2x1_ASAP7_75t_R _15238_ (.A(_01097_),
    .Y(_08174_),
    .B(_08173_));
 AND4x1_ASAP7_75t_R _15239_ (.A(_08055_),
    .B(_08062_),
    .C(_08068_),
    .D(_08174_),
    .Y(_08175_));
 AND3x1_ASAP7_75t_R _15240_ (.A(_08063_),
    .B(_08140_),
    .C(_08174_),
    .Y(_08176_));
 AO221x1_ASAP7_75t_R _15241_ (.A1(_08082_),
    .A2(_08161_),
    .B1(_08162_),
    .B2(_08087_),
    .C(_08176_),
    .Y(_08177_));
 OR3x4_ASAP7_75t_R _15242_ (.A(_08163_),
    .B(_08175_),
    .C(_08177_),
    .Y(_08178_));
 BUFx4f_ASAP7_75t_R _15243_ (.A(_08151_),
    .Y(_08179_));
 AND4x1_ASAP7_75t_R _15244_ (.A(\readdata[7] ),
    .B(_03218_),
    .C(_06942_),
    .D(_07000_),
    .Y(_08180_));
 OR2x2_ASAP7_75t_R _15245_ (.A(_06935_),
    .B(_08180_),
    .Y(_08181_));
 BUFx3_ASAP7_75t_R _15246_ (.A(_08181_),
    .Y(_08182_));
 AO21x1_ASAP7_75t_R _15247_ (.A1(\readdata[11] ),
    .A2(_08179_),
    .B(_08182_),
    .Y(_08183_));
 OAI21x1_ASAP7_75t_R _15248_ (.A1(_08150_),
    .A2(net34),
    .B(_08183_),
    .Y(_08184_));
 BUFx10_ASAP7_75t_R _15249_ (.A(_08184_),
    .Y(_08185_));
 AOI22x1_ASAP7_75t_R _15250_ (.A1(_00709_),
    .A2(_08144_),
    .B1(_08148_),
    .B2(_08185_),
    .Y(_08186_));
 OA21x2_ASAP7_75t_R _15251_ (.A1(_08121_),
    .A2(_08178_),
    .B(_08186_),
    .Y(_01256_));
 INVx1_ASAP7_75t_R _15252_ (.A(_00676_),
    .Y(_08187_));
 BUFx3_ASAP7_75t_R _15253_ (.A(_08151_),
    .Y(_08188_));
 AO21x1_ASAP7_75t_R _15254_ (.A1(\readdata[12] ),
    .A2(_08188_),
    .B(_08182_),
    .Y(_08189_));
 OA21x2_ASAP7_75t_R _15255_ (.A1(_08150_),
    .A2(net35),
    .B(_08189_),
    .Y(_08190_));
 BUFx4f_ASAP7_75t_R _15256_ (.A(_08190_),
    .Y(_08191_));
 OR3x1_ASAP7_75t_R _15257_ (.A(_01093_),
    .B(_01096_),
    .C(_08125_),
    .Y(_08192_));
 XNOR2x1_ASAP7_75t_R _15258_ (.B(_08192_),
    .Y(_08193_),
    .A(net68));
 AND2x2_ASAP7_75t_R _15259_ (.A(_05776_),
    .B(_08193_),
    .Y(_08194_));
 AND2x2_ASAP7_75t_R _15260_ (.A(_08078_),
    .B(_08194_),
    .Y(_08195_));
 BUFx6f_ASAP7_75t_R _15261_ (.A(_08054_),
    .Y(_08196_));
 BUFx3_ASAP7_75t_R _15262_ (.A(_08061_),
    .Y(_08197_));
 OA21x2_ASAP7_75t_R _15263_ (.A1(_01094_),
    .A2(_08137_),
    .B(_01098_),
    .Y(_08198_));
 OA21x2_ASAP7_75t_R _15264_ (.A1(_01097_),
    .A2(_08198_),
    .B(_01101_),
    .Y(_08199_));
 XOR2x1_ASAP7_75t_R _15265_ (.A(_01100_),
    .Y(_08200_),
    .B(_08199_));
 AND4x1_ASAP7_75t_R _15266_ (.A(_08196_),
    .B(_08197_),
    .C(_08140_),
    .D(_08200_),
    .Y(_08201_));
 BUFx3_ASAP7_75t_R _15267_ (.A(_08081_),
    .Y(_08202_));
 BUFx4f_ASAP7_75t_R _15268_ (.A(_03256_),
    .Y(_08203_));
 AND3x1_ASAP7_75t_R _15269_ (.A(_08203_),
    .B(_08067_),
    .C(_08200_),
    .Y(_08204_));
 AO221x1_ASAP7_75t_R _15270_ (.A1(_08202_),
    .A2(_08193_),
    .B1(_08194_),
    .B2(_08080_),
    .C(_08204_),
    .Y(_08205_));
 OR3x4_ASAP7_75t_R _15271_ (.A(_08195_),
    .B(_08201_),
    .C(_08205_),
    .Y(_08206_));
 OA222x2_ASAP7_75t_R _15272_ (.A1(_08187_),
    .A2(_08103_),
    .B1(_08116_),
    .B2(_08191_),
    .C1(_08206_),
    .C2(_08107_),
    .Y(_01257_));
 INVx1_ASAP7_75t_R _15273_ (.A(_00643_),
    .Y(_08207_));
 AO21x1_ASAP7_75t_R _15274_ (.A1(\readdata[13] ),
    .A2(_08179_),
    .B(_08152_),
    .Y(_08208_));
 AND2x2_ASAP7_75t_R _15275_ (.A(_08149_),
    .B(_08208_),
    .Y(_08209_));
 AO21x2_ASAP7_75t_R _15276_ (.A1(_08108_),
    .A2(net36),
    .B(_08209_),
    .Y(_08210_));
 BUFx3_ASAP7_75t_R _15277_ (.A(_08210_),
    .Y(_08211_));
 OR3x1_ASAP7_75t_R _15278_ (.A(_01078_),
    .B(_08122_),
    .C(_08158_),
    .Y(_08212_));
 BUFx4f_ASAP7_75t_R _15279_ (.A(_08212_),
    .Y(_08213_));
 OR4x1_ASAP7_75t_R _15280_ (.A(_01093_),
    .B(_01096_),
    .C(_01099_),
    .D(_08213_),
    .Y(_08214_));
 XNOR2x1_ASAP7_75t_R _15281_ (.B(_08214_),
    .Y(_08215_),
    .A(net69));
 AND2x2_ASAP7_75t_R _15282_ (.A(_05776_),
    .B(_08215_),
    .Y(_08216_));
 AND2x2_ASAP7_75t_R _15283_ (.A(_08078_),
    .B(_08216_),
    .Y(_08217_));
 OA21x2_ASAP7_75t_R _15284_ (.A1(_01097_),
    .A2(_08173_),
    .B(_01101_),
    .Y(_08218_));
 OA21x2_ASAP7_75t_R _15285_ (.A1(_01100_),
    .A2(_08218_),
    .B(_01104_),
    .Y(_08219_));
 XOR2x1_ASAP7_75t_R _15286_ (.A(_01103_),
    .Y(_08220_),
    .B(_08219_));
 AND4x1_ASAP7_75t_R _15287_ (.A(_08196_),
    .B(_08197_),
    .C(_08140_),
    .D(_08220_),
    .Y(_08221_));
 AND3x1_ASAP7_75t_R _15288_ (.A(_08203_),
    .B(_08088_),
    .C(_08220_),
    .Y(_08222_));
 AO221x1_ASAP7_75t_R _15289_ (.A1(_08202_),
    .A2(_08215_),
    .B1(_08216_),
    .B2(_08080_),
    .C(_08222_),
    .Y(_08223_));
 OR3x4_ASAP7_75t_R _15290_ (.A(_08217_),
    .B(_08221_),
    .C(_08223_),
    .Y(_08224_));
 OA222x2_ASAP7_75t_R _15291_ (.A1(_08207_),
    .A2(_08103_),
    .B1(_08116_),
    .B2(_08211_),
    .C1(_08224_),
    .C2(_08107_),
    .Y(_01258_));
 OR4x1_ASAP7_75t_R _15292_ (.A(_01093_),
    .B(_01096_),
    .C(_01099_),
    .D(_01102_),
    .Y(_08225_));
 OR3x1_ASAP7_75t_R _15293_ (.A(_08122_),
    .B(_08123_),
    .C(_08225_),
    .Y(_08226_));
 XNOR2x1_ASAP7_75t_R _15294_ (.B(_08226_),
    .Y(_08227_),
    .A(net70));
 AND2x2_ASAP7_75t_R _15295_ (.A(_05777_),
    .B(_08227_),
    .Y(_08228_));
 AND2x2_ASAP7_75t_R _15296_ (.A(_08084_),
    .B(_08228_),
    .Y(_08229_));
 OR5x2_ASAP7_75t_R _15297_ (.A(_01091_),
    .B(_01094_),
    .C(_01097_),
    .D(_01100_),
    .E(_01103_),
    .Y(_08230_));
 OA21x2_ASAP7_75t_R _15298_ (.A1(_01098_),
    .A2(_01097_),
    .B(_01101_),
    .Y(_08231_));
 OR4x1_ASAP7_75t_R _15299_ (.A(_01095_),
    .B(_01094_),
    .C(_01097_),
    .D(_01100_),
    .Y(_08232_));
 OA211x2_ASAP7_75t_R _15300_ (.A1(_01100_),
    .A2(_08231_),
    .B(_08232_),
    .C(_01104_),
    .Y(_08233_));
 OA21x2_ASAP7_75t_R _15301_ (.A1(_01103_),
    .A2(_08233_),
    .B(_01107_),
    .Y(_08234_));
 OA21x2_ASAP7_75t_R _15302_ (.A1(_08136_),
    .A2(_08230_),
    .B(_08234_),
    .Y(_08235_));
 XOR2x1_ASAP7_75t_R _15303_ (.A(_01106_),
    .Y(_08236_),
    .B(_08235_));
 AND4x1_ASAP7_75t_R _15304_ (.A(_08055_),
    .B(_08062_),
    .C(_08068_),
    .D(_08236_),
    .Y(_08237_));
 AND3x1_ASAP7_75t_R _15305_ (.A(_08063_),
    .B(_08140_),
    .C(_08236_),
    .Y(_08238_));
 AO221x1_ASAP7_75t_R _15306_ (.A1(_08082_),
    .A2(_08227_),
    .B1(_08228_),
    .B2(_08087_),
    .C(_08238_),
    .Y(_08239_));
 OR3x4_ASAP7_75t_R _15307_ (.A(_08229_),
    .B(_08237_),
    .C(_08239_),
    .Y(_08240_));
 AO21x1_ASAP7_75t_R _15308_ (.A1(\readdata[14] ),
    .A2(_08179_),
    .B(_08182_),
    .Y(_08241_));
 OAI21x1_ASAP7_75t_R _15309_ (.A1(_08150_),
    .A2(net37),
    .B(_08241_),
    .Y(_08242_));
 BUFx6f_ASAP7_75t_R _15310_ (.A(_08242_),
    .Y(_08243_));
 AOI22x1_ASAP7_75t_R _15311_ (.A1(_00610_),
    .A2(_08144_),
    .B1(_08148_),
    .B2(_08243_),
    .Y(_08244_));
 OA21x2_ASAP7_75t_R _15312_ (.A1(_08121_),
    .A2(_08240_),
    .B(_08244_),
    .Y(_01259_));
 OR3x1_ASAP7_75t_R _15313_ (.A(_01105_),
    .B(_08213_),
    .C(_08225_),
    .Y(_08245_));
 XNOR2x1_ASAP7_75t_R _15314_ (.B(_08245_),
    .Y(_08246_),
    .A(net71));
 AND2x2_ASAP7_75t_R _15315_ (.A(_05777_),
    .B(_08246_),
    .Y(_08247_));
 AND2x2_ASAP7_75t_R _15316_ (.A(_08084_),
    .B(_08247_),
    .Y(_08248_));
 BUFx3_ASAP7_75t_R _15317_ (.A(_08067_),
    .Y(_08249_));
 OA21x2_ASAP7_75t_R _15318_ (.A1(_08171_),
    .A2(_08230_),
    .B(_08234_),
    .Y(_08250_));
 OA21x2_ASAP7_75t_R _15319_ (.A1(_01106_),
    .A2(_08250_),
    .B(_01110_),
    .Y(_08251_));
 XOR2x1_ASAP7_75t_R _15320_ (.A(_01109_),
    .Y(_08252_),
    .B(_08251_));
 AND4x1_ASAP7_75t_R _15321_ (.A(_08055_),
    .B(_08062_),
    .C(_08249_),
    .D(_08252_),
    .Y(_08253_));
 AND3x1_ASAP7_75t_R _15322_ (.A(_08063_),
    .B(_08140_),
    .C(_08252_),
    .Y(_08254_));
 AO221x1_ASAP7_75t_R _15323_ (.A1(_08082_),
    .A2(_08246_),
    .B1(_08247_),
    .B2(_08087_),
    .C(_08254_),
    .Y(_08255_));
 OR3x4_ASAP7_75t_R _15324_ (.A(_08248_),
    .B(_08253_),
    .C(_08255_),
    .Y(_08256_));
 AO21x1_ASAP7_75t_R _15325_ (.A1(\readdata[15] ),
    .A2(_08179_),
    .B(_08182_),
    .Y(_08257_));
 OAI21x1_ASAP7_75t_R _15326_ (.A1(_08150_),
    .A2(net38),
    .B(_08257_),
    .Y(_08258_));
 BUFx6f_ASAP7_75t_R _15327_ (.A(_08258_),
    .Y(_08259_));
 AOI22x1_ASAP7_75t_R _15328_ (.A1(_00576_),
    .A2(_08144_),
    .B1(_08148_),
    .B2(_08259_),
    .Y(_08260_));
 OA21x2_ASAP7_75t_R _15329_ (.A1(_08121_),
    .A2(_08256_),
    .B(_08260_),
    .Y(_01260_));
 OR3x2_ASAP7_75t_R _15330_ (.A(_01105_),
    .B(_01108_),
    .C(_08225_),
    .Y(_08261_));
 NOR2x1_ASAP7_75t_R _15331_ (.A(_08125_),
    .B(_08261_),
    .Y(_08262_));
 XNOR2x1_ASAP7_75t_R _15332_ (.B(_08262_),
    .Y(_08263_),
    .A(_01111_));
 AND2x2_ASAP7_75t_R _15333_ (.A(_05777_),
    .B(_08263_),
    .Y(_08264_));
 AND2x2_ASAP7_75t_R _15334_ (.A(_08084_),
    .B(_08264_),
    .Y(_08265_));
 OR3x1_ASAP7_75t_R _15335_ (.A(_01085_),
    .B(_01088_),
    .C(_08230_),
    .Y(_08266_));
 OR2x2_ASAP7_75t_R _15336_ (.A(_01089_),
    .B(_01088_),
    .Y(_08267_));
 AO21x1_ASAP7_75t_R _15337_ (.A1(_01092_),
    .A2(_08267_),
    .B(_08230_),
    .Y(_08268_));
 AND3x1_ASAP7_75t_R _15338_ (.A(_01110_),
    .B(_01113_),
    .C(_08234_),
    .Y(_08269_));
 OA211x2_ASAP7_75t_R _15339_ (.A1(_08134_),
    .A2(_08266_),
    .B(_08268_),
    .C(_08269_),
    .Y(_08270_));
 AND3x1_ASAP7_75t_R _15340_ (.A(_01106_),
    .B(_01110_),
    .C(_01113_),
    .Y(_08271_));
 AO21x2_ASAP7_75t_R _15341_ (.A1(_01109_),
    .A2(_01113_),
    .B(_08271_),
    .Y(_08272_));
 NOR2x1_ASAP7_75t_R _15342_ (.A(_08270_),
    .B(_08272_),
    .Y(_08273_));
 XNOR2x1_ASAP7_75t_R _15343_ (.B(_08273_),
    .Y(_08274_),
    .A(_01112_));
 AND4x1_ASAP7_75t_R _15344_ (.A(_08055_),
    .B(_08062_),
    .C(_08249_),
    .D(_08274_),
    .Y(_08275_));
 BUFx3_ASAP7_75t_R _15345_ (.A(_08066_),
    .Y(_08276_));
 AND3x1_ASAP7_75t_R _15346_ (.A(_08063_),
    .B(_08276_),
    .C(_08274_),
    .Y(_08277_));
 AO221x1_ASAP7_75t_R _15347_ (.A1(_08082_),
    .A2(_08263_),
    .B1(_08264_),
    .B2(_08087_),
    .C(_08277_),
    .Y(_08278_));
 OR3x4_ASAP7_75t_R _15348_ (.A(_08265_),
    .B(_08275_),
    .C(_08278_),
    .Y(_08279_));
 OR4x2_ASAP7_75t_R _15349_ (.A(_03713_),
    .B(_03212_),
    .C(_06929_),
    .D(_06935_),
    .Y(_08280_));
 BUFx3_ASAP7_75t_R _15350_ (.A(_08280_),
    .Y(_08281_));
 AND4x2_ASAP7_75t_R _15351_ (.A(\readdata[15] ),
    .B(_08149_),
    .C(_06826_),
    .D(_06928_),
    .Y(_08282_));
 BUFx3_ASAP7_75t_R _15352_ (.A(_08282_),
    .Y(_08283_));
 AO21x1_ASAP7_75t_R _15353_ (.A1(\readdata[16] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08284_));
 AO21x1_ASAP7_75t_R _15354_ (.A1(_08188_),
    .A2(_08284_),
    .B(_08182_),
    .Y(_08285_));
 OAI21x1_ASAP7_75t_R _15355_ (.A1(_08150_),
    .A2(net39),
    .B(_08285_),
    .Y(_08286_));
 BUFx6f_ASAP7_75t_R _15356_ (.A(_08286_),
    .Y(_08287_));
 AOI22x1_ASAP7_75t_R _15357_ (.A1(_00543_),
    .A2(_08144_),
    .B1(_08148_),
    .B2(_08287_),
    .Y(_08288_));
 OA21x2_ASAP7_75t_R _15358_ (.A1(_08121_),
    .A2(_08279_),
    .B(_08288_),
    .Y(_01261_));
 BUFx3_ASAP7_75t_R _15359_ (.A(_08077_),
    .Y(_08289_));
 OR3x1_ASAP7_75t_R _15360_ (.A(_01111_),
    .B(_08213_),
    .C(_08261_),
    .Y(_08290_));
 XNOR2x1_ASAP7_75t_R _15361_ (.B(_08290_),
    .Y(_08291_),
    .A(net73));
 AND2x2_ASAP7_75t_R _15362_ (.A(_05777_),
    .B(_08291_),
    .Y(_08292_));
 AND2x2_ASAP7_75t_R _15363_ (.A(_08289_),
    .B(_08292_),
    .Y(_08293_));
 OA211x2_ASAP7_75t_R _15364_ (.A1(_08169_),
    .A2(_08266_),
    .B(_08268_),
    .C(_08269_),
    .Y(_08294_));
 OR3x1_ASAP7_75t_R _15365_ (.A(_01112_),
    .B(_08272_),
    .C(_08294_),
    .Y(_08295_));
 NAND2x1_ASAP7_75t_R _15366_ (.A(_01116_),
    .B(_08295_),
    .Y(_08296_));
 XNOR2x1_ASAP7_75t_R _15367_ (.B(_08296_),
    .Y(_08297_),
    .A(_01115_));
 AND4x1_ASAP7_75t_R _15368_ (.A(_08055_),
    .B(_08062_),
    .C(_08249_),
    .D(_08297_),
    .Y(_08298_));
 AND3x1_ASAP7_75t_R _15369_ (.A(_08063_),
    .B(_08276_),
    .C(_08297_),
    .Y(_08299_));
 AO221x1_ASAP7_75t_R _15370_ (.A1(_08082_),
    .A2(_08291_),
    .B1(_08292_),
    .B2(_08087_),
    .C(_08299_),
    .Y(_08300_));
 OR3x4_ASAP7_75t_R _15371_ (.A(_08293_),
    .B(_08298_),
    .C(_08300_),
    .Y(_08301_));
 BUFx12_ASAP7_75t_R _15372_ (.A(_08118_),
    .Y(_08302_));
 AO21x1_ASAP7_75t_R _15373_ (.A1(\readdata[17] ),
    .A2(_08280_),
    .B(_08282_),
    .Y(_08303_));
 BUFx4f_ASAP7_75t_R _15374_ (.A(_08181_),
    .Y(_08304_));
 AOI21x1_ASAP7_75t_R _15375_ (.A1(_08179_),
    .A2(_08303_),
    .B(_08304_),
    .Y(_08305_));
 AO21x1_ASAP7_75t_R _15376_ (.A1(_08108_),
    .A2(_07579_),
    .B(_08305_),
    .Y(_08306_));
 BUFx6f_ASAP7_75t_R _15377_ (.A(_08306_),
    .Y(_08307_));
 BUFx6f_ASAP7_75t_R _15378_ (.A(_08307_),
    .Y(_08308_));
 AOI22x1_ASAP7_75t_R _15379_ (.A1(_00510_),
    .A2(_08302_),
    .B1(_08148_),
    .B2(_08308_),
    .Y(_08309_));
 OA21x2_ASAP7_75t_R _15380_ (.A1(_08121_),
    .A2(_08301_),
    .B(_08309_),
    .Y(_01262_));
 OR4x1_ASAP7_75t_R _15381_ (.A(_01111_),
    .B(_01114_),
    .C(_08125_),
    .D(_08261_),
    .Y(_08310_));
 XNOR2x1_ASAP7_75t_R _15382_ (.B(_08310_),
    .Y(_08311_),
    .A(net74));
 AND2x2_ASAP7_75t_R _15383_ (.A(_05777_),
    .B(_08311_),
    .Y(_08312_));
 AND2x2_ASAP7_75t_R _15384_ (.A(_08289_),
    .B(_08312_),
    .Y(_08313_));
 OR2x2_ASAP7_75t_R _15385_ (.A(_01112_),
    .B(_01115_),
    .Y(_08314_));
 OR2x2_ASAP7_75t_R _15386_ (.A(_01116_),
    .B(_01115_),
    .Y(_08315_));
 AND2x2_ASAP7_75t_R _15387_ (.A(_01119_),
    .B(_08315_),
    .Y(_08316_));
 OA31x2_ASAP7_75t_R _15388_ (.A1(_08270_),
    .A2(_08272_),
    .A3(_08314_),
    .B1(_08316_),
    .Y(_08317_));
 XOR2x2_ASAP7_75t_R _15389_ (.A(_01118_),
    .B(_08317_),
    .Y(_08318_));
 AND4x1_ASAP7_75t_R _15390_ (.A(_08055_),
    .B(_08062_),
    .C(_08249_),
    .D(_08318_),
    .Y(_08319_));
 BUFx3_ASAP7_75t_R _15391_ (.A(_08081_),
    .Y(_08320_));
 AND3x1_ASAP7_75t_R _15392_ (.A(_08063_),
    .B(_08276_),
    .C(_08318_),
    .Y(_08321_));
 AO221x1_ASAP7_75t_R _15393_ (.A1(_08320_),
    .A2(_08311_),
    .B1(_08312_),
    .B2(_08087_),
    .C(_08321_),
    .Y(_08322_));
 OR3x4_ASAP7_75t_R _15394_ (.A(_08313_),
    .B(_08319_),
    .C(_08322_),
    .Y(_08323_));
 AO21x1_ASAP7_75t_R _15395_ (.A1(\readdata[18] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08324_));
 AO21x1_ASAP7_75t_R _15396_ (.A1(_08188_),
    .A2(_08324_),
    .B(_08182_),
    .Y(_08325_));
 OAI21x1_ASAP7_75t_R _15397_ (.A1(_08150_),
    .A2(net41),
    .B(_08325_),
    .Y(_08326_));
 BUFx6f_ASAP7_75t_R _15398_ (.A(_08326_),
    .Y(_08327_));
 AOI22x1_ASAP7_75t_R _15399_ (.A1(_00477_),
    .A2(_08302_),
    .B1(_08148_),
    .B2(_08327_),
    .Y(_08328_));
 OA21x2_ASAP7_75t_R _15400_ (.A1(_08121_),
    .A2(_08323_),
    .B(_08328_),
    .Y(_01263_));
 BUFx3_ASAP7_75t_R _15401_ (.A(_05775_),
    .Y(_08329_));
 OR4x2_ASAP7_75t_R _15402_ (.A(_01111_),
    .B(_01114_),
    .C(_01117_),
    .D(_08261_),
    .Y(_08330_));
 NOR2x1_ASAP7_75t_R _15403_ (.A(_08213_),
    .B(_08330_),
    .Y(_08331_));
 XNOR2x1_ASAP7_75t_R _15404_ (.B(_08331_),
    .Y(_08332_),
    .A(_01120_));
 AND2x2_ASAP7_75t_R _15405_ (.A(_08329_),
    .B(_08332_),
    .Y(_08333_));
 AND2x2_ASAP7_75t_R _15406_ (.A(_08289_),
    .B(_08333_),
    .Y(_08334_));
 BUFx4f_ASAP7_75t_R _15407_ (.A(_08054_),
    .Y(_08335_));
 OR4x1_ASAP7_75t_R _15408_ (.A(_01118_),
    .B(_08272_),
    .C(_08294_),
    .D(_08314_),
    .Y(_08336_));
 AO21x1_ASAP7_75t_R _15409_ (.A1(_01119_),
    .A2(_08315_),
    .B(_01118_),
    .Y(_08337_));
 AND3x1_ASAP7_75t_R _15410_ (.A(_01122_),
    .B(_08336_),
    .C(_08337_),
    .Y(_08338_));
 XOR2x1_ASAP7_75t_R _15411_ (.A(_01121_),
    .Y(_08339_),
    .B(_08338_));
 AND4x1_ASAP7_75t_R _15412_ (.A(_08335_),
    .B(_08062_),
    .C(_08249_),
    .D(_08339_),
    .Y(_08340_));
 BUFx4f_ASAP7_75t_R _15413_ (.A(_03256_),
    .Y(_08341_));
 AND3x1_ASAP7_75t_R _15414_ (.A(_08341_),
    .B(_08276_),
    .C(_08339_),
    .Y(_08342_));
 AO221x1_ASAP7_75t_R _15415_ (.A1(_08320_),
    .A2(_08332_),
    .B1(_08333_),
    .B2(_08087_),
    .C(_08342_),
    .Y(_08343_));
 OR3x4_ASAP7_75t_R _15416_ (.A(_08334_),
    .B(_08340_),
    .C(_08343_),
    .Y(_08344_));
 AO21x1_ASAP7_75t_R _15417_ (.A1(\readdata[19] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08345_));
 AO21x1_ASAP7_75t_R _15418_ (.A1(_08188_),
    .A2(_08345_),
    .B(_08182_),
    .Y(_08346_));
 OAI21x1_ASAP7_75t_R _15419_ (.A1(_08150_),
    .A2(net42),
    .B(_08346_),
    .Y(_08347_));
 BUFx6f_ASAP7_75t_R _15420_ (.A(_08347_),
    .Y(_08348_));
 AOI22x1_ASAP7_75t_R _15421_ (.A1(_00444_),
    .A2(_08302_),
    .B1(_08148_),
    .B2(_08348_),
    .Y(_08349_));
 OA21x2_ASAP7_75t_R _15422_ (.A1(_08121_),
    .A2(_08344_),
    .B(_08349_),
    .Y(_01264_));
 AND4x1_ASAP7_75t_R _15423_ (.A(_06826_),
    .B(_06930_),
    .C(_08022_),
    .D(_08057_),
    .Y(_08350_));
 OR3x1_ASAP7_75t_R _15424_ (.A(_03713_),
    .B(_06927_),
    .C(_06929_),
    .Y(_08351_));
 AOI21x1_ASAP7_75t_R _15425_ (.A1(_08022_),
    .A2(_08057_),
    .B(_08351_),
    .Y(_08352_));
 OR4x1_ASAP7_75t_R _15426_ (.A(_08075_),
    .B(_08350_),
    .C(_08352_),
    .D(_08081_),
    .Y(_08353_));
 OR3x1_ASAP7_75t_R _15427_ (.A(net76),
    .B(_03249_),
    .C(_03254_),
    .Y(_08354_));
 AO31x2_ASAP7_75t_R _15428_ (.A1(_08021_),
    .A2(_08048_),
    .A3(_08053_),
    .B(_08354_),
    .Y(_08355_));
 NAND2x1_ASAP7_75t_R _15429_ (.A(_01070_),
    .B(_03256_),
    .Y(_08356_));
 AO211x2_ASAP7_75t_R _15430_ (.A1(_08043_),
    .A2(_08065_),
    .B(_08356_),
    .C(_05467_),
    .Y(_08357_));
 OA21x2_ASAP7_75t_R _15431_ (.A1(net76),
    .A2(_08088_),
    .B(_08357_),
    .Y(_08358_));
 OA31x2_ASAP7_75t_R _15432_ (.A1(_08058_),
    .A2(_08060_),
    .A3(_08354_),
    .B1(_08358_),
    .Y(_08359_));
 OA211x2_ASAP7_75t_R _15433_ (.A1(_08084_),
    .A2(_08353_),
    .B(_08355_),
    .C(_08359_),
    .Y(_08360_));
 BUFx6f_ASAP7_75t_R _15434_ (.A(_08149_),
    .Y(_08361_));
 OA21x2_ASAP7_75t_R _15435_ (.A1(\readdata[1] ),
    .A2(_06935_),
    .B(_08113_),
    .Y(_08362_));
 OA21x2_ASAP7_75t_R _15436_ (.A1(_08361_),
    .A2(net43),
    .B(_08362_),
    .Y(_08363_));
 AO21x2_ASAP7_75t_R _15437_ (.A1(_08106_),
    .A2(_08360_),
    .B(_08363_),
    .Y(_08364_));
 NAND2x1_ASAP7_75t_R _15438_ (.A(_01042_),
    .B(_08144_),
    .Y(_08365_));
 OA21x2_ASAP7_75t_R _15439_ (.A1(_08144_),
    .A2(_08364_),
    .B(_08365_),
    .Y(_01265_));
 OR3x1_ASAP7_75t_R _15440_ (.A(_01120_),
    .B(_08125_),
    .C(_08330_),
    .Y(_08366_));
 XNOR2x1_ASAP7_75t_R _15441_ (.B(_08366_),
    .Y(_08367_),
    .A(net77));
 AND2x2_ASAP7_75t_R _15442_ (.A(_08329_),
    .B(_08367_),
    .Y(_08368_));
 AND2x2_ASAP7_75t_R _15443_ (.A(_08289_),
    .B(_08368_),
    .Y(_08369_));
 BUFx4f_ASAP7_75t_R _15444_ (.A(_08061_),
    .Y(_08370_));
 OA21x2_ASAP7_75t_R _15445_ (.A1(_01118_),
    .A2(_08317_),
    .B(_01122_),
    .Y(_08371_));
 OA21x2_ASAP7_75t_R _15446_ (.A1(_01121_),
    .A2(_08371_),
    .B(_01125_),
    .Y(_08372_));
 XOR2x1_ASAP7_75t_R _15447_ (.A(_01124_),
    .Y(_08373_),
    .B(_08372_));
 AND4x1_ASAP7_75t_R _15448_ (.A(_08335_),
    .B(_08370_),
    .C(_08249_),
    .D(_08373_),
    .Y(_08374_));
 BUFx3_ASAP7_75t_R _15449_ (.A(_08079_),
    .Y(_08375_));
 AND3x1_ASAP7_75t_R _15450_ (.A(_08341_),
    .B(_08276_),
    .C(_08373_),
    .Y(_08376_));
 AO221x1_ASAP7_75t_R _15451_ (.A1(_08320_),
    .A2(_08367_),
    .B1(_08368_),
    .B2(_08375_),
    .C(_08376_),
    .Y(_08377_));
 OR3x4_ASAP7_75t_R _15452_ (.A(_08369_),
    .B(_08374_),
    .C(_08377_),
    .Y(_08378_));
 AO21x1_ASAP7_75t_R _15453_ (.A1(\readdata[20] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08379_));
 AO21x1_ASAP7_75t_R _15454_ (.A1(_08188_),
    .A2(_08379_),
    .B(_08182_),
    .Y(_08380_));
 OAI21x1_ASAP7_75t_R _15455_ (.A1(_08361_),
    .A2(net44),
    .B(_08380_),
    .Y(_08381_));
 BUFx6f_ASAP7_75t_R _15456_ (.A(_08381_),
    .Y(_08382_));
 AOI22x1_ASAP7_75t_R _15457_ (.A1(_00411_),
    .A2(_08302_),
    .B1(_08148_),
    .B2(_08382_),
    .Y(_08383_));
 OA21x2_ASAP7_75t_R _15458_ (.A1(_08121_),
    .A2(_08378_),
    .B(_08383_),
    .Y(_01266_));
 OR4x1_ASAP7_75t_R _15459_ (.A(_01120_),
    .B(_01123_),
    .C(_08213_),
    .D(_08330_),
    .Y(_08384_));
 XNOR2x2_ASAP7_75t_R _15460_ (.A(net78),
    .B(_08384_),
    .Y(_08385_));
 AND2x2_ASAP7_75t_R _15461_ (.A(_05776_),
    .B(_08385_),
    .Y(_08386_));
 AND2x2_ASAP7_75t_R _15462_ (.A(_08077_),
    .B(_08386_),
    .Y(_08387_));
 AND3x1_ASAP7_75t_R _15463_ (.A(_01122_),
    .B(_01125_),
    .C(_01128_),
    .Y(_08388_));
 AND3x1_ASAP7_75t_R _15464_ (.A(_01121_),
    .B(_01125_),
    .C(_01128_),
    .Y(_08389_));
 AO21x1_ASAP7_75t_R _15465_ (.A1(_01124_),
    .A2(_01128_),
    .B(_08389_),
    .Y(_08390_));
 AO31x2_ASAP7_75t_R _15466_ (.A1(_08336_),
    .A2(_08337_),
    .A3(_08388_),
    .B(_08390_),
    .Y(_08391_));
 XOR2x2_ASAP7_75t_R _15467_ (.A(_01127_),
    .B(_08391_),
    .Y(_08392_));
 AND4x1_ASAP7_75t_R _15468_ (.A(_08196_),
    .B(_08197_),
    .C(_08140_),
    .D(_08392_),
    .Y(_08393_));
 AND3x1_ASAP7_75t_R _15469_ (.A(_08203_),
    .B(_08088_),
    .C(_08392_),
    .Y(_08394_));
 AO221x1_ASAP7_75t_R _15470_ (.A1(_08202_),
    .A2(_08385_),
    .B1(_08386_),
    .B2(_08080_),
    .C(_08394_),
    .Y(_08395_));
 OR3x4_ASAP7_75t_R _15471_ (.A(_08387_),
    .B(_08393_),
    .C(_08395_),
    .Y(_08396_));
 AO21x1_ASAP7_75t_R _15472_ (.A1(\readdata[21] ),
    .A2(_08280_),
    .B(_08282_),
    .Y(_08397_));
 AO21x1_ASAP7_75t_R _15473_ (.A1(_08151_),
    .A2(_08397_),
    .B(_08152_),
    .Y(_08398_));
 AND2x2_ASAP7_75t_R _15474_ (.A(_08149_),
    .B(_08398_),
    .Y(_08399_));
 AO211x2_ASAP7_75t_R _15475_ (.A1(_08108_),
    .A2(net45),
    .B(_08106_),
    .C(_08399_),
    .Y(_08400_));
 BUFx6f_ASAP7_75t_R _15476_ (.A(_08400_),
    .Y(_08401_));
 BUFx6f_ASAP7_75t_R _15477_ (.A(_08118_),
    .Y(_08402_));
 NAND2x1_ASAP7_75t_R _15478_ (.A(_00378_),
    .B(_08402_),
    .Y(_08403_));
 OA221x2_ASAP7_75t_R _15479_ (.A1(_08107_),
    .A2(_08396_),
    .B1(_08401_),
    .B2(_08144_),
    .C(_08403_),
    .Y(_01267_));
 OR5x2_ASAP7_75t_R _15480_ (.A(_01120_),
    .B(_01123_),
    .C(_01126_),
    .D(_08125_),
    .E(_08330_),
    .Y(_08404_));
 XNOR2x1_ASAP7_75t_R _15481_ (.B(_08404_),
    .Y(_08405_),
    .A(net79));
 AND2x2_ASAP7_75t_R _15482_ (.A(_08329_),
    .B(_08405_),
    .Y(_08406_));
 AND2x2_ASAP7_75t_R _15483_ (.A(_08289_),
    .B(_08406_),
    .Y(_08407_));
 OA21x2_ASAP7_75t_R _15484_ (.A1(_01118_),
    .A2(_08317_),
    .B(_08388_),
    .Y(_08408_));
 OR3x1_ASAP7_75t_R _15485_ (.A(_01127_),
    .B(_08390_),
    .C(_08408_),
    .Y(_08409_));
 NAND2x1_ASAP7_75t_R _15486_ (.A(_01131_),
    .B(_08409_),
    .Y(_08410_));
 XNOR2x1_ASAP7_75t_R _15487_ (.B(_08410_),
    .Y(_08411_),
    .A(_01130_));
 AND4x1_ASAP7_75t_R _15488_ (.A(_08335_),
    .B(_08370_),
    .C(_08249_),
    .D(_08411_),
    .Y(_08412_));
 AND3x1_ASAP7_75t_R _15489_ (.A(_08341_),
    .B(_08276_),
    .C(_08411_),
    .Y(_08413_));
 AO221x1_ASAP7_75t_R _15490_ (.A1(_08320_),
    .A2(_08405_),
    .B1(_08406_),
    .B2(_08375_),
    .C(_08413_),
    .Y(_08414_));
 OR3x4_ASAP7_75t_R _15491_ (.A(_08407_),
    .B(_08412_),
    .C(_08414_),
    .Y(_08415_));
 BUFx6f_ASAP7_75t_R _15492_ (.A(_08147_),
    .Y(_08416_));
 AO21x1_ASAP7_75t_R _15493_ (.A1(\readdata[22] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08417_));
 AO21x1_ASAP7_75t_R _15494_ (.A1(_08188_),
    .A2(_08417_),
    .B(_08304_),
    .Y(_08418_));
 OAI21x1_ASAP7_75t_R _15495_ (.A1(_08361_),
    .A2(net46),
    .B(_08418_),
    .Y(_08419_));
 BUFx6f_ASAP7_75t_R _15496_ (.A(_08419_),
    .Y(_08420_));
 AOI22x1_ASAP7_75t_R _15497_ (.A1(_00345_),
    .A2(_08302_),
    .B1(_08416_),
    .B2(_08420_),
    .Y(_08421_));
 OA21x2_ASAP7_75t_R _15498_ (.A1(_08121_),
    .A2(_08415_),
    .B(_08421_),
    .Y(_01268_));
 BUFx4f_ASAP7_75t_R _15499_ (.A(_08107_),
    .Y(_08422_));
 OR5x2_ASAP7_75t_R _15500_ (.A(_01120_),
    .B(_01123_),
    .C(_01126_),
    .D(_01129_),
    .E(_08330_),
    .Y(_08423_));
 NOR2x1_ASAP7_75t_R _15501_ (.A(_08213_),
    .B(_08423_),
    .Y(_08424_));
 XNOR2x1_ASAP7_75t_R _15502_ (.B(_08424_),
    .Y(_08425_),
    .A(_01132_));
 AND2x2_ASAP7_75t_R _15503_ (.A(_08329_),
    .B(_08425_),
    .Y(_08426_));
 AND2x2_ASAP7_75t_R _15504_ (.A(_08289_),
    .B(_08426_),
    .Y(_08427_));
 OA21x2_ASAP7_75t_R _15505_ (.A1(_01127_),
    .A2(_08391_),
    .B(_01131_),
    .Y(_08428_));
 OA21x2_ASAP7_75t_R _15506_ (.A1(_01130_),
    .A2(_08428_),
    .B(_01134_),
    .Y(_08429_));
 XOR2x1_ASAP7_75t_R _15507_ (.A(_01133_),
    .Y(_08430_),
    .B(_08429_));
 AND4x1_ASAP7_75t_R _15508_ (.A(_08335_),
    .B(_08370_),
    .C(_08249_),
    .D(_08430_),
    .Y(_08431_));
 AND3x1_ASAP7_75t_R _15509_ (.A(_08341_),
    .B(_08276_),
    .C(_08430_),
    .Y(_08432_));
 AO221x1_ASAP7_75t_R _15510_ (.A1(_08320_),
    .A2(_08425_),
    .B1(_08426_),
    .B2(_08375_),
    .C(_08432_),
    .Y(_08433_));
 OR3x4_ASAP7_75t_R _15511_ (.A(_08427_),
    .B(_08431_),
    .C(_08433_),
    .Y(_08434_));
 AO21x1_ASAP7_75t_R _15512_ (.A1(\readdata[23] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08435_));
 AO21x1_ASAP7_75t_R _15513_ (.A1(_08188_),
    .A2(_08435_),
    .B(_08304_),
    .Y(_08436_));
 OAI21x1_ASAP7_75t_R _15514_ (.A1(_08361_),
    .A2(net47),
    .B(_08436_),
    .Y(_08437_));
 BUFx6f_ASAP7_75t_R _15515_ (.A(_08437_),
    .Y(_08438_));
 AOI22x1_ASAP7_75t_R _15516_ (.A1(_00311_),
    .A2(_08302_),
    .B1(_08416_),
    .B2(_08438_),
    .Y(_08439_));
 OA21x2_ASAP7_75t_R _15517_ (.A1(_08422_),
    .A2(_08434_),
    .B(_08439_),
    .Y(_01269_));
 OR2x2_ASAP7_75t_R _15518_ (.A(_01132_),
    .B(_08423_),
    .Y(_08440_));
 NOR2x1_ASAP7_75t_R _15519_ (.A(_08125_),
    .B(_08440_),
    .Y(_08441_));
 XNOR2x1_ASAP7_75t_R _15520_ (.B(_08441_),
    .Y(_08442_),
    .A(_01135_));
 AND2x2_ASAP7_75t_R _15521_ (.A(_08329_),
    .B(_08442_),
    .Y(_08443_));
 AND2x2_ASAP7_75t_R _15522_ (.A(_08289_),
    .B(_08443_),
    .Y(_08444_));
 OR3x1_ASAP7_75t_R _15523_ (.A(_01127_),
    .B(_01130_),
    .C(_01133_),
    .Y(_08445_));
 OR3x1_ASAP7_75t_R _15524_ (.A(_08390_),
    .B(_08408_),
    .C(_08445_),
    .Y(_08446_));
 OR2x2_ASAP7_75t_R _15525_ (.A(_01131_),
    .B(_01130_),
    .Y(_08447_));
 AO21x1_ASAP7_75t_R _15526_ (.A1(_01134_),
    .A2(_08447_),
    .B(_01133_),
    .Y(_08448_));
 AND2x2_ASAP7_75t_R _15527_ (.A(_08446_),
    .B(_08448_),
    .Y(_08449_));
 NAND2x1_ASAP7_75t_R _15528_ (.A(_01137_),
    .B(_08449_),
    .Y(_08450_));
 XNOR2x1_ASAP7_75t_R _15529_ (.B(_08450_),
    .Y(_08451_),
    .A(_01136_));
 AND4x1_ASAP7_75t_R _15530_ (.A(_08335_),
    .B(_08370_),
    .C(_08249_),
    .D(_08451_),
    .Y(_08452_));
 AND3x1_ASAP7_75t_R _15531_ (.A(_08341_),
    .B(_08276_),
    .C(_08451_),
    .Y(_08453_));
 AO221x1_ASAP7_75t_R _15532_ (.A1(_08320_),
    .A2(_08442_),
    .B1(_08443_),
    .B2(_08375_),
    .C(_08453_),
    .Y(_08454_));
 OR3x4_ASAP7_75t_R _15533_ (.A(_08444_),
    .B(_08452_),
    .C(_08454_),
    .Y(_08455_));
 AO21x1_ASAP7_75t_R _15534_ (.A1(\readdata[24] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08456_));
 AO21x1_ASAP7_75t_R _15535_ (.A1(_08188_),
    .A2(_08456_),
    .B(_08304_),
    .Y(_08457_));
 OAI21x1_ASAP7_75t_R _15536_ (.A1(_08361_),
    .A2(net48),
    .B(_08457_),
    .Y(_08458_));
 BUFx6f_ASAP7_75t_R _15537_ (.A(_08458_),
    .Y(_08459_));
 AOI22x1_ASAP7_75t_R _15538_ (.A1(_00278_),
    .A2(_08302_),
    .B1(_08416_),
    .B2(_08459_),
    .Y(_08460_));
 OA21x2_ASAP7_75t_R _15539_ (.A1(_08422_),
    .A2(_08455_),
    .B(_08460_),
    .Y(_01270_));
 OR3x1_ASAP7_75t_R _15540_ (.A(_01135_),
    .B(_08213_),
    .C(_08440_),
    .Y(_08461_));
 XNOR2x1_ASAP7_75t_R _15541_ (.B(_08461_),
    .Y(_08462_),
    .A(net82));
 AND2x2_ASAP7_75t_R _15542_ (.A(_08329_),
    .B(_08462_),
    .Y(_08463_));
 AND2x2_ASAP7_75t_R _15543_ (.A(_08289_),
    .B(_08463_),
    .Y(_08464_));
 OA21x2_ASAP7_75t_R _15544_ (.A1(_08391_),
    .A2(_08445_),
    .B(_08448_),
    .Y(_08465_));
 AO21x1_ASAP7_75t_R _15545_ (.A1(_01137_),
    .A2(_08465_),
    .B(_01136_),
    .Y(_08466_));
 AND2x2_ASAP7_75t_R _15546_ (.A(_01140_),
    .B(_08466_),
    .Y(_08467_));
 XOR2x1_ASAP7_75t_R _15547_ (.A(_01139_),
    .Y(_08468_),
    .B(_08467_));
 AND4x1_ASAP7_75t_R _15548_ (.A(_08335_),
    .B(_08370_),
    .C(_08249_),
    .D(_08468_),
    .Y(_08469_));
 AND3x1_ASAP7_75t_R _15549_ (.A(_08341_),
    .B(_08276_),
    .C(_08468_),
    .Y(_08470_));
 AO221x1_ASAP7_75t_R _15550_ (.A1(_08320_),
    .A2(_08462_),
    .B1(_08463_),
    .B2(_08375_),
    .C(_08470_),
    .Y(_08471_));
 OR3x4_ASAP7_75t_R _15551_ (.A(_08464_),
    .B(_08469_),
    .C(_08471_),
    .Y(_08472_));
 AO21x1_ASAP7_75t_R _15552_ (.A1(\readdata[25] ),
    .A2(_08280_),
    .B(_08282_),
    .Y(_08473_));
 AOI21x1_ASAP7_75t_R _15553_ (.A1(_08179_),
    .A2(_08473_),
    .B(_08304_),
    .Y(_08474_));
 AO21x1_ASAP7_75t_R _15554_ (.A1(_08108_),
    .A2(_07743_),
    .B(_08474_),
    .Y(_08475_));
 BUFx12f_ASAP7_75t_R _15555_ (.A(_08475_),
    .Y(_08476_));
 BUFx6f_ASAP7_75t_R _15556_ (.A(_08476_),
    .Y(_08477_));
 AOI22x1_ASAP7_75t_R _15557_ (.A1(_00245_),
    .A2(_08302_),
    .B1(_08416_),
    .B2(_08477_),
    .Y(_08478_));
 OA21x2_ASAP7_75t_R _15558_ (.A1(_08422_),
    .A2(_08472_),
    .B(_08478_),
    .Y(_01271_));
 OR4x1_ASAP7_75t_R _15559_ (.A(_01135_),
    .B(_01138_),
    .C(_08125_),
    .D(_08440_),
    .Y(_08479_));
 XNOR2x1_ASAP7_75t_R _15560_ (.B(_08479_),
    .Y(_08480_),
    .A(net83));
 AND2x2_ASAP7_75t_R _15561_ (.A(_08329_),
    .B(_08480_),
    .Y(_08481_));
 AND2x2_ASAP7_75t_R _15562_ (.A(_08289_),
    .B(_08481_),
    .Y(_08482_));
 AND3x1_ASAP7_75t_R _15563_ (.A(_01137_),
    .B(_01140_),
    .C(_01143_),
    .Y(_08483_));
 AND3x1_ASAP7_75t_R _15564_ (.A(_01136_),
    .B(_01140_),
    .C(_01143_),
    .Y(_08484_));
 AO21x1_ASAP7_75t_R _15565_ (.A1(_01139_),
    .A2(_01143_),
    .B(_08484_),
    .Y(_08485_));
 AO21x1_ASAP7_75t_R _15566_ (.A1(_08449_),
    .A2(_08483_),
    .B(_08485_),
    .Y(_08486_));
 XOR2x1_ASAP7_75t_R _15567_ (.A(_01142_),
    .Y(_08487_),
    .B(_08486_));
 AND4x1_ASAP7_75t_R _15568_ (.A(_08335_),
    .B(_08370_),
    .C(_08089_),
    .D(_08487_),
    .Y(_08488_));
 AND3x1_ASAP7_75t_R _15569_ (.A(_08341_),
    .B(_08276_),
    .C(_08487_),
    .Y(_08489_));
 AO221x1_ASAP7_75t_R _15570_ (.A1(_08320_),
    .A2(_08480_),
    .B1(_08481_),
    .B2(_08375_),
    .C(_08489_),
    .Y(_08490_));
 OR3x4_ASAP7_75t_R _15571_ (.A(_08482_),
    .B(_08488_),
    .C(_08490_),
    .Y(_08491_));
 AO21x1_ASAP7_75t_R _15572_ (.A1(\readdata[26] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08492_));
 AO21x1_ASAP7_75t_R _15573_ (.A1(_08179_),
    .A2(_08492_),
    .B(_08304_),
    .Y(_08493_));
 OAI21x1_ASAP7_75t_R _15574_ (.A1(_08361_),
    .A2(net50),
    .B(_08493_),
    .Y(_08494_));
 BUFx6f_ASAP7_75t_R _15575_ (.A(_08494_),
    .Y(_08495_));
 AOI22x1_ASAP7_75t_R _15576_ (.A1(_00211_),
    .A2(_08302_),
    .B1(_08416_),
    .B2(_08495_),
    .Y(_08496_));
 OA21x2_ASAP7_75t_R _15577_ (.A1(_08422_),
    .A2(_08491_),
    .B(_08496_),
    .Y(_01272_));
 OR4x1_ASAP7_75t_R _15578_ (.A(_01135_),
    .B(_01138_),
    .C(_01141_),
    .D(_08440_),
    .Y(_08497_));
 NOR2x1_ASAP7_75t_R _15579_ (.A(_08213_),
    .B(_08497_),
    .Y(_08498_));
 XNOR2x1_ASAP7_75t_R _15580_ (.B(_08498_),
    .Y(_08499_),
    .A(_01144_));
 AND2x2_ASAP7_75t_R _15581_ (.A(_08329_),
    .B(_08499_),
    .Y(_08500_));
 AND2x2_ASAP7_75t_R _15582_ (.A(_08289_),
    .B(_08500_),
    .Y(_08501_));
 AO21x1_ASAP7_75t_R _15583_ (.A1(_08465_),
    .A2(_08483_),
    .B(_08485_),
    .Y(_08502_));
 OA21x2_ASAP7_75t_R _15584_ (.A1(_01142_),
    .A2(_08502_),
    .B(_01146_),
    .Y(_08503_));
 XOR2x1_ASAP7_75t_R _15585_ (.A(_01145_),
    .Y(_08504_),
    .B(_08503_));
 AND4x1_ASAP7_75t_R _15586_ (.A(_08335_),
    .B(_08370_),
    .C(_08089_),
    .D(_08504_),
    .Y(_08505_));
 AND3x1_ASAP7_75t_R _15587_ (.A(_08341_),
    .B(_08067_),
    .C(_08504_),
    .Y(_08506_));
 AO221x1_ASAP7_75t_R _15588_ (.A1(_08320_),
    .A2(_08499_),
    .B1(_08500_),
    .B2(_08375_),
    .C(_08506_),
    .Y(_08507_));
 OR3x4_ASAP7_75t_R _15589_ (.A(_08501_),
    .B(_08505_),
    .C(_08507_),
    .Y(_08508_));
 AO21x1_ASAP7_75t_R _15590_ (.A1(\readdata[27] ),
    .A2(_08280_),
    .B(_08282_),
    .Y(_08509_));
 AO21x1_ASAP7_75t_R _15591_ (.A1(_08179_),
    .A2(_08509_),
    .B(_08304_),
    .Y(_08510_));
 OAI21x1_ASAP7_75t_R _15592_ (.A1(_08361_),
    .A2(net51),
    .B(_08510_),
    .Y(_08511_));
 BUFx6f_ASAP7_75t_R _15593_ (.A(_08511_),
    .Y(_08512_));
 AOI22x1_ASAP7_75t_R _15594_ (.A1(_00178_),
    .A2(_08302_),
    .B1(_08416_),
    .B2(_08512_),
    .Y(_08513_));
 OA21x2_ASAP7_75t_R _15595_ (.A1(_08422_),
    .A2(_08508_),
    .B(_08513_),
    .Y(_01273_));
 INVx1_ASAP7_75t_R _15596_ (.A(_00144_),
    .Y(_08514_));
 AO21x1_ASAP7_75t_R _15597_ (.A1(\readdata[28] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08515_));
 AO21x1_ASAP7_75t_R _15598_ (.A1(_08188_),
    .A2(_08515_),
    .B(_08182_),
    .Y(_08516_));
 OA21x2_ASAP7_75t_R _15599_ (.A1(_08150_),
    .A2(net52),
    .B(_08516_),
    .Y(_08517_));
 BUFx4f_ASAP7_75t_R _15600_ (.A(_08517_),
    .Y(_08518_));
 OR2x2_ASAP7_75t_R _15601_ (.A(_01144_),
    .B(_08497_),
    .Y(_08519_));
 NOR2x1_ASAP7_75t_R _15602_ (.A(_08125_),
    .B(_08519_),
    .Y(_08520_));
 XNOR2x1_ASAP7_75t_R _15603_ (.B(_08520_),
    .Y(_08521_),
    .A(net85));
 NOR2x1_ASAP7_75t_R _15604_ (.A(_08203_),
    .B(_08521_),
    .Y(_08522_));
 AND2x2_ASAP7_75t_R _15605_ (.A(_08078_),
    .B(_08522_),
    .Y(_08523_));
 OA21x2_ASAP7_75t_R _15606_ (.A1(_01142_),
    .A2(_08486_),
    .B(_01146_),
    .Y(_08524_));
 OA21x2_ASAP7_75t_R _15607_ (.A1(_01145_),
    .A2(_08524_),
    .B(_01149_),
    .Y(_08525_));
 XOR2x2_ASAP7_75t_R _15608_ (.A(_01148_),
    .B(_08525_),
    .Y(_08526_));
 AND4x1_ASAP7_75t_R _15609_ (.A(_08196_),
    .B(_08197_),
    .C(_08140_),
    .D(_08526_),
    .Y(_08527_));
 INVx1_ASAP7_75t_R _15610_ (.A(_08521_),
    .Y(_08528_));
 AND3x1_ASAP7_75t_R _15611_ (.A(_08203_),
    .B(_08088_),
    .C(_08526_),
    .Y(_08529_));
 AO221x1_ASAP7_75t_R _15612_ (.A1(_08202_),
    .A2(_08528_),
    .B1(_08522_),
    .B2(_08080_),
    .C(_08529_),
    .Y(_08530_));
 OR3x4_ASAP7_75t_R _15613_ (.A(_08523_),
    .B(_08527_),
    .C(_08530_),
    .Y(_08531_));
 OA222x2_ASAP7_75t_R _15614_ (.A1(_08514_),
    .A2(_08103_),
    .B1(_08116_),
    .B2(_08518_),
    .C1(_08531_),
    .C2(_08107_),
    .Y(_01274_));
 OR3x2_ASAP7_75t_R _15615_ (.A(_01147_),
    .B(_08213_),
    .C(_08519_),
    .Y(_08532_));
 XNOR2x1_ASAP7_75t_R _15616_ (.B(_08532_),
    .Y(_08533_),
    .A(net86));
 AND2x2_ASAP7_75t_R _15617_ (.A(_08329_),
    .B(_08533_),
    .Y(_08534_));
 AND2x2_ASAP7_75t_R _15618_ (.A(_08078_),
    .B(_08534_),
    .Y(_08535_));
 OA21x2_ASAP7_75t_R _15619_ (.A1(_01145_),
    .A2(_08503_),
    .B(_01149_),
    .Y(_08536_));
 OA21x2_ASAP7_75t_R _15620_ (.A1(_01148_),
    .A2(_08536_),
    .B(_01152_),
    .Y(_08537_));
 XOR2x1_ASAP7_75t_R _15621_ (.A(_01151_),
    .Y(_08538_),
    .B(_08537_));
 AND4x1_ASAP7_75t_R _15622_ (.A(_08335_),
    .B(_08370_),
    .C(_08089_),
    .D(_08538_),
    .Y(_08539_));
 AND3x1_ASAP7_75t_R _15623_ (.A(_08341_),
    .B(_08067_),
    .C(_08538_),
    .Y(_08540_));
 AO221x1_ASAP7_75t_R _15624_ (.A1(_08320_),
    .A2(_08533_),
    .B1(_08534_),
    .B2(_08375_),
    .C(_08540_),
    .Y(_08541_));
 OR3x4_ASAP7_75t_R _15625_ (.A(_08535_),
    .B(_08539_),
    .C(_08541_),
    .Y(_08542_));
 AO21x1_ASAP7_75t_R _15626_ (.A1(\readdata[29] ),
    .A2(_08280_),
    .B(_08282_),
    .Y(_08543_));
 AO21x1_ASAP7_75t_R _15627_ (.A1(_08179_),
    .A2(_08543_),
    .B(_08304_),
    .Y(_08544_));
 OAI21x1_ASAP7_75t_R _15628_ (.A1(_08361_),
    .A2(net53),
    .B(_08544_),
    .Y(_08545_));
 BUFx6f_ASAP7_75t_R _15629_ (.A(_08545_),
    .Y(_08546_));
 AOI22x1_ASAP7_75t_R _15630_ (.A1(_00111_),
    .A2(_08402_),
    .B1(_08416_),
    .B2(_08546_),
    .Y(_08547_));
 OA21x2_ASAP7_75t_R _15631_ (.A1(_08422_),
    .A2(_08542_),
    .B(_08547_),
    .Y(_01275_));
 XOR2x2_ASAP7_75t_R _15632_ (.A(_01071_),
    .B(_01159_),
    .Y(_08548_));
 NAND2x1_ASAP7_75t_R _15633_ (.A(_08067_),
    .B(_08548_),
    .Y(_08549_));
 OR3x1_ASAP7_75t_R _15634_ (.A(_08350_),
    .B(_08352_),
    .C(_08549_),
    .Y(_08550_));
 OR3x1_ASAP7_75t_R _15635_ (.A(net87),
    .B(_03249_),
    .C(_03254_),
    .Y(_08551_));
 AO31x2_ASAP7_75t_R _15636_ (.A1(_08021_),
    .A2(_08048_),
    .A3(_08053_),
    .B(_08551_),
    .Y(_08552_));
 NAND2x1_ASAP7_75t_R _15637_ (.A(_03256_),
    .B(_08548_),
    .Y(_08553_));
 AO211x2_ASAP7_75t_R _15638_ (.A1(_08043_),
    .A2(_08065_),
    .B(_08553_),
    .C(_05467_),
    .Y(_08554_));
 OA21x2_ASAP7_75t_R _15639_ (.A1(net87),
    .A2(_08088_),
    .B(_08554_),
    .Y(_08555_));
 OA31x2_ASAP7_75t_R _15640_ (.A1(_08058_),
    .A2(_08060_),
    .A3(_08551_),
    .B1(_08555_),
    .Y(_08556_));
 OA211x2_ASAP7_75t_R _15641_ (.A1(_08084_),
    .A2(_08550_),
    .B(_08552_),
    .C(_08556_),
    .Y(_08557_));
 AO21x1_ASAP7_75t_R _15642_ (.A1(\readdata[2] ),
    .A2(_08361_),
    .B(_08105_),
    .Y(_08558_));
 AOI21x1_ASAP7_75t_R _15643_ (.A1(_08108_),
    .A2(net54),
    .B(_08558_),
    .Y(_08559_));
 AOI21x1_ASAP7_75t_R _15644_ (.A1(_08106_),
    .A2(_08557_),
    .B(_08559_),
    .Y(_08560_));
 NOR2x1_ASAP7_75t_R _15645_ (.A(_01009_),
    .B(_08103_),
    .Y(_08561_));
 AO21x1_ASAP7_75t_R _15646_ (.A1(_08103_),
    .A2(_08560_),
    .B(_08561_),
    .Y(_01276_));
 AO21x1_ASAP7_75t_R _15647_ (.A1(\readdata[30] ),
    .A2(_08280_),
    .B(_08282_),
    .Y(_08562_));
 AO21x1_ASAP7_75t_R _15648_ (.A1(_08151_),
    .A2(_08562_),
    .B(_08304_),
    .Y(_08563_));
 OA211x2_ASAP7_75t_R _15649_ (.A1(_08149_),
    .A2(net55),
    .B(_08113_),
    .C(_08563_),
    .Y(_08564_));
 BUFx4f_ASAP7_75t_R _15650_ (.A(_08564_),
    .Y(_08565_));
 OR4x1_ASAP7_75t_R _15651_ (.A(_01147_),
    .B(_01150_),
    .C(_08125_),
    .D(_08519_),
    .Y(_08566_));
 XNOR2x1_ASAP7_75t_R _15652_ (.B(_08566_),
    .Y(_08567_),
    .A(net88));
 AND2x2_ASAP7_75t_R _15653_ (.A(_05776_),
    .B(_08567_),
    .Y(_08568_));
 AND2x2_ASAP7_75t_R _15654_ (.A(_08078_),
    .B(_08568_),
    .Y(_08569_));
 OA21x2_ASAP7_75t_R _15655_ (.A1(_01148_),
    .A2(_08525_),
    .B(_01152_),
    .Y(_08570_));
 OA21x2_ASAP7_75t_R _15656_ (.A1(_01151_),
    .A2(_08570_),
    .B(_01155_),
    .Y(_08571_));
 XOR2x2_ASAP7_75t_R _15657_ (.A(_01154_),
    .B(_08571_),
    .Y(_08572_));
 AND4x1_ASAP7_75t_R _15658_ (.A(_08196_),
    .B(_08197_),
    .C(_08089_),
    .D(_08572_),
    .Y(_08573_));
 AND2x2_ASAP7_75t_R _15659_ (.A(_08203_),
    .B(_08088_),
    .Y(_08574_));
 AO222x2_ASAP7_75t_R _15660_ (.A1(_08202_),
    .A2(_08567_),
    .B1(_08574_),
    .B2(_08572_),
    .C1(_08568_),
    .C2(_08080_),
    .Y(_08575_));
 OR3x4_ASAP7_75t_R _15661_ (.A(_08569_),
    .B(_08573_),
    .C(_08575_),
    .Y(_08576_));
 BUFx6f_ASAP7_75t_R _15662_ (.A(_08106_),
    .Y(_08577_));
 AND3x1_ASAP7_75t_R _15663_ (.A(_08145_),
    .B(_08146_),
    .C(_08577_),
    .Y(_08578_));
 NOR2x1_ASAP7_75t_R _15664_ (.A(_00077_),
    .B(_08103_),
    .Y(_08579_));
 AO221x1_ASAP7_75t_R _15665_ (.A1(_08103_),
    .A2(_08565_),
    .B1(_08576_),
    .B2(_08578_),
    .C(_08579_),
    .Y(_01277_));
 OR3x1_ASAP7_75t_R _15666_ (.A(_01150_),
    .B(_01153_),
    .C(_08532_),
    .Y(_08580_));
 XNOR2x1_ASAP7_75t_R _15667_ (.B(_08580_),
    .Y(_08581_),
    .A(_03025_));
 AND2x2_ASAP7_75t_R _15668_ (.A(_05776_),
    .B(_08581_),
    .Y(_08582_));
 OA21x2_ASAP7_75t_R _15669_ (.A1(_01151_),
    .A2(_08537_),
    .B(_01155_),
    .Y(_08583_));
 OA21x2_ASAP7_75t_R _15670_ (.A1(_01154_),
    .A2(_08583_),
    .B(_01156_),
    .Y(_08584_));
 OR2x2_ASAP7_75t_R _15671_ (.A(_09561_),
    .B(_07888_),
    .Y(_08585_));
 XNOR2x1_ASAP7_75t_R _15672_ (.B(_08585_),
    .Y(_08586_),
    .A(_03642_));
 XNOR2x2_ASAP7_75t_R _15673_ (.A(_08584_),
    .B(_08586_),
    .Y(_08587_));
 AND4x1_ASAP7_75t_R _15674_ (.A(_08196_),
    .B(_08197_),
    .C(_08089_),
    .D(_08587_),
    .Y(_08588_));
 AO222x2_ASAP7_75t_R _15675_ (.A1(_08574_),
    .A2(_08587_),
    .B1(_08581_),
    .B2(_08082_),
    .C1(_08080_),
    .C2(_08582_),
    .Y(_08589_));
 AOI211x1_ASAP7_75t_R _15676_ (.A1(_08084_),
    .A2(_08582_),
    .B(_08588_),
    .C(_08589_),
    .Y(_08590_));
 BUFx6f_ASAP7_75t_R _15677_ (.A(_08590_),
    .Y(_08591_));
 AO21x1_ASAP7_75t_R _15678_ (.A1(\readdata[31] ),
    .A2(_08281_),
    .B(_08283_),
    .Y(_08592_));
 AO21x1_ASAP7_75t_R _15679_ (.A1(_08188_),
    .A2(_08592_),
    .B(_08182_),
    .Y(_08593_));
 OAI21x1_ASAP7_75t_R _15680_ (.A1(_08150_),
    .A2(net56),
    .B(_08593_),
    .Y(_08594_));
 AND2x2_ASAP7_75t_R _15681_ (.A(_00045_),
    .B(_08402_),
    .Y(_08595_));
 AOI221x1_ASAP7_75t_R _15682_ (.A1(_08578_),
    .A2(_08591_),
    .B1(_08594_),
    .B2(_08148_),
    .C(_08595_),
    .Y(_01278_));
 AND2x2_ASAP7_75t_R _15683_ (.A(_01217_),
    .B(_05777_),
    .Y(_08596_));
 XNOR2x2_ASAP7_75t_R _15684_ (.A(_01073_),
    .B(_08165_),
    .Y(_08597_));
 AND3x1_ASAP7_75t_R _15685_ (.A(_08063_),
    .B(_08140_),
    .C(_08597_),
    .Y(_08598_));
 AO221x1_ASAP7_75t_R _15686_ (.A1(_01217_),
    .A2(_08082_),
    .B1(_08596_),
    .B2(_08087_),
    .C(_08598_),
    .Y(_08599_));
 AND4x1_ASAP7_75t_R _15687_ (.A(_08055_),
    .B(_08062_),
    .C(_08068_),
    .D(_08597_),
    .Y(_08600_));
 AOI211x1_ASAP7_75t_R _15688_ (.A1(_08084_),
    .A2(_08596_),
    .B(_08599_),
    .C(_08600_),
    .Y(_08601_));
 AND3x1_ASAP7_75t_R _15689_ (.A(\readdata[3] ),
    .B(_03222_),
    .C(_03224_),
    .Y(_08602_));
 AOI21x1_ASAP7_75t_R _15690_ (.A1(_08108_),
    .A2(net57),
    .B(_08602_),
    .Y(_08603_));
 BUFx6f_ASAP7_75t_R _15691_ (.A(_08603_),
    .Y(_08604_));
 AOI22x1_ASAP7_75t_R _15692_ (.A1(_00976_),
    .A2(_08402_),
    .B1(_08416_),
    .B2(_08604_),
    .Y(_08605_));
 OA21x2_ASAP7_75t_R _15693_ (.A1(_08422_),
    .A2(_08601_),
    .B(_08605_),
    .Y(_01279_));
 BUFx16f_ASAP7_75t_R _15694_ (.A(_08105_),
    .Y(_08606_));
 AND3x1_ASAP7_75t_R _15695_ (.A(\readdata[4] ),
    .B(_03222_),
    .C(_03224_),
    .Y(_08607_));
 AO21x2_ASAP7_75t_R _15696_ (.A1(_08108_),
    .A2(net58),
    .B(_08607_),
    .Y(_08608_));
 OR2x6_ASAP7_75t_R _15697_ (.A(_08606_),
    .B(_08608_),
    .Y(_08609_));
 XOR2x1_ASAP7_75t_R _15698_ (.A(_01075_),
    .Y(_08610_),
    .B(_01218_));
 OR3x1_ASAP7_75t_R _15699_ (.A(_03249_),
    .B(_03254_),
    .C(_08610_),
    .Y(_08611_));
 XOR2x1_ASAP7_75t_R _15700_ (.A(_01076_),
    .Y(_08612_),
    .B(_08130_));
 OR4x1_ASAP7_75t_R _15701_ (.A(_08077_),
    .B(_08079_),
    .C(_08081_),
    .D(_08612_),
    .Y(_08613_));
 OR3x1_ASAP7_75t_R _15702_ (.A(_05775_),
    .B(_08081_),
    .C(_08612_),
    .Y(_08614_));
 OA21x2_ASAP7_75t_R _15703_ (.A1(_08088_),
    .A2(_08610_),
    .B(_08614_),
    .Y(_08615_));
 OA21x2_ASAP7_75t_R _15704_ (.A1(_08197_),
    .A2(_08611_),
    .B(_08615_),
    .Y(_08616_));
 OA211x2_ASAP7_75t_R _15705_ (.A1(_08055_),
    .A2(_08611_),
    .B(_08613_),
    .C(_08616_),
    .Y(_08617_));
 BUFx10_ASAP7_75t_R _15706_ (.A(_08617_),
    .Y(_08618_));
 BUFx6f_ASAP7_75t_R _15707_ (.A(_08618_),
    .Y(_08619_));
 NAND2x1_ASAP7_75t_R _15708_ (.A(_00943_),
    .B(_08402_),
    .Y(_08620_));
 OA221x2_ASAP7_75t_R _15709_ (.A1(_08144_),
    .A2(_08609_),
    .B1(_08619_),
    .B2(_08107_),
    .C(_08620_),
    .Y(_01280_));
 XNOR2x1_ASAP7_75t_R _15710_ (.B(_08158_),
    .Y(_08621_),
    .A(net92));
 AND2x2_ASAP7_75t_R _15711_ (.A(_05776_),
    .B(_08621_),
    .Y(_08622_));
 AND2x2_ASAP7_75t_R _15712_ (.A(_08077_),
    .B(_08622_),
    .Y(_08623_));
 XOR2x2_ASAP7_75t_R _15713_ (.A(_01079_),
    .B(_08168_),
    .Y(_08624_));
 AND4x1_ASAP7_75t_R _15714_ (.A(_08196_),
    .B(_08197_),
    .C(_08140_),
    .D(_08624_),
    .Y(_08625_));
 AND3x1_ASAP7_75t_R _15715_ (.A(_08203_),
    .B(_08088_),
    .C(_08624_),
    .Y(_08626_));
 AO221x1_ASAP7_75t_R _15716_ (.A1(_08202_),
    .A2(_08621_),
    .B1(_08622_),
    .B2(_08080_),
    .C(_08626_),
    .Y(_08627_));
 OR3x4_ASAP7_75t_R _15717_ (.A(_08623_),
    .B(_08625_),
    .C(_08627_),
    .Y(_08628_));
 AND3x1_ASAP7_75t_R _15718_ (.A(\readdata[5] ),
    .B(_03222_),
    .C(_03224_),
    .Y(_08629_));
 AO211x2_ASAP7_75t_R _15719_ (.A1(_08108_),
    .A2(net59),
    .B(_08106_),
    .C(_08629_),
    .Y(_08630_));
 BUFx6f_ASAP7_75t_R _15720_ (.A(_08630_),
    .Y(_08631_));
 NAND2x1_ASAP7_75t_R _15721_ (.A(_00909_),
    .B(_08402_),
    .Y(_08632_));
 OA221x2_ASAP7_75t_R _15722_ (.A1(_08107_),
    .A2(_08628_),
    .B1(_08631_),
    .B2(_08144_),
    .C(_08632_),
    .Y(_01281_));
 XNOR2x1_ASAP7_75t_R _15723_ (.B(_08123_),
    .Y(_08633_),
    .A(net93));
 AND2x2_ASAP7_75t_R _15724_ (.A(_08329_),
    .B(_08633_),
    .Y(_08634_));
 AND2x2_ASAP7_75t_R _15725_ (.A(_08078_),
    .B(_08634_),
    .Y(_08635_));
 OA21x2_ASAP7_75t_R _15726_ (.A1(_01079_),
    .A2(_08131_),
    .B(_01083_),
    .Y(_08636_));
 XOR2x2_ASAP7_75t_R _15727_ (.A(_01082_),
    .B(_08636_),
    .Y(_08637_));
 AND4x1_ASAP7_75t_R _15728_ (.A(_08335_),
    .B(_08370_),
    .C(_08089_),
    .D(_08637_),
    .Y(_08638_));
 AND3x1_ASAP7_75t_R _15729_ (.A(_08341_),
    .B(_08067_),
    .C(_08637_),
    .Y(_08639_));
 AO221x1_ASAP7_75t_R _15730_ (.A1(_08202_),
    .A2(_08633_),
    .B1(_08634_),
    .B2(_08375_),
    .C(_08639_),
    .Y(_08640_));
 OR3x4_ASAP7_75t_R _15731_ (.A(_08635_),
    .B(_08638_),
    .C(_08640_),
    .Y(_08641_));
 AND3x1_ASAP7_75t_R _15732_ (.A(\readdata[6] ),
    .B(_03222_),
    .C(_03224_),
    .Y(_08642_));
 AOI21x1_ASAP7_75t_R _15733_ (.A1(_08108_),
    .A2(net60),
    .B(_08642_),
    .Y(_08643_));
 BUFx6f_ASAP7_75t_R _15734_ (.A(_08643_),
    .Y(_08644_));
 AOI22x1_ASAP7_75t_R _15735_ (.A1(_00876_),
    .A2(_08402_),
    .B1(_08416_),
    .B2(_08644_),
    .Y(_08645_));
 OA21x2_ASAP7_75t_R _15736_ (.A1(_08422_),
    .A2(_08641_),
    .B(_08645_),
    .Y(_01282_));
 NOR2x1_ASAP7_75t_R _15737_ (.A(_01081_),
    .B(_08159_),
    .Y(_08646_));
 XNOR2x1_ASAP7_75t_R _15738_ (.B(_08646_),
    .Y(_08647_),
    .A(_01084_));
 AND2x2_ASAP7_75t_R _15739_ (.A(_05776_),
    .B(_08647_),
    .Y(_08648_));
 AND2x2_ASAP7_75t_R _15740_ (.A(_08078_),
    .B(_08648_),
    .Y(_08649_));
 XOR2x2_ASAP7_75t_R _15741_ (.A(_01085_),
    .B(_08169_),
    .Y(_08650_));
 AND4x1_ASAP7_75t_R _15742_ (.A(_08196_),
    .B(_08370_),
    .C(_08089_),
    .D(_08650_),
    .Y(_08651_));
 AND3x1_ASAP7_75t_R _15743_ (.A(_08203_),
    .B(_08067_),
    .C(_08650_),
    .Y(_08652_));
 AO221x1_ASAP7_75t_R _15744_ (.A1(_08202_),
    .A2(_08647_),
    .B1(_08648_),
    .B2(_08375_),
    .C(_08652_),
    .Y(_08653_));
 OR3x4_ASAP7_75t_R _15745_ (.A(_08649_),
    .B(_08651_),
    .C(_08653_),
    .Y(_08654_));
 AND2x2_ASAP7_75t_R _15746_ (.A(_06935_),
    .B(_07336_),
    .Y(_08655_));
 AO221x2_ASAP7_75t_R _15747_ (.A1(\readdata[7] ),
    .A2(_08149_),
    .B1(_07328_),
    .B2(_08655_),
    .C(_08105_),
    .Y(_08656_));
 NAND2x1_ASAP7_75t_R _15748_ (.A(_00842_),
    .B(_08118_),
    .Y(_08657_));
 OA21x2_ASAP7_75t_R _15749_ (.A1(_08402_),
    .A2(_08656_),
    .B(_08657_),
    .Y(_08658_));
 OA21x2_ASAP7_75t_R _15750_ (.A1(_08422_),
    .A2(_08654_),
    .B(_08658_),
    .Y(_01283_));
 OR3x1_ASAP7_75t_R _15751_ (.A(_01081_),
    .B(_01084_),
    .C(_08123_),
    .Y(_08659_));
 XNOR2x1_ASAP7_75t_R _15752_ (.B(_08659_),
    .Y(_08660_),
    .A(net95));
 AND2x2_ASAP7_75t_R _15753_ (.A(_05776_),
    .B(_08660_),
    .Y(_08661_));
 AND2x2_ASAP7_75t_R _15754_ (.A(_08078_),
    .B(_08661_),
    .Y(_08662_));
 XOR2x2_ASAP7_75t_R _15755_ (.A(_01088_),
    .B(_08135_),
    .Y(_08663_));
 AND4x1_ASAP7_75t_R _15756_ (.A(_08196_),
    .B(_08197_),
    .C(_08089_),
    .D(_08663_),
    .Y(_08664_));
 AND3x1_ASAP7_75t_R _15757_ (.A(_08203_),
    .B(_08067_),
    .C(_08663_),
    .Y(_08665_));
 AO221x1_ASAP7_75t_R _15758_ (.A1(_08202_),
    .A2(_08660_),
    .B1(_08661_),
    .B2(_08080_),
    .C(_08665_),
    .Y(_08666_));
 OR3x4_ASAP7_75t_R _15759_ (.A(_08662_),
    .B(_08664_),
    .C(_08666_),
    .Y(_08667_));
 AO21x1_ASAP7_75t_R _15760_ (.A1(\readdata[8] ),
    .A2(_08179_),
    .B(_08304_),
    .Y(_08668_));
 OAI21x1_ASAP7_75t_R _15761_ (.A1(_08361_),
    .A2(net62),
    .B(_08668_),
    .Y(_08669_));
 BUFx6f_ASAP7_75t_R _15762_ (.A(_08669_),
    .Y(_08670_));
 AOI22x1_ASAP7_75t_R _15763_ (.A1(_00809_),
    .A2(_08402_),
    .B1(_08416_),
    .B2(_08670_),
    .Y(_08671_));
 OA21x2_ASAP7_75t_R _15764_ (.A1(_08422_),
    .A2(_08667_),
    .B(_08671_),
    .Y(_01284_));
 OR4x1_ASAP7_75t_R _15765_ (.A(_01081_),
    .B(_01084_),
    .C(_01087_),
    .D(_08159_),
    .Y(_08672_));
 XNOR2x1_ASAP7_75t_R _15766_ (.B(_08672_),
    .Y(_08673_),
    .A(net96));
 AND2x2_ASAP7_75t_R _15767_ (.A(_05776_),
    .B(_08673_),
    .Y(_08674_));
 AND2x2_ASAP7_75t_R _15768_ (.A(_08078_),
    .B(_08674_),
    .Y(_08675_));
 XOR2x1_ASAP7_75t_R _15769_ (.A(_01091_),
    .Y(_08676_),
    .B(_08171_));
 AND4x1_ASAP7_75t_R _15770_ (.A(_08196_),
    .B(_08197_),
    .C(_08089_),
    .D(_08676_),
    .Y(_08677_));
 AND3x1_ASAP7_75t_R _15771_ (.A(_08203_),
    .B(_08067_),
    .C(_08676_),
    .Y(_08678_));
 AO221x1_ASAP7_75t_R _15772_ (.A1(_08202_),
    .A2(_08673_),
    .B1(_08674_),
    .B2(_08080_),
    .C(_08678_),
    .Y(_08679_));
 OR3x4_ASAP7_75t_R _15773_ (.A(_08675_),
    .B(_08677_),
    .C(_08679_),
    .Y(_08680_));
 NAND2x1_ASAP7_75t_R _15774_ (.A(_06935_),
    .B(_08112_),
    .Y(_08681_));
 AO21x1_ASAP7_75t_R _15775_ (.A1(\readdata[9] ),
    .A2(_08151_),
    .B(_08152_),
    .Y(_08682_));
 OA22x2_ASAP7_75t_R _15776_ (.A1(_07373_),
    .A2(_08681_),
    .B1(_08682_),
    .B2(_06935_),
    .Y(_08683_));
 OA21x2_ASAP7_75t_R _15777_ (.A1(_07392_),
    .A2(_08681_),
    .B(_08683_),
    .Y(_08684_));
 NAND2x1_ASAP7_75t_R _15778_ (.A(_00775_),
    .B(_08118_),
    .Y(_08685_));
 OA21x2_ASAP7_75t_R _15779_ (.A1(_08402_),
    .A2(_08684_),
    .B(_08685_),
    .Y(_08686_));
 OA21x2_ASAP7_75t_R _15780_ (.A1(_08107_),
    .A2(_08680_),
    .B(_08686_),
    .Y(_01285_));
 BUFx16f_ASAP7_75t_R _15781_ (.A(_08105_),
    .Y(_08687_));
 AND3x2_ASAP7_75t_R _15782_ (.A(_03279_),
    .B(_06715_),
    .C(_08096_),
    .Y(_08688_));
 BUFx16f_ASAP7_75t_R _15783_ (.A(_08688_),
    .Y(_08689_));
 AND2x6_ASAP7_75t_R _15784_ (.A(_08102_),
    .B(_08689_),
    .Y(_08690_));
 NAND2x2_ASAP7_75t_R _15785_ (.A(_08687_),
    .B(_08690_),
    .Y(_08691_));
 BUFx4f_ASAP7_75t_R _15786_ (.A(_08691_),
    .Y(_08692_));
 NAND2x2_ASAP7_75t_R _15787_ (.A(_08115_),
    .B(_08690_),
    .Y(_08693_));
 BUFx16f_ASAP7_75t_R _15788_ (.A(_08689_),
    .Y(_08694_));
 NAND2x2_ASAP7_75t_R _15789_ (.A(_08102_),
    .B(_08694_),
    .Y(_08695_));
 BUFx6f_ASAP7_75t_R _15790_ (.A(_08695_),
    .Y(_08696_));
 NAND2x1_ASAP7_75t_R _15791_ (.A(_00011_),
    .B(_08696_),
    .Y(_08697_));
 OA21x2_ASAP7_75t_R _15792_ (.A1(_08111_),
    .A2(_08693_),
    .B(_08697_),
    .Y(_08698_));
 OA21x2_ASAP7_75t_R _15793_ (.A1(_08093_),
    .A2(_08692_),
    .B(_08698_),
    .Y(_01286_));
 BUFx4f_ASAP7_75t_R _15794_ (.A(_08143_),
    .Y(_08699_));
 BUFx10_ASAP7_75t_R _15795_ (.A(_08695_),
    .Y(_08700_));
 BUFx6f_ASAP7_75t_R _15796_ (.A(_08113_),
    .Y(_08701_));
 AND3x2_ASAP7_75t_R _15797_ (.A(_08146_),
    .B(_08701_),
    .C(_08694_),
    .Y(_08702_));
 BUFx10_ASAP7_75t_R _15798_ (.A(_08702_),
    .Y(_08703_));
 AOI22x1_ASAP7_75t_R _15799_ (.A1(_00743_),
    .A2(_08700_),
    .B1(_08703_),
    .B2(_08156_),
    .Y(_08704_));
 OA21x2_ASAP7_75t_R _15800_ (.A1(_08699_),
    .A2(_08692_),
    .B(_08704_),
    .Y(_01287_));
 BUFx4f_ASAP7_75t_R _15801_ (.A(_08178_),
    .Y(_08705_));
 AOI22x1_ASAP7_75t_R _15802_ (.A1(_00710_),
    .A2(_08700_),
    .B1(_08703_),
    .B2(_08185_),
    .Y(_08706_));
 OA21x2_ASAP7_75t_R _15803_ (.A1(_08705_),
    .A2(_08692_),
    .B(_08706_),
    .Y(_01288_));
 BUFx3_ASAP7_75t_R _15804_ (.A(_08206_),
    .Y(_08707_));
 OA222x2_ASAP7_75t_R _15805_ (.A1(_05737_),
    .A2(_08690_),
    .B1(_08691_),
    .B2(_08707_),
    .C1(_08693_),
    .C2(_08191_),
    .Y(_01289_));
 INVx1_ASAP7_75t_R _15806_ (.A(_00644_),
    .Y(_08708_));
 BUFx3_ASAP7_75t_R _15807_ (.A(_08224_),
    .Y(_08709_));
 OA222x2_ASAP7_75t_R _15808_ (.A1(_08708_),
    .A2(_08690_),
    .B1(_08691_),
    .B2(_08709_),
    .C1(_08693_),
    .C2(_08211_),
    .Y(_01290_));
 BUFx4f_ASAP7_75t_R _15809_ (.A(_08240_),
    .Y(_08710_));
 AOI22x1_ASAP7_75t_R _15810_ (.A1(_00611_),
    .A2(_08700_),
    .B1(_08703_),
    .B2(_08243_),
    .Y(_08711_));
 OA21x2_ASAP7_75t_R _15811_ (.A1(_08710_),
    .A2(_08692_),
    .B(_08711_),
    .Y(_01291_));
 BUFx4f_ASAP7_75t_R _15812_ (.A(_08256_),
    .Y(_08712_));
 AOI22x1_ASAP7_75t_R _15813_ (.A1(_00577_),
    .A2(_08700_),
    .B1(_08703_),
    .B2(_08259_),
    .Y(_08713_));
 OA21x2_ASAP7_75t_R _15814_ (.A1(_08712_),
    .A2(_08692_),
    .B(_08713_),
    .Y(_01292_));
 BUFx4f_ASAP7_75t_R _15815_ (.A(_08279_),
    .Y(_08714_));
 AOI22x1_ASAP7_75t_R _15816_ (.A1(_00544_),
    .A2(_08700_),
    .B1(_08703_),
    .B2(_08287_),
    .Y(_08715_));
 OA21x2_ASAP7_75t_R _15817_ (.A1(_08714_),
    .A2(_08692_),
    .B(_08715_),
    .Y(_01293_));
 BUFx3_ASAP7_75t_R _15818_ (.A(_08301_),
    .Y(_08716_));
 BUFx12_ASAP7_75t_R _15819_ (.A(_08695_),
    .Y(_08717_));
 AOI22x1_ASAP7_75t_R _15820_ (.A1(_00511_),
    .A2(_08717_),
    .B1(_08703_),
    .B2(_08308_),
    .Y(_08718_));
 OA21x2_ASAP7_75t_R _15821_ (.A1(_08716_),
    .A2(_08692_),
    .B(_08718_),
    .Y(_01294_));
 BUFx3_ASAP7_75t_R _15822_ (.A(_08323_),
    .Y(_08719_));
 AOI22x1_ASAP7_75t_R _15823_ (.A1(_00478_),
    .A2(_08717_),
    .B1(_08703_),
    .B2(_08327_),
    .Y(_08720_));
 OA21x2_ASAP7_75t_R _15824_ (.A1(_08719_),
    .A2(_08692_),
    .B(_08720_),
    .Y(_01295_));
 BUFx3_ASAP7_75t_R _15825_ (.A(_08344_),
    .Y(_08721_));
 AOI22x1_ASAP7_75t_R _15826_ (.A1(_00445_),
    .A2(_08717_),
    .B1(_08703_),
    .B2(_08348_),
    .Y(_08722_));
 OA21x2_ASAP7_75t_R _15827_ (.A1(_08721_),
    .A2(_08692_),
    .B(_08722_),
    .Y(_01296_));
 BUFx4f_ASAP7_75t_R _15828_ (.A(_08364_),
    .Y(_08723_));
 NAND2x1_ASAP7_75t_R _15829_ (.A(_01043_),
    .B(_08700_),
    .Y(_08724_));
 OA21x2_ASAP7_75t_R _15830_ (.A1(_08723_),
    .A2(_08700_),
    .B(_08724_),
    .Y(_01297_));
 BUFx3_ASAP7_75t_R _15831_ (.A(_08378_),
    .Y(_08725_));
 AOI22x1_ASAP7_75t_R _15832_ (.A1(_00412_),
    .A2(_08717_),
    .B1(_08703_),
    .B2(_08382_),
    .Y(_08726_));
 OA21x2_ASAP7_75t_R _15833_ (.A1(_08725_),
    .A2(_08692_),
    .B(_08726_),
    .Y(_01298_));
 BUFx6f_ASAP7_75t_R _15834_ (.A(_08396_),
    .Y(_08727_));
 NAND2x1_ASAP7_75t_R _15835_ (.A(_00379_),
    .B(_08696_),
    .Y(_08728_));
 OA221x2_ASAP7_75t_R _15836_ (.A1(_08401_),
    .A2(_08700_),
    .B1(_08691_),
    .B2(_08727_),
    .C(_08728_),
    .Y(_01299_));
 BUFx3_ASAP7_75t_R _15837_ (.A(_08415_),
    .Y(_08729_));
 BUFx4f_ASAP7_75t_R _15838_ (.A(_08691_),
    .Y(_08730_));
 BUFx6f_ASAP7_75t_R _15839_ (.A(_08702_),
    .Y(_08731_));
 AOI22x1_ASAP7_75t_R _15840_ (.A1(_00346_),
    .A2(_08717_),
    .B1(_08731_),
    .B2(_08420_),
    .Y(_08732_));
 OA21x2_ASAP7_75t_R _15841_ (.A1(_08729_),
    .A2(_08730_),
    .B(_08732_),
    .Y(_01300_));
 BUFx3_ASAP7_75t_R _15842_ (.A(_08434_),
    .Y(_08733_));
 AOI22x1_ASAP7_75t_R _15843_ (.A1(_00312_),
    .A2(_08717_),
    .B1(_08731_),
    .B2(_08438_),
    .Y(_08734_));
 OA21x2_ASAP7_75t_R _15844_ (.A1(_08733_),
    .A2(_08730_),
    .B(_08734_),
    .Y(_01301_));
 BUFx4f_ASAP7_75t_R _15845_ (.A(_08455_),
    .Y(_08735_));
 AOI22x1_ASAP7_75t_R _15846_ (.A1(_00279_),
    .A2(_08717_),
    .B1(_08731_),
    .B2(_08459_),
    .Y(_08736_));
 OA21x2_ASAP7_75t_R _15847_ (.A1(_08735_),
    .A2(_08730_),
    .B(_08736_),
    .Y(_01302_));
 BUFx4f_ASAP7_75t_R _15848_ (.A(_08472_),
    .Y(_08737_));
 AOI22x1_ASAP7_75t_R _15849_ (.A1(_00246_),
    .A2(_08717_),
    .B1(_08731_),
    .B2(_08477_),
    .Y(_08738_));
 OA21x2_ASAP7_75t_R _15850_ (.A1(_08737_),
    .A2(_08730_),
    .B(_08738_),
    .Y(_01303_));
 BUFx4f_ASAP7_75t_R _15851_ (.A(_08491_),
    .Y(_08739_));
 AOI22x1_ASAP7_75t_R _15852_ (.A1(_00212_),
    .A2(_08717_),
    .B1(_08731_),
    .B2(_08495_),
    .Y(_08740_));
 OA21x2_ASAP7_75t_R _15853_ (.A1(_08739_),
    .A2(_08730_),
    .B(_08740_),
    .Y(_01304_));
 BUFx4f_ASAP7_75t_R _15854_ (.A(_08508_),
    .Y(_08741_));
 AOI22x1_ASAP7_75t_R _15855_ (.A1(_00179_),
    .A2(_08717_),
    .B1(_08731_),
    .B2(_08512_),
    .Y(_08742_));
 OA21x2_ASAP7_75t_R _15856_ (.A1(_08741_),
    .A2(_08730_),
    .B(_08742_),
    .Y(_01305_));
 INVx1_ASAP7_75t_R _15857_ (.A(_00145_),
    .Y(_08743_));
 BUFx4f_ASAP7_75t_R _15858_ (.A(_08531_),
    .Y(_08744_));
 OA222x2_ASAP7_75t_R _15859_ (.A1(_08743_),
    .A2(_08690_),
    .B1(_08691_),
    .B2(_08744_),
    .C1(_08693_),
    .C2(_08518_),
    .Y(_01306_));
 BUFx4f_ASAP7_75t_R _15860_ (.A(_08542_),
    .Y(_08745_));
 AOI22x1_ASAP7_75t_R _15861_ (.A1(_00112_),
    .A2(_08696_),
    .B1(_08731_),
    .B2(_08546_),
    .Y(_08746_));
 OA21x2_ASAP7_75t_R _15862_ (.A1(_08745_),
    .A2(_08730_),
    .B(_08746_),
    .Y(_01307_));
 BUFx4f_ASAP7_75t_R _15863_ (.A(_08560_),
    .Y(_08747_));
 NOR2x1_ASAP7_75t_R _15864_ (.A(_01010_),
    .B(_08690_),
    .Y(_08748_));
 AO21x1_ASAP7_75t_R _15865_ (.A1(_08747_),
    .A2(_08690_),
    .B(_08748_),
    .Y(_01308_));
 BUFx10_ASAP7_75t_R _15866_ (.A(_08689_),
    .Y(_08749_));
 BUFx6f_ASAP7_75t_R _15867_ (.A(_08749_),
    .Y(_08750_));
 AND3x1_ASAP7_75t_R _15868_ (.A(_08146_),
    .B(_08577_),
    .C(_08750_),
    .Y(_08751_));
 BUFx3_ASAP7_75t_R _15869_ (.A(_08576_),
    .Y(_08752_));
 NOR2x1_ASAP7_75t_R _15870_ (.A(_00078_),
    .B(_08690_),
    .Y(_08753_));
 AO221x1_ASAP7_75t_R _15871_ (.A1(_08565_),
    .A2(_08690_),
    .B1(_08751_),
    .B2(_08752_),
    .C(_08753_),
    .Y(_01309_));
 BUFx6f_ASAP7_75t_R _15872_ (.A(_08594_),
    .Y(_08754_));
 AND2x2_ASAP7_75t_R _15873_ (.A(_00046_),
    .B(_08696_),
    .Y(_08755_));
 AOI221x1_ASAP7_75t_R _15874_ (.A1(_08591_),
    .A2(_08751_),
    .B1(_08703_),
    .B2(_08754_),
    .C(_08755_),
    .Y(_01310_));
 BUFx4f_ASAP7_75t_R _15875_ (.A(_08601_),
    .Y(_08756_));
 AOI22x1_ASAP7_75t_R _15876_ (.A1(_00977_),
    .A2(_08696_),
    .B1(_08731_),
    .B2(_08604_),
    .Y(_08757_));
 OA21x2_ASAP7_75t_R _15877_ (.A1(_08756_),
    .A2(_08730_),
    .B(_08757_),
    .Y(_01311_));
 BUFx6f_ASAP7_75t_R _15878_ (.A(_08609_),
    .Y(_08758_));
 AO21x1_ASAP7_75t_R _15879_ (.A1(_08146_),
    .A2(_08750_),
    .B(_06491_),
    .Y(_08759_));
 OA221x2_ASAP7_75t_R _15880_ (.A1(_08758_),
    .A2(_08700_),
    .B1(_08691_),
    .B2(_08619_),
    .C(_08759_),
    .Y(_01312_));
 BUFx6f_ASAP7_75t_R _15881_ (.A(_08628_),
    .Y(_08760_));
 NAND2x1_ASAP7_75t_R _15882_ (.A(_00910_),
    .B(_08696_),
    .Y(_08761_));
 OA221x2_ASAP7_75t_R _15883_ (.A1(_08631_),
    .A2(_08700_),
    .B1(_08691_),
    .B2(_08760_),
    .C(_08761_),
    .Y(_01313_));
 BUFx4f_ASAP7_75t_R _15884_ (.A(_08641_),
    .Y(_08762_));
 AOI22x1_ASAP7_75t_R _15885_ (.A1(_00877_),
    .A2(_08696_),
    .B1(_08731_),
    .B2(_08644_),
    .Y(_08763_));
 OA21x2_ASAP7_75t_R _15886_ (.A1(_08762_),
    .A2(_08730_),
    .B(_08763_),
    .Y(_01314_));
 BUFx4f_ASAP7_75t_R _15887_ (.A(_08654_),
    .Y(_08764_));
 BUFx4f_ASAP7_75t_R _15888_ (.A(_08656_),
    .Y(_08765_));
 NAND2x1_ASAP7_75t_R _15889_ (.A(_00843_),
    .B(_08695_),
    .Y(_08766_));
 OA21x2_ASAP7_75t_R _15890_ (.A1(_08765_),
    .A2(_08696_),
    .B(_08766_),
    .Y(_08767_));
 OA21x2_ASAP7_75t_R _15891_ (.A1(_08764_),
    .A2(_08730_),
    .B(_08767_),
    .Y(_01315_));
 BUFx4f_ASAP7_75t_R _15892_ (.A(_08667_),
    .Y(_08768_));
 AOI22x1_ASAP7_75t_R _15893_ (.A1(_00810_),
    .A2(_08696_),
    .B1(_08731_),
    .B2(_08670_),
    .Y(_08769_));
 OA21x2_ASAP7_75t_R _15894_ (.A1(_08768_),
    .A2(_08691_),
    .B(_08769_),
    .Y(_01316_));
 BUFx4f_ASAP7_75t_R _15895_ (.A(_08680_),
    .Y(_08770_));
 BUFx4f_ASAP7_75t_R _15896_ (.A(_08684_),
    .Y(_08771_));
 NAND2x1_ASAP7_75t_R _15897_ (.A(_00776_),
    .B(_08695_),
    .Y(_08772_));
 OA21x2_ASAP7_75t_R _15898_ (.A1(_08771_),
    .A2(_08696_),
    .B(_08772_),
    .Y(_08773_));
 OA21x2_ASAP7_75t_R _15899_ (.A1(_08770_),
    .A2(_08691_),
    .B(_08773_),
    .Y(_01317_));
 AOI21x1_ASAP7_75t_R _15900_ (.A1(_03025_),
    .A2(net29),
    .B(_03238_),
    .Y(_08774_));
 NAND2x1_ASAP7_75t_R _15901_ (.A(_08774_),
    .B(_08096_),
    .Y(_08775_));
 OA21x2_ASAP7_75t_R _15902_ (.A1(net5),
    .A2(net2),
    .B(_03024_),
    .Y(_08776_));
 NOR2x2_ASAP7_75t_R _15903_ (.A(_06618_),
    .B(_08776_),
    .Y(_08777_));
 OR3x4_ASAP7_75t_R _15904_ (.A(_03279_),
    .B(_08775_),
    .C(_08777_),
    .Y(_08778_));
 INVx1_ASAP7_75t_R _15905_ (.A(net2),
    .Y(_08779_));
 OR4x2_ASAP7_75t_R _15906_ (.A(_03713_),
    .B(net5),
    .C(_08779_),
    .D(_08100_),
    .Y(_08780_));
 OR3x1_ASAP7_75t_R _15907_ (.A(_08113_),
    .B(_08778_),
    .C(_08780_),
    .Y(_08781_));
 BUFx6f_ASAP7_75t_R _15908_ (.A(_08781_),
    .Y(_08782_));
 BUFx6f_ASAP7_75t_R _15909_ (.A(_08782_),
    .Y(_08783_));
 INVx1_ASAP7_75t_R _15910_ (.A(_00012_),
    .Y(_08784_));
 INVx1_ASAP7_75t_R _15911_ (.A(_08777_),
    .Y(_08785_));
 AND4x2_ASAP7_75t_R _15912_ (.A(_08094_),
    .B(_08774_),
    .C(_08096_),
    .D(_08785_),
    .Y(_08786_));
 BUFx16f_ASAP7_75t_R _15913_ (.A(_08786_),
    .Y(_08787_));
 BUFx6f_ASAP7_75t_R _15914_ (.A(_08787_),
    .Y(_08788_));
 INVx6_ASAP7_75t_R _15915_ (.A(_08780_),
    .Y(_08789_));
 BUFx4f_ASAP7_75t_R _15916_ (.A(_08789_),
    .Y(_08790_));
 AND2x6_ASAP7_75t_R _15917_ (.A(_08788_),
    .B(_08790_),
    .Y(_08791_));
 OR3x2_ASAP7_75t_R _15918_ (.A(_08106_),
    .B(_08778_),
    .C(_08780_),
    .Y(_08792_));
 BUFx6f_ASAP7_75t_R _15919_ (.A(_08110_),
    .Y(_08793_));
 OA22x2_ASAP7_75t_R _15920_ (.A1(_08784_),
    .A2(_08791_),
    .B1(_08792_),
    .B2(_08793_),
    .Y(_08794_));
 OA21x2_ASAP7_75t_R _15921_ (.A1(_08093_),
    .A2(_08783_),
    .B(_08794_),
    .Y(_01318_));
 BUFx12f_ASAP7_75t_R _15922_ (.A(_08787_),
    .Y(_08795_));
 NAND2x2_ASAP7_75t_R _15923_ (.A(_08795_),
    .B(_08790_),
    .Y(_08796_));
 BUFx10_ASAP7_75t_R _15924_ (.A(_08796_),
    .Y(_08797_));
 BUFx6f_ASAP7_75t_R _15925_ (.A(_08113_),
    .Y(_08798_));
 AND3x2_ASAP7_75t_R _15926_ (.A(_08798_),
    .B(_08788_),
    .C(_08790_),
    .Y(_08799_));
 BUFx10_ASAP7_75t_R _15927_ (.A(_08799_),
    .Y(_08800_));
 AOI22x1_ASAP7_75t_R _15928_ (.A1(_00744_),
    .A2(_08797_),
    .B1(_08800_),
    .B2(_08156_),
    .Y(_08801_));
 OA21x2_ASAP7_75t_R _15929_ (.A1(_08699_),
    .A2(_08783_),
    .B(_08801_),
    .Y(_01319_));
 AOI22x1_ASAP7_75t_R _15930_ (.A1(_00711_),
    .A2(_08797_),
    .B1(_08800_),
    .B2(_08185_),
    .Y(_08802_));
 OA21x2_ASAP7_75t_R _15931_ (.A1(_08705_),
    .A2(_08783_),
    .B(_08802_),
    .Y(_01320_));
 OA222x2_ASAP7_75t_R _15932_ (.A1(_05732_),
    .A2(_08791_),
    .B1(_08782_),
    .B2(_08707_),
    .C1(_08792_),
    .C2(_08191_),
    .Y(_01321_));
 OA222x2_ASAP7_75t_R _15933_ (.A1(_05656_),
    .A2(_08791_),
    .B1(_08782_),
    .B2(_08709_),
    .C1(_08792_),
    .C2(_08211_),
    .Y(_01322_));
 AOI22x1_ASAP7_75t_R _15934_ (.A1(_00612_),
    .A2(_08797_),
    .B1(_08800_),
    .B2(_08243_),
    .Y(_08803_));
 OA21x2_ASAP7_75t_R _15935_ (.A1(_08710_),
    .A2(_08783_),
    .B(_08803_),
    .Y(_01323_));
 AOI22x1_ASAP7_75t_R _15936_ (.A1(_00578_),
    .A2(_08797_),
    .B1(_08800_),
    .B2(_08259_),
    .Y(_08804_));
 OA21x2_ASAP7_75t_R _15937_ (.A1(_08712_),
    .A2(_08783_),
    .B(_08804_),
    .Y(_01324_));
 AOI22x1_ASAP7_75t_R _15938_ (.A1(_00545_),
    .A2(_08797_),
    .B1(_08800_),
    .B2(_08287_),
    .Y(_08805_));
 OA21x2_ASAP7_75t_R _15939_ (.A1(_08714_),
    .A2(_08783_),
    .B(_08805_),
    .Y(_01325_));
 BUFx12_ASAP7_75t_R _15940_ (.A(_08796_),
    .Y(_08806_));
 AOI22x1_ASAP7_75t_R _15941_ (.A1(_00512_),
    .A2(_08806_),
    .B1(_08800_),
    .B2(_08308_),
    .Y(_08807_));
 OA21x2_ASAP7_75t_R _15942_ (.A1(_08716_),
    .A2(_08783_),
    .B(_08807_),
    .Y(_01326_));
 AOI22x1_ASAP7_75t_R _15943_ (.A1(_00479_),
    .A2(_08806_),
    .B1(_08800_),
    .B2(_08327_),
    .Y(_08808_));
 OA21x2_ASAP7_75t_R _15944_ (.A1(_08719_),
    .A2(_08783_),
    .B(_08808_),
    .Y(_01327_));
 AOI22x1_ASAP7_75t_R _15945_ (.A1(_00446_),
    .A2(_08806_),
    .B1(_08800_),
    .B2(_08348_),
    .Y(_08809_));
 OA21x2_ASAP7_75t_R _15946_ (.A1(_08721_),
    .A2(_08783_),
    .B(_08809_),
    .Y(_01328_));
 NAND2x1_ASAP7_75t_R _15947_ (.A(_01044_),
    .B(_08797_),
    .Y(_08810_));
 OA21x2_ASAP7_75t_R _15948_ (.A1(_08723_),
    .A2(_08797_),
    .B(_08810_),
    .Y(_01329_));
 AOI22x1_ASAP7_75t_R _15949_ (.A1(_00413_),
    .A2(_08806_),
    .B1(_08800_),
    .B2(_08382_),
    .Y(_08811_));
 OA21x2_ASAP7_75t_R _15950_ (.A1(_08725_),
    .A2(_08783_),
    .B(_08811_),
    .Y(_01330_));
 BUFx6f_ASAP7_75t_R _15951_ (.A(_08796_),
    .Y(_08812_));
 NAND2x1_ASAP7_75t_R _15952_ (.A(_00380_),
    .B(_08812_),
    .Y(_08813_));
 OA221x2_ASAP7_75t_R _15953_ (.A1(_08401_),
    .A2(_08797_),
    .B1(_08782_),
    .B2(_08727_),
    .C(_08813_),
    .Y(_01331_));
 BUFx4f_ASAP7_75t_R _15954_ (.A(_08782_),
    .Y(_08814_));
 BUFx6f_ASAP7_75t_R _15955_ (.A(_08799_),
    .Y(_08815_));
 AOI22x1_ASAP7_75t_R _15956_ (.A1(_00347_),
    .A2(_08806_),
    .B1(_08815_),
    .B2(_08420_),
    .Y(_08816_));
 OA21x2_ASAP7_75t_R _15957_ (.A1(_08729_),
    .A2(_08814_),
    .B(_08816_),
    .Y(_01332_));
 AOI22x1_ASAP7_75t_R _15958_ (.A1(_00313_),
    .A2(_08806_),
    .B1(_08815_),
    .B2(_08438_),
    .Y(_08817_));
 OA21x2_ASAP7_75t_R _15959_ (.A1(_08733_),
    .A2(_08814_),
    .B(_08817_),
    .Y(_01333_));
 AOI22x1_ASAP7_75t_R _15960_ (.A1(_00280_),
    .A2(_08806_),
    .B1(_08815_),
    .B2(_08459_),
    .Y(_08818_));
 OA21x2_ASAP7_75t_R _15961_ (.A1(_08735_),
    .A2(_08814_),
    .B(_08818_),
    .Y(_01334_));
 AOI22x1_ASAP7_75t_R _15962_ (.A1(_00247_),
    .A2(_08806_),
    .B1(_08815_),
    .B2(_08477_),
    .Y(_08819_));
 OA21x2_ASAP7_75t_R _15963_ (.A1(_08737_),
    .A2(_08814_),
    .B(_08819_),
    .Y(_01335_));
 AOI22x1_ASAP7_75t_R _15964_ (.A1(_00213_),
    .A2(_08806_),
    .B1(_08815_),
    .B2(_08495_),
    .Y(_08820_));
 OA21x2_ASAP7_75t_R _15965_ (.A1(_08739_),
    .A2(_08814_),
    .B(_08820_),
    .Y(_01336_));
 AOI22x1_ASAP7_75t_R _15966_ (.A1(_00180_),
    .A2(_08806_),
    .B1(_08815_),
    .B2(_08512_),
    .Y(_08821_));
 OA21x2_ASAP7_75t_R _15967_ (.A1(_08741_),
    .A2(_08814_),
    .B(_08821_),
    .Y(_01337_));
 OA222x2_ASAP7_75t_R _15968_ (.A1(_04032_),
    .A2(_08791_),
    .B1(_08782_),
    .B2(_08744_),
    .C1(_08792_),
    .C2(_08518_),
    .Y(_01338_));
 AOI22x1_ASAP7_75t_R _15969_ (.A1(_00113_),
    .A2(_08812_),
    .B1(_08815_),
    .B2(_08546_),
    .Y(_08822_));
 OA21x2_ASAP7_75t_R _15970_ (.A1(_08745_),
    .A2(_08814_),
    .B(_08822_),
    .Y(_01339_));
 NOR2x1_ASAP7_75t_R _15971_ (.A(_01011_),
    .B(_08791_),
    .Y(_08823_));
 AO21x1_ASAP7_75t_R _15972_ (.A1(_08747_),
    .A2(_08791_),
    .B(_08823_),
    .Y(_01340_));
 BUFx4f_ASAP7_75t_R _15973_ (.A(_08106_),
    .Y(_08824_));
 AND3x1_ASAP7_75t_R _15974_ (.A(_08824_),
    .B(_08788_),
    .C(_08790_),
    .Y(_08825_));
 NOR2x1_ASAP7_75t_R _15975_ (.A(_00079_),
    .B(_08791_),
    .Y(_08826_));
 AO221x1_ASAP7_75t_R _15976_ (.A1(_08565_),
    .A2(_08791_),
    .B1(_08825_),
    .B2(_08752_),
    .C(_08826_),
    .Y(_01341_));
 AND2x2_ASAP7_75t_R _15977_ (.A(_00047_),
    .B(_08812_),
    .Y(_08827_));
 AOI221x1_ASAP7_75t_R _15978_ (.A1(_08591_),
    .A2(_08825_),
    .B1(_08800_),
    .B2(_08754_),
    .C(_08827_),
    .Y(_01342_));
 AOI22x1_ASAP7_75t_R _15979_ (.A1(_00978_),
    .A2(_08812_),
    .B1(_08815_),
    .B2(_08604_),
    .Y(_08828_));
 OA21x2_ASAP7_75t_R _15980_ (.A1(_08756_),
    .A2(_08814_),
    .B(_08828_),
    .Y(_01343_));
 NAND2x1_ASAP7_75t_R _15981_ (.A(_00945_),
    .B(_08812_),
    .Y(_08829_));
 OA221x2_ASAP7_75t_R _15982_ (.A1(_08758_),
    .A2(_08797_),
    .B1(_08782_),
    .B2(_08619_),
    .C(_08829_),
    .Y(_01344_));
 NAND2x1_ASAP7_75t_R _15983_ (.A(_00911_),
    .B(_08812_),
    .Y(_08830_));
 OA221x2_ASAP7_75t_R _15984_ (.A1(_08631_),
    .A2(_08797_),
    .B1(_08782_),
    .B2(_08760_),
    .C(_08830_),
    .Y(_01345_));
 AOI22x1_ASAP7_75t_R _15985_ (.A1(_00878_),
    .A2(_08812_),
    .B1(_08815_),
    .B2(_08644_),
    .Y(_08831_));
 OA21x2_ASAP7_75t_R _15986_ (.A1(_08762_),
    .A2(_08814_),
    .B(_08831_),
    .Y(_01346_));
 NAND2x1_ASAP7_75t_R _15987_ (.A(_00844_),
    .B(_08796_),
    .Y(_08832_));
 OA21x2_ASAP7_75t_R _15988_ (.A1(_08765_),
    .A2(_08812_),
    .B(_08832_),
    .Y(_08833_));
 OA21x2_ASAP7_75t_R _15989_ (.A1(_08764_),
    .A2(_08814_),
    .B(_08833_),
    .Y(_01347_));
 AOI22x1_ASAP7_75t_R _15990_ (.A1(_00811_),
    .A2(_08812_),
    .B1(_08815_),
    .B2(_08670_),
    .Y(_08834_));
 OA21x2_ASAP7_75t_R _15991_ (.A1(_08768_),
    .A2(_08782_),
    .B(_08834_),
    .Y(_01348_));
 NAND2x1_ASAP7_75t_R _15992_ (.A(_00777_),
    .B(_08796_),
    .Y(_08835_));
 OA21x2_ASAP7_75t_R _15993_ (.A1(_08771_),
    .A2(_08812_),
    .B(_08835_),
    .Y(_08836_));
 OA21x2_ASAP7_75t_R _15994_ (.A1(_08770_),
    .A2(_08782_),
    .B(_08836_),
    .Y(_01349_));
 AND3x4_ASAP7_75t_R _15995_ (.A(_03279_),
    .B(_08774_),
    .C(_08096_),
    .Y(_08837_));
 BUFx16f_ASAP7_75t_R _15996_ (.A(_08837_),
    .Y(_08838_));
 AND2x6_ASAP7_75t_R _15997_ (.A(_08789_),
    .B(_08838_),
    .Y(_08839_));
 NAND2x2_ASAP7_75t_R _15998_ (.A(_08687_),
    .B(_08839_),
    .Y(_08840_));
 BUFx4f_ASAP7_75t_R _15999_ (.A(_08840_),
    .Y(_08841_));
 NAND2x2_ASAP7_75t_R _16000_ (.A(_08115_),
    .B(_08839_),
    .Y(_08842_));
 NAND2x2_ASAP7_75t_R _16001_ (.A(_08789_),
    .B(_08838_),
    .Y(_08843_));
 NAND2x1_ASAP7_75t_R _16002_ (.A(_00013_),
    .B(_08843_),
    .Y(_08844_));
 OA21x2_ASAP7_75t_R _16003_ (.A1(_08111_),
    .A2(_08842_),
    .B(_08844_),
    .Y(_08845_));
 OA21x2_ASAP7_75t_R _16004_ (.A1(_08093_),
    .A2(_08841_),
    .B(_08845_),
    .Y(_01350_));
 BUFx10_ASAP7_75t_R _16005_ (.A(_08843_),
    .Y(_08846_));
 BUFx12_ASAP7_75t_R _16006_ (.A(_08837_),
    .Y(_08847_));
 AND3x2_ASAP7_75t_R _16007_ (.A(_08798_),
    .B(_08790_),
    .C(_08847_),
    .Y(_08848_));
 BUFx10_ASAP7_75t_R _16008_ (.A(_08848_),
    .Y(_08849_));
 AOI22x1_ASAP7_75t_R _16009_ (.A1(_00745_),
    .A2(_08846_),
    .B1(_08849_),
    .B2(_08156_),
    .Y(_08850_));
 OA21x2_ASAP7_75t_R _16010_ (.A1(_08699_),
    .A2(_08841_),
    .B(_08850_),
    .Y(_01351_));
 AOI22x1_ASAP7_75t_R _16011_ (.A1(_00712_),
    .A2(_08846_),
    .B1(_08849_),
    .B2(_08185_),
    .Y(_08851_));
 OA21x2_ASAP7_75t_R _16012_ (.A1(_08705_),
    .A2(_08841_),
    .B(_08851_),
    .Y(_01352_));
 OA222x2_ASAP7_75t_R _16013_ (.A1(_05731_),
    .A2(_08839_),
    .B1(_08840_),
    .B2(_08707_),
    .C1(_08842_),
    .C2(_08191_),
    .Y(_01353_));
 OA222x2_ASAP7_75t_R _16014_ (.A1(_05655_),
    .A2(_08839_),
    .B1(_08840_),
    .B2(_08709_),
    .C1(_08842_),
    .C2(_08211_),
    .Y(_01354_));
 AOI22x1_ASAP7_75t_R _16015_ (.A1(_00613_),
    .A2(_08846_),
    .B1(_08849_),
    .B2(_08243_),
    .Y(_08852_));
 OA21x2_ASAP7_75t_R _16016_ (.A1(_08710_),
    .A2(_08841_),
    .B(_08852_),
    .Y(_01355_));
 AOI22x1_ASAP7_75t_R _16017_ (.A1(_00579_),
    .A2(_08846_),
    .B1(_08849_),
    .B2(_08259_),
    .Y(_08853_));
 OA21x2_ASAP7_75t_R _16018_ (.A1(_08712_),
    .A2(_08841_),
    .B(_08853_),
    .Y(_01356_));
 AOI22x1_ASAP7_75t_R _16019_ (.A1(_00546_),
    .A2(_08846_),
    .B1(_08849_),
    .B2(_08287_),
    .Y(_08854_));
 OA21x2_ASAP7_75t_R _16020_ (.A1(_08714_),
    .A2(_08841_),
    .B(_08854_),
    .Y(_01357_));
 BUFx12_ASAP7_75t_R _16021_ (.A(_08843_),
    .Y(_08855_));
 AOI22x1_ASAP7_75t_R _16022_ (.A1(_00513_),
    .A2(_08855_),
    .B1(_08849_),
    .B2(_08308_),
    .Y(_08856_));
 OA21x2_ASAP7_75t_R _16023_ (.A1(_08716_),
    .A2(_08841_),
    .B(_08856_),
    .Y(_01358_));
 AOI22x1_ASAP7_75t_R _16024_ (.A1(_00480_),
    .A2(_08855_),
    .B1(_08849_),
    .B2(_08327_),
    .Y(_08857_));
 OA21x2_ASAP7_75t_R _16025_ (.A1(_08719_),
    .A2(_08841_),
    .B(_08857_),
    .Y(_01359_));
 AOI22x1_ASAP7_75t_R _16026_ (.A1(_00447_),
    .A2(_08855_),
    .B1(_08849_),
    .B2(_08348_),
    .Y(_08858_));
 OA21x2_ASAP7_75t_R _16027_ (.A1(_08721_),
    .A2(_08841_),
    .B(_08858_),
    .Y(_01360_));
 NAND2x1_ASAP7_75t_R _16028_ (.A(_01045_),
    .B(_08846_),
    .Y(_08859_));
 OA21x2_ASAP7_75t_R _16029_ (.A1(_08723_),
    .A2(_08846_),
    .B(_08859_),
    .Y(_01361_));
 AOI22x1_ASAP7_75t_R _16030_ (.A1(_00414_),
    .A2(_08855_),
    .B1(_08849_),
    .B2(_08382_),
    .Y(_08860_));
 OA21x2_ASAP7_75t_R _16031_ (.A1(_08725_),
    .A2(_08841_),
    .B(_08860_),
    .Y(_01362_));
 BUFx6f_ASAP7_75t_R _16032_ (.A(_08843_),
    .Y(_08861_));
 NAND2x1_ASAP7_75t_R _16033_ (.A(_00381_),
    .B(_08861_),
    .Y(_08862_));
 OA221x2_ASAP7_75t_R _16034_ (.A1(_08401_),
    .A2(_08846_),
    .B1(_08840_),
    .B2(_08727_),
    .C(_08862_),
    .Y(_01363_));
 BUFx4f_ASAP7_75t_R _16035_ (.A(_08840_),
    .Y(_08863_));
 BUFx6f_ASAP7_75t_R _16036_ (.A(_08848_),
    .Y(_08864_));
 AOI22x1_ASAP7_75t_R _16037_ (.A1(_00348_),
    .A2(_08855_),
    .B1(_08864_),
    .B2(_08420_),
    .Y(_08865_));
 OA21x2_ASAP7_75t_R _16038_ (.A1(_08729_),
    .A2(_08863_),
    .B(_08865_),
    .Y(_01364_));
 AOI22x1_ASAP7_75t_R _16039_ (.A1(_00314_),
    .A2(_08855_),
    .B1(_08864_),
    .B2(_08438_),
    .Y(_08866_));
 OA21x2_ASAP7_75t_R _16040_ (.A1(_08733_),
    .A2(_08863_),
    .B(_08866_),
    .Y(_01365_));
 AOI22x1_ASAP7_75t_R _16041_ (.A1(_00281_),
    .A2(_08855_),
    .B1(_08864_),
    .B2(_08459_),
    .Y(_08867_));
 OA21x2_ASAP7_75t_R _16042_ (.A1(_08735_),
    .A2(_08863_),
    .B(_08867_),
    .Y(_01366_));
 AOI22x1_ASAP7_75t_R _16043_ (.A1(_00248_),
    .A2(_08855_),
    .B1(_08864_),
    .B2(_08477_),
    .Y(_08868_));
 OA21x2_ASAP7_75t_R _16044_ (.A1(_08737_),
    .A2(_08863_),
    .B(_08868_),
    .Y(_01367_));
 AOI22x1_ASAP7_75t_R _16045_ (.A1(_00214_),
    .A2(_08855_),
    .B1(_08864_),
    .B2(_08495_),
    .Y(_08869_));
 OA21x2_ASAP7_75t_R _16046_ (.A1(_08739_),
    .A2(_08863_),
    .B(_08869_),
    .Y(_01368_));
 AOI22x1_ASAP7_75t_R _16047_ (.A1(_00181_),
    .A2(_08855_),
    .B1(_08864_),
    .B2(_08512_),
    .Y(_08870_));
 OA21x2_ASAP7_75t_R _16048_ (.A1(_08741_),
    .A2(_08863_),
    .B(_08870_),
    .Y(_01369_));
 OA222x2_ASAP7_75t_R _16049_ (.A1(_04031_),
    .A2(_08839_),
    .B1(_08840_),
    .B2(_08744_),
    .C1(_08842_),
    .C2(_08518_),
    .Y(_01370_));
 AOI22x1_ASAP7_75t_R _16050_ (.A1(_00114_),
    .A2(_08861_),
    .B1(_08864_),
    .B2(_08546_),
    .Y(_08871_));
 OA21x2_ASAP7_75t_R _16051_ (.A1(_08745_),
    .A2(_08863_),
    .B(_08871_),
    .Y(_01371_));
 NOR2x1_ASAP7_75t_R _16052_ (.A(_01012_),
    .B(_08839_),
    .Y(_08872_));
 AO21x1_ASAP7_75t_R _16053_ (.A1(_08747_),
    .A2(_08839_),
    .B(_08872_),
    .Y(_01372_));
 BUFx10_ASAP7_75t_R _16054_ (.A(_08838_),
    .Y(_08873_));
 AND3x1_ASAP7_75t_R _16055_ (.A(_08824_),
    .B(_08790_),
    .C(_08873_),
    .Y(_08874_));
 NOR2x1_ASAP7_75t_R _16056_ (.A(_00080_),
    .B(_08839_),
    .Y(_08875_));
 AO221x1_ASAP7_75t_R _16057_ (.A1(_08565_),
    .A2(_08839_),
    .B1(_08874_),
    .B2(_08752_),
    .C(_08875_),
    .Y(_01373_));
 AND2x2_ASAP7_75t_R _16058_ (.A(_00048_),
    .B(_08861_),
    .Y(_08876_));
 AOI221x1_ASAP7_75t_R _16059_ (.A1(_08591_),
    .A2(_08874_),
    .B1(_08849_),
    .B2(_08754_),
    .C(_08876_),
    .Y(_01374_));
 AOI22x1_ASAP7_75t_R _16060_ (.A1(_00979_),
    .A2(_08861_),
    .B1(_08864_),
    .B2(_08604_),
    .Y(_08877_));
 OA21x2_ASAP7_75t_R _16061_ (.A1(_08756_),
    .A2(_08863_),
    .B(_08877_),
    .Y(_01375_));
 NAND2x1_ASAP7_75t_R _16062_ (.A(_00946_),
    .B(_08861_),
    .Y(_08878_));
 OA221x2_ASAP7_75t_R _16063_ (.A1(_08758_),
    .A2(_08846_),
    .B1(_08840_),
    .B2(_08619_),
    .C(_08878_),
    .Y(_01376_));
 NAND2x1_ASAP7_75t_R _16064_ (.A(_00912_),
    .B(_08861_),
    .Y(_08879_));
 OA221x2_ASAP7_75t_R _16065_ (.A1(_08631_),
    .A2(_08846_),
    .B1(_08840_),
    .B2(_08760_),
    .C(_08879_),
    .Y(_01377_));
 AOI22x1_ASAP7_75t_R _16066_ (.A1(_00879_),
    .A2(_08861_),
    .B1(_08864_),
    .B2(_08644_),
    .Y(_08880_));
 OA21x2_ASAP7_75t_R _16067_ (.A1(_08762_),
    .A2(_08863_),
    .B(_08880_),
    .Y(_01378_));
 NAND2x1_ASAP7_75t_R _16068_ (.A(_00845_),
    .B(_08843_),
    .Y(_08881_));
 OA21x2_ASAP7_75t_R _16069_ (.A1(_08765_),
    .A2(_08861_),
    .B(_08881_),
    .Y(_08882_));
 OA21x2_ASAP7_75t_R _16070_ (.A1(_08764_),
    .A2(_08863_),
    .B(_08882_),
    .Y(_01379_));
 AOI22x1_ASAP7_75t_R _16071_ (.A1(_00812_),
    .A2(_08861_),
    .B1(_08864_),
    .B2(_08670_),
    .Y(_08883_));
 OA21x2_ASAP7_75t_R _16072_ (.A1(_08768_),
    .A2(_08840_),
    .B(_08883_),
    .Y(_01380_));
 NAND2x1_ASAP7_75t_R _16073_ (.A(_00778_),
    .B(_08843_),
    .Y(_08884_));
 OA21x2_ASAP7_75t_R _16074_ (.A1(_08771_),
    .A2(_08861_),
    .B(_08884_),
    .Y(_08885_));
 OA21x2_ASAP7_75t_R _16075_ (.A1(_08770_),
    .A2(_08840_),
    .B(_08885_),
    .Y(_01381_));
 AND2x6_ASAP7_75t_R _16076_ (.A(_08098_),
    .B(_08789_),
    .Y(_08886_));
 NAND2x2_ASAP7_75t_R _16077_ (.A(_08687_),
    .B(_08886_),
    .Y(_08887_));
 BUFx4f_ASAP7_75t_R _16078_ (.A(_08887_),
    .Y(_08888_));
 NAND2x2_ASAP7_75t_R _16079_ (.A(_08115_),
    .B(_08886_),
    .Y(_08889_));
 NAND2x2_ASAP7_75t_R _16080_ (.A(_08117_),
    .B(_08789_),
    .Y(_08890_));
 NAND2x1_ASAP7_75t_R _16081_ (.A(_00014_),
    .B(_08890_),
    .Y(_08891_));
 OA21x2_ASAP7_75t_R _16082_ (.A1(_08111_),
    .A2(_08889_),
    .B(_08891_),
    .Y(_08892_));
 OA21x2_ASAP7_75t_R _16083_ (.A1(_08093_),
    .A2(_08888_),
    .B(_08892_),
    .Y(_01382_));
 BUFx10_ASAP7_75t_R _16084_ (.A(_08890_),
    .Y(_08893_));
 AND3x2_ASAP7_75t_R _16085_ (.A(_08145_),
    .B(_08701_),
    .C(_08790_),
    .Y(_08894_));
 BUFx10_ASAP7_75t_R _16086_ (.A(_08894_),
    .Y(_08895_));
 AOI22x1_ASAP7_75t_R _16087_ (.A1(_00746_),
    .A2(_08893_),
    .B1(_08895_),
    .B2(_08156_),
    .Y(_08896_));
 OA21x2_ASAP7_75t_R _16088_ (.A1(_08699_),
    .A2(_08888_),
    .B(_08896_),
    .Y(_01383_));
 AOI22x1_ASAP7_75t_R _16089_ (.A1(_00713_),
    .A2(_08893_),
    .B1(_08895_),
    .B2(_08185_),
    .Y(_08897_));
 OA21x2_ASAP7_75t_R _16090_ (.A1(_08705_),
    .A2(_08888_),
    .B(_08897_),
    .Y(_01384_));
 INVx1_ASAP7_75t_R _16091_ (.A(_00680_),
    .Y(_08898_));
 OA222x2_ASAP7_75t_R _16092_ (.A1(_08898_),
    .A2(_08886_),
    .B1(_08887_),
    .B2(_08707_),
    .C1(_08889_),
    .C2(_08191_),
    .Y(_01385_));
 INVx1_ASAP7_75t_R _16093_ (.A(_00647_),
    .Y(_08899_));
 OA222x2_ASAP7_75t_R _16094_ (.A1(_08899_),
    .A2(_08886_),
    .B1(_08887_),
    .B2(_08709_),
    .C1(_08889_),
    .C2(_08211_),
    .Y(_01386_));
 AOI22x1_ASAP7_75t_R _16095_ (.A1(_00614_),
    .A2(_08893_),
    .B1(_08895_),
    .B2(_08243_),
    .Y(_08900_));
 OA21x2_ASAP7_75t_R _16096_ (.A1(_08710_),
    .A2(_08888_),
    .B(_08900_),
    .Y(_01387_));
 AOI22x1_ASAP7_75t_R _16097_ (.A1(_00580_),
    .A2(_08893_),
    .B1(_08895_),
    .B2(_08259_),
    .Y(_08901_));
 OA21x2_ASAP7_75t_R _16098_ (.A1(_08712_),
    .A2(_08888_),
    .B(_08901_),
    .Y(_01388_));
 AOI22x1_ASAP7_75t_R _16099_ (.A1(_00547_),
    .A2(_08893_),
    .B1(_08895_),
    .B2(_08287_),
    .Y(_08902_));
 OA21x2_ASAP7_75t_R _16100_ (.A1(_08714_),
    .A2(_08888_),
    .B(_08902_),
    .Y(_01389_));
 BUFx12_ASAP7_75t_R _16101_ (.A(_08890_),
    .Y(_08903_));
 AOI22x1_ASAP7_75t_R _16102_ (.A1(_00514_),
    .A2(_08903_),
    .B1(_08895_),
    .B2(_08308_),
    .Y(_08904_));
 OA21x2_ASAP7_75t_R _16103_ (.A1(_08716_),
    .A2(_08888_),
    .B(_08904_),
    .Y(_01390_));
 AOI22x1_ASAP7_75t_R _16104_ (.A1(_00481_),
    .A2(_08903_),
    .B1(_08895_),
    .B2(_08327_),
    .Y(_08905_));
 OA21x2_ASAP7_75t_R _16105_ (.A1(_08719_),
    .A2(_08888_),
    .B(_08905_),
    .Y(_01391_));
 AOI22x1_ASAP7_75t_R _16106_ (.A1(_00448_),
    .A2(_08903_),
    .B1(_08895_),
    .B2(_08348_),
    .Y(_08906_));
 OA21x2_ASAP7_75t_R _16107_ (.A1(_08721_),
    .A2(_08888_),
    .B(_08906_),
    .Y(_01392_));
 NAND2x1_ASAP7_75t_R _16108_ (.A(_01046_),
    .B(_08893_),
    .Y(_08907_));
 OA21x2_ASAP7_75t_R _16109_ (.A1(_08723_),
    .A2(_08893_),
    .B(_08907_),
    .Y(_01393_));
 AOI22x1_ASAP7_75t_R _16110_ (.A1(_00415_),
    .A2(_08903_),
    .B1(_08895_),
    .B2(_08382_),
    .Y(_08908_));
 OA21x2_ASAP7_75t_R _16111_ (.A1(_08725_),
    .A2(_08888_),
    .B(_08908_),
    .Y(_01394_));
 BUFx6f_ASAP7_75t_R _16112_ (.A(_08890_),
    .Y(_08909_));
 NAND2x1_ASAP7_75t_R _16113_ (.A(_00382_),
    .B(_08909_),
    .Y(_08910_));
 OA221x2_ASAP7_75t_R _16114_ (.A1(_08401_),
    .A2(_08893_),
    .B1(_08887_),
    .B2(_08727_),
    .C(_08910_),
    .Y(_01395_));
 BUFx4f_ASAP7_75t_R _16115_ (.A(_08887_),
    .Y(_08911_));
 BUFx6f_ASAP7_75t_R _16116_ (.A(_08894_),
    .Y(_08912_));
 AOI22x1_ASAP7_75t_R _16117_ (.A1(_00349_),
    .A2(_08903_),
    .B1(_08912_),
    .B2(_08420_),
    .Y(_08913_));
 OA21x2_ASAP7_75t_R _16118_ (.A1(_08729_),
    .A2(_08911_),
    .B(_08913_),
    .Y(_01396_));
 AOI22x1_ASAP7_75t_R _16119_ (.A1(_00315_),
    .A2(_08903_),
    .B1(_08912_),
    .B2(_08438_),
    .Y(_08914_));
 OA21x2_ASAP7_75t_R _16120_ (.A1(_08733_),
    .A2(_08911_),
    .B(_08914_),
    .Y(_01397_));
 AOI22x1_ASAP7_75t_R _16121_ (.A1(_00282_),
    .A2(_08903_),
    .B1(_08912_),
    .B2(_08459_),
    .Y(_08915_));
 OA21x2_ASAP7_75t_R _16122_ (.A1(_08735_),
    .A2(_08911_),
    .B(_08915_),
    .Y(_01398_));
 AOI22x1_ASAP7_75t_R _16123_ (.A1(_00249_),
    .A2(_08903_),
    .B1(_08912_),
    .B2(_08477_),
    .Y(_08916_));
 OA21x2_ASAP7_75t_R _16124_ (.A1(_08737_),
    .A2(_08911_),
    .B(_08916_),
    .Y(_01399_));
 AOI22x1_ASAP7_75t_R _16125_ (.A1(_00215_),
    .A2(_08903_),
    .B1(_08912_),
    .B2(_08495_),
    .Y(_08917_));
 OA21x2_ASAP7_75t_R _16126_ (.A1(_08739_),
    .A2(_08911_),
    .B(_08917_),
    .Y(_01400_));
 AOI22x1_ASAP7_75t_R _16127_ (.A1(_00182_),
    .A2(_08903_),
    .B1(_08912_),
    .B2(_08512_),
    .Y(_08918_));
 OA21x2_ASAP7_75t_R _16128_ (.A1(_08741_),
    .A2(_08911_),
    .B(_08918_),
    .Y(_01401_));
 INVx1_ASAP7_75t_R _16129_ (.A(_00148_),
    .Y(_08919_));
 OA222x2_ASAP7_75t_R _16130_ (.A1(_08919_),
    .A2(_08886_),
    .B1(_08887_),
    .B2(_08744_),
    .C1(_08889_),
    .C2(_08518_),
    .Y(_01402_));
 AOI22x1_ASAP7_75t_R _16131_ (.A1(_00115_),
    .A2(_08909_),
    .B1(_08912_),
    .B2(_08546_),
    .Y(_08920_));
 OA21x2_ASAP7_75t_R _16132_ (.A1(_08745_),
    .A2(_08911_),
    .B(_08920_),
    .Y(_01403_));
 NOR2x1_ASAP7_75t_R _16133_ (.A(_01013_),
    .B(_08886_),
    .Y(_08921_));
 AO21x1_ASAP7_75t_R _16134_ (.A1(_08747_),
    .A2(_08886_),
    .B(_08921_),
    .Y(_01404_));
 AND3x1_ASAP7_75t_R _16135_ (.A(_08145_),
    .B(_08577_),
    .C(_08790_),
    .Y(_08922_));
 NOR2x1_ASAP7_75t_R _16136_ (.A(_00081_),
    .B(_08886_),
    .Y(_08923_));
 AO221x1_ASAP7_75t_R _16137_ (.A1(_08565_),
    .A2(_08886_),
    .B1(_08922_),
    .B2(_08752_),
    .C(_08923_),
    .Y(_01405_));
 AND2x2_ASAP7_75t_R _16138_ (.A(_00049_),
    .B(_08909_),
    .Y(_08924_));
 AOI221x1_ASAP7_75t_R _16139_ (.A1(_08591_),
    .A2(_08922_),
    .B1(_08895_),
    .B2(_08754_),
    .C(_08924_),
    .Y(_01406_));
 AOI22x1_ASAP7_75t_R _16140_ (.A1(_00980_),
    .A2(_08909_),
    .B1(_08912_),
    .B2(_08604_),
    .Y(_08925_));
 OA21x2_ASAP7_75t_R _16141_ (.A1(_08756_),
    .A2(_08911_),
    .B(_08925_),
    .Y(_01407_));
 NAND2x1_ASAP7_75t_R _16142_ (.A(_00947_),
    .B(_08909_),
    .Y(_08926_));
 OA221x2_ASAP7_75t_R _16143_ (.A1(_08758_),
    .A2(_08893_),
    .B1(_08887_),
    .B2(_08619_),
    .C(_08926_),
    .Y(_01408_));
 NAND2x1_ASAP7_75t_R _16144_ (.A(_00913_),
    .B(_08909_),
    .Y(_08927_));
 OA221x2_ASAP7_75t_R _16145_ (.A1(_08631_),
    .A2(_08893_),
    .B1(_08887_),
    .B2(_08760_),
    .C(_08927_),
    .Y(_01409_));
 AOI22x1_ASAP7_75t_R _16146_ (.A1(_00880_),
    .A2(_08909_),
    .B1(_08912_),
    .B2(_08644_),
    .Y(_08928_));
 OA21x2_ASAP7_75t_R _16147_ (.A1(_08762_),
    .A2(_08911_),
    .B(_08928_),
    .Y(_01410_));
 NAND2x1_ASAP7_75t_R _16148_ (.A(_00846_),
    .B(_08890_),
    .Y(_08929_));
 OA21x2_ASAP7_75t_R _16149_ (.A1(_08765_),
    .A2(_08909_),
    .B(_08929_),
    .Y(_08930_));
 OA21x2_ASAP7_75t_R _16150_ (.A1(_08764_),
    .A2(_08911_),
    .B(_08930_),
    .Y(_01411_));
 AOI22x1_ASAP7_75t_R _16151_ (.A1(_00813_),
    .A2(_08909_),
    .B1(_08912_),
    .B2(_08670_),
    .Y(_08931_));
 OA21x2_ASAP7_75t_R _16152_ (.A1(_08768_),
    .A2(_08887_),
    .B(_08931_),
    .Y(_01412_));
 NAND2x1_ASAP7_75t_R _16153_ (.A(_00779_),
    .B(_08890_),
    .Y(_08932_));
 OA21x2_ASAP7_75t_R _16154_ (.A1(_08771_),
    .A2(_08909_),
    .B(_08932_),
    .Y(_08933_));
 OA21x2_ASAP7_75t_R _16155_ (.A1(_08770_),
    .A2(_08887_),
    .B(_08933_),
    .Y(_01413_));
 AND2x6_ASAP7_75t_R _16156_ (.A(_08689_),
    .B(_08789_),
    .Y(_08934_));
 NAND2x2_ASAP7_75t_R _16157_ (.A(_08687_),
    .B(_08934_),
    .Y(_08935_));
 BUFx4f_ASAP7_75t_R _16158_ (.A(_08935_),
    .Y(_08936_));
 BUFx16f_ASAP7_75t_R _16159_ (.A(_08798_),
    .Y(_08937_));
 NAND2x2_ASAP7_75t_R _16160_ (.A(_08937_),
    .B(_08934_),
    .Y(_08938_));
 OA22x2_ASAP7_75t_R _16161_ (.A1(_03150_),
    .A2(_08934_),
    .B1(_08938_),
    .B2(_08793_),
    .Y(_08939_));
 OA21x2_ASAP7_75t_R _16162_ (.A1(_08093_),
    .A2(_08936_),
    .B(_08939_),
    .Y(_01414_));
 NAND2x2_ASAP7_75t_R _16163_ (.A(_08694_),
    .B(_08789_),
    .Y(_08940_));
 BUFx10_ASAP7_75t_R _16164_ (.A(_08940_),
    .Y(_08941_));
 AND3x2_ASAP7_75t_R _16165_ (.A(_08798_),
    .B(_08749_),
    .C(_08790_),
    .Y(_08942_));
 BUFx10_ASAP7_75t_R _16166_ (.A(_08942_),
    .Y(_08943_));
 AOI22x1_ASAP7_75t_R _16167_ (.A1(_00747_),
    .A2(_08941_),
    .B1(_08943_),
    .B2(_08156_),
    .Y(_08944_));
 OA21x2_ASAP7_75t_R _16168_ (.A1(_08699_),
    .A2(_08936_),
    .B(_08944_),
    .Y(_01415_));
 AOI22x1_ASAP7_75t_R _16169_ (.A1(_00714_),
    .A2(_08941_),
    .B1(_08943_),
    .B2(_08185_),
    .Y(_08945_));
 OA21x2_ASAP7_75t_R _16170_ (.A1(_08705_),
    .A2(_08936_),
    .B(_08945_),
    .Y(_01416_));
 INVx1_ASAP7_75t_R _16171_ (.A(_00681_),
    .Y(_08946_));
 OA222x2_ASAP7_75t_R _16172_ (.A1(_08946_),
    .A2(_08934_),
    .B1(_08935_),
    .B2(_08707_),
    .C1(_08938_),
    .C2(_08191_),
    .Y(_01417_));
 INVx1_ASAP7_75t_R _16173_ (.A(_00648_),
    .Y(_08947_));
 OA222x2_ASAP7_75t_R _16174_ (.A1(_08947_),
    .A2(_08934_),
    .B1(_08935_),
    .B2(_08709_),
    .C1(_08938_),
    .C2(_08211_),
    .Y(_01418_));
 AOI22x1_ASAP7_75t_R _16175_ (.A1(_00615_),
    .A2(_08941_),
    .B1(_08943_),
    .B2(_08243_),
    .Y(_08948_));
 OA21x2_ASAP7_75t_R _16176_ (.A1(_08710_),
    .A2(_08936_),
    .B(_08948_),
    .Y(_01419_));
 AOI22x1_ASAP7_75t_R _16177_ (.A1(_00581_),
    .A2(_08941_),
    .B1(_08943_),
    .B2(_08259_),
    .Y(_08949_));
 OA21x2_ASAP7_75t_R _16178_ (.A1(_08712_),
    .A2(_08936_),
    .B(_08949_),
    .Y(_01420_));
 AOI22x1_ASAP7_75t_R _16179_ (.A1(_00548_),
    .A2(_08941_),
    .B1(_08943_),
    .B2(_08287_),
    .Y(_08950_));
 OA21x2_ASAP7_75t_R _16180_ (.A1(_08714_),
    .A2(_08936_),
    .B(_08950_),
    .Y(_01421_));
 BUFx12_ASAP7_75t_R _16181_ (.A(_08940_),
    .Y(_08951_));
 AOI22x1_ASAP7_75t_R _16182_ (.A1(_00515_),
    .A2(_08951_),
    .B1(_08943_),
    .B2(_08308_),
    .Y(_08952_));
 OA21x2_ASAP7_75t_R _16183_ (.A1(_08716_),
    .A2(_08936_),
    .B(_08952_),
    .Y(_01422_));
 AOI22x1_ASAP7_75t_R _16184_ (.A1(_00482_),
    .A2(_08951_),
    .B1(_08943_),
    .B2(_08327_),
    .Y(_08953_));
 OA21x2_ASAP7_75t_R _16185_ (.A1(_08719_),
    .A2(_08936_),
    .B(_08953_),
    .Y(_01423_));
 AOI22x1_ASAP7_75t_R _16186_ (.A1(_00449_),
    .A2(_08951_),
    .B1(_08943_),
    .B2(_08348_),
    .Y(_08954_));
 OA21x2_ASAP7_75t_R _16187_ (.A1(_08721_),
    .A2(_08936_),
    .B(_08954_),
    .Y(_01424_));
 NAND2x1_ASAP7_75t_R _16188_ (.A(_01047_),
    .B(_08941_),
    .Y(_08955_));
 OA21x2_ASAP7_75t_R _16189_ (.A1(_08723_),
    .A2(_08941_),
    .B(_08955_),
    .Y(_01425_));
 AOI22x1_ASAP7_75t_R _16190_ (.A1(_00416_),
    .A2(_08951_),
    .B1(_08943_),
    .B2(_08382_),
    .Y(_08956_));
 OA21x2_ASAP7_75t_R _16191_ (.A1(_08725_),
    .A2(_08936_),
    .B(_08956_),
    .Y(_01426_));
 BUFx6f_ASAP7_75t_R _16192_ (.A(_08940_),
    .Y(_08957_));
 NAND2x1_ASAP7_75t_R _16193_ (.A(_00383_),
    .B(_08957_),
    .Y(_08958_));
 OA221x2_ASAP7_75t_R _16194_ (.A1(_08401_),
    .A2(_08941_),
    .B1(_08935_),
    .B2(_08727_),
    .C(_08958_),
    .Y(_01427_));
 BUFx4f_ASAP7_75t_R _16195_ (.A(_08935_),
    .Y(_08959_));
 BUFx10_ASAP7_75t_R _16196_ (.A(_08942_),
    .Y(_08960_));
 AOI22x1_ASAP7_75t_R _16197_ (.A1(_00350_),
    .A2(_08951_),
    .B1(_08960_),
    .B2(_08420_),
    .Y(_08961_));
 OA21x2_ASAP7_75t_R _16198_ (.A1(_08729_),
    .A2(_08959_),
    .B(_08961_),
    .Y(_01428_));
 AOI22x1_ASAP7_75t_R _16199_ (.A1(_00316_),
    .A2(_08951_),
    .B1(_08960_),
    .B2(_08438_),
    .Y(_08962_));
 OA21x2_ASAP7_75t_R _16200_ (.A1(_08733_),
    .A2(_08959_),
    .B(_08962_),
    .Y(_01429_));
 AOI22x1_ASAP7_75t_R _16201_ (.A1(_00283_),
    .A2(_08951_),
    .B1(_08960_),
    .B2(_08459_),
    .Y(_08963_));
 OA21x2_ASAP7_75t_R _16202_ (.A1(_08735_),
    .A2(_08959_),
    .B(_08963_),
    .Y(_01430_));
 AOI22x1_ASAP7_75t_R _16203_ (.A1(_00250_),
    .A2(_08951_),
    .B1(_08960_),
    .B2(_08477_),
    .Y(_08964_));
 OA21x2_ASAP7_75t_R _16204_ (.A1(_08737_),
    .A2(_08959_),
    .B(_08964_),
    .Y(_01431_));
 AOI22x1_ASAP7_75t_R _16205_ (.A1(_00216_),
    .A2(_08951_),
    .B1(_08960_),
    .B2(_08495_),
    .Y(_08965_));
 OA21x2_ASAP7_75t_R _16206_ (.A1(_08739_),
    .A2(_08959_),
    .B(_08965_),
    .Y(_01432_));
 AOI22x1_ASAP7_75t_R _16207_ (.A1(_00183_),
    .A2(_08951_),
    .B1(_08960_),
    .B2(_08512_),
    .Y(_08966_));
 OA21x2_ASAP7_75t_R _16208_ (.A1(_08741_),
    .A2(_08959_),
    .B(_08966_),
    .Y(_01433_));
 INVx1_ASAP7_75t_R _16209_ (.A(_00149_),
    .Y(_08967_));
 OA222x2_ASAP7_75t_R _16210_ (.A1(_08967_),
    .A2(_08934_),
    .B1(_08935_),
    .B2(_08744_),
    .C1(_08938_),
    .C2(_08518_),
    .Y(_01434_));
 AOI22x1_ASAP7_75t_R _16211_ (.A1(_00116_),
    .A2(_08957_),
    .B1(_08960_),
    .B2(_08546_),
    .Y(_08968_));
 OA21x2_ASAP7_75t_R _16212_ (.A1(_08745_),
    .A2(_08959_),
    .B(_08968_),
    .Y(_01435_));
 NOR2x1_ASAP7_75t_R _16213_ (.A(_01014_),
    .B(_08934_),
    .Y(_08969_));
 AO21x1_ASAP7_75t_R _16214_ (.A1(_08747_),
    .A2(_08934_),
    .B(_08969_),
    .Y(_01436_));
 AND3x1_ASAP7_75t_R _16215_ (.A(_08824_),
    .B(_08750_),
    .C(_08790_),
    .Y(_08970_));
 NOR2x1_ASAP7_75t_R _16216_ (.A(_00082_),
    .B(_08934_),
    .Y(_08971_));
 AO221x1_ASAP7_75t_R _16217_ (.A1(_08565_),
    .A2(_08934_),
    .B1(_08970_),
    .B2(_08752_),
    .C(_08971_),
    .Y(_01437_));
 AND2x2_ASAP7_75t_R _16218_ (.A(_00050_),
    .B(_08957_),
    .Y(_08972_));
 AOI221x1_ASAP7_75t_R _16219_ (.A1(_08591_),
    .A2(_08970_),
    .B1(_08943_),
    .B2(_08754_),
    .C(_08972_),
    .Y(_01438_));
 AOI22x1_ASAP7_75t_R _16220_ (.A1(_00981_),
    .A2(_08957_),
    .B1(_08960_),
    .B2(_08604_),
    .Y(_08973_));
 OA21x2_ASAP7_75t_R _16221_ (.A1(_08756_),
    .A2(_08959_),
    .B(_08973_),
    .Y(_01439_));
 NAND2x1_ASAP7_75t_R _16222_ (.A(_00948_),
    .B(_08957_),
    .Y(_08974_));
 OA221x2_ASAP7_75t_R _16223_ (.A1(_08758_),
    .A2(_08941_),
    .B1(_08935_),
    .B2(_08619_),
    .C(_08974_),
    .Y(_01440_));
 NAND2x1_ASAP7_75t_R _16224_ (.A(_00914_),
    .B(_08957_),
    .Y(_08975_));
 OA221x2_ASAP7_75t_R _16225_ (.A1(_08631_),
    .A2(_08941_),
    .B1(_08935_),
    .B2(_08760_),
    .C(_08975_),
    .Y(_01441_));
 AOI22x1_ASAP7_75t_R _16226_ (.A1(_00881_),
    .A2(_08957_),
    .B1(_08960_),
    .B2(_08644_),
    .Y(_08976_));
 OA21x2_ASAP7_75t_R _16227_ (.A1(_08762_),
    .A2(_08959_),
    .B(_08976_),
    .Y(_01442_));
 NAND2x1_ASAP7_75t_R _16228_ (.A(_00847_),
    .B(_08940_),
    .Y(_08977_));
 OA21x2_ASAP7_75t_R _16229_ (.A1(_08765_),
    .A2(_08957_),
    .B(_08977_),
    .Y(_08978_));
 OA21x2_ASAP7_75t_R _16230_ (.A1(_08764_),
    .A2(_08959_),
    .B(_08978_),
    .Y(_01443_));
 AOI22x1_ASAP7_75t_R _16231_ (.A1(_00814_),
    .A2(_08957_),
    .B1(_08960_),
    .B2(_08670_),
    .Y(_08979_));
 OA21x2_ASAP7_75t_R _16232_ (.A1(_08768_),
    .A2(_08935_),
    .B(_08979_),
    .Y(_01444_));
 NAND2x1_ASAP7_75t_R _16233_ (.A(_00780_),
    .B(_08940_),
    .Y(_08980_));
 OA21x2_ASAP7_75t_R _16234_ (.A1(_08771_),
    .A2(_08957_),
    .B(_08980_),
    .Y(_08981_));
 OA21x2_ASAP7_75t_R _16235_ (.A1(_08770_),
    .A2(_08935_),
    .B(_08981_),
    .Y(_01445_));
 AND4x1_ASAP7_75t_R _16236_ (.A(_03025_),
    .B(net5),
    .C(_08779_),
    .D(_08100_),
    .Y(_08982_));
 BUFx4f_ASAP7_75t_R _16237_ (.A(_08982_),
    .Y(_08983_));
 AND2x6_ASAP7_75t_R _16238_ (.A(_08787_),
    .B(_08983_),
    .Y(_08984_));
 NAND2x2_ASAP7_75t_R _16239_ (.A(_08687_),
    .B(_08984_),
    .Y(_08985_));
 BUFx4f_ASAP7_75t_R _16240_ (.A(_08985_),
    .Y(_08986_));
 NAND2x2_ASAP7_75t_R _16241_ (.A(_08937_),
    .B(_08984_),
    .Y(_08987_));
 OA22x2_ASAP7_75t_R _16242_ (.A1(_03108_),
    .A2(_08984_),
    .B1(_08987_),
    .B2(_08793_),
    .Y(_08988_));
 OA21x2_ASAP7_75t_R _16243_ (.A1(_08093_),
    .A2(_08986_),
    .B(_08988_),
    .Y(_01446_));
 BUFx6f_ASAP7_75t_R _16244_ (.A(_08983_),
    .Y(_08989_));
 NAND2x2_ASAP7_75t_R _16245_ (.A(_08795_),
    .B(_08989_),
    .Y(_08990_));
 BUFx10_ASAP7_75t_R _16246_ (.A(_08990_),
    .Y(_08991_));
 AND3x2_ASAP7_75t_R _16247_ (.A(_08798_),
    .B(_08795_),
    .C(_08989_),
    .Y(_08992_));
 BUFx10_ASAP7_75t_R _16248_ (.A(_08992_),
    .Y(_08993_));
 AOI22x1_ASAP7_75t_R _16249_ (.A1(_00748_),
    .A2(_08991_),
    .B1(_08993_),
    .B2(_08156_),
    .Y(_08994_));
 OA21x2_ASAP7_75t_R _16250_ (.A1(_08699_),
    .A2(_08986_),
    .B(_08994_),
    .Y(_01447_));
 AOI22x1_ASAP7_75t_R _16251_ (.A1(_00715_),
    .A2(_08991_),
    .B1(_08993_),
    .B2(_08185_),
    .Y(_08995_));
 OA21x2_ASAP7_75t_R _16252_ (.A1(_08705_),
    .A2(_08986_),
    .B(_08995_),
    .Y(_01448_));
 OA222x2_ASAP7_75t_R _16253_ (.A1(_05744_),
    .A2(_08984_),
    .B1(_08985_),
    .B2(_08707_),
    .C1(_08987_),
    .C2(_08191_),
    .Y(_01449_));
 INVx1_ASAP7_75t_R _16254_ (.A(_00649_),
    .Y(_08996_));
 OA222x2_ASAP7_75t_R _16255_ (.A1(_08996_),
    .A2(_08984_),
    .B1(_08985_),
    .B2(_08709_),
    .C1(_08987_),
    .C2(_08211_),
    .Y(_01450_));
 AOI22x1_ASAP7_75t_R _16256_ (.A1(_00616_),
    .A2(_08991_),
    .B1(_08993_),
    .B2(_08243_),
    .Y(_08997_));
 OA21x2_ASAP7_75t_R _16257_ (.A1(_08710_),
    .A2(_08986_),
    .B(_08997_),
    .Y(_01451_));
 AOI22x1_ASAP7_75t_R _16258_ (.A1(_00582_),
    .A2(_08991_),
    .B1(_08993_),
    .B2(_08259_),
    .Y(_08998_));
 OA21x2_ASAP7_75t_R _16259_ (.A1(_08712_),
    .A2(_08986_),
    .B(_08998_),
    .Y(_01452_));
 AOI22x1_ASAP7_75t_R _16260_ (.A1(_00549_),
    .A2(_08991_),
    .B1(_08993_),
    .B2(_08287_),
    .Y(_08999_));
 OA21x2_ASAP7_75t_R _16261_ (.A1(_08714_),
    .A2(_08986_),
    .B(_08999_),
    .Y(_01453_));
 BUFx12_ASAP7_75t_R _16262_ (.A(_08990_),
    .Y(_09000_));
 AOI22x1_ASAP7_75t_R _16263_ (.A1(_00516_),
    .A2(_09000_),
    .B1(_08993_),
    .B2(_08308_),
    .Y(_09001_));
 OA21x2_ASAP7_75t_R _16264_ (.A1(_08716_),
    .A2(_08986_),
    .B(_09001_),
    .Y(_01454_));
 AOI22x1_ASAP7_75t_R _16265_ (.A1(_00483_),
    .A2(_09000_),
    .B1(_08993_),
    .B2(_08327_),
    .Y(_09002_));
 OA21x2_ASAP7_75t_R _16266_ (.A1(_08719_),
    .A2(_08986_),
    .B(_09002_),
    .Y(_01455_));
 AOI22x1_ASAP7_75t_R _16267_ (.A1(_00450_),
    .A2(_09000_),
    .B1(_08993_),
    .B2(_08348_),
    .Y(_09003_));
 OA21x2_ASAP7_75t_R _16268_ (.A1(_08721_),
    .A2(_08986_),
    .B(_09003_),
    .Y(_01456_));
 NAND2x1_ASAP7_75t_R _16269_ (.A(_01048_),
    .B(_08991_),
    .Y(_09004_));
 OA21x2_ASAP7_75t_R _16270_ (.A1(_08723_),
    .A2(_08991_),
    .B(_09004_),
    .Y(_01457_));
 AOI22x1_ASAP7_75t_R _16271_ (.A1(_00417_),
    .A2(_09000_),
    .B1(_08993_),
    .B2(_08382_),
    .Y(_09005_));
 OA21x2_ASAP7_75t_R _16272_ (.A1(_08725_),
    .A2(_08986_),
    .B(_09005_),
    .Y(_01458_));
 BUFx6f_ASAP7_75t_R _16273_ (.A(_08990_),
    .Y(_09006_));
 NAND2x1_ASAP7_75t_R _16274_ (.A(_00384_),
    .B(_09006_),
    .Y(_09007_));
 OA221x2_ASAP7_75t_R _16275_ (.A1(_08401_),
    .A2(_08991_),
    .B1(_08985_),
    .B2(_08727_),
    .C(_09007_),
    .Y(_01459_));
 BUFx4f_ASAP7_75t_R _16276_ (.A(_08985_),
    .Y(_09008_));
 BUFx6f_ASAP7_75t_R _16277_ (.A(_08992_),
    .Y(_09009_));
 AOI22x1_ASAP7_75t_R _16278_ (.A1(_00351_),
    .A2(_09000_),
    .B1(_09009_),
    .B2(_08420_),
    .Y(_09010_));
 OA21x2_ASAP7_75t_R _16279_ (.A1(_08729_),
    .A2(_09008_),
    .B(_09010_),
    .Y(_01460_));
 AOI22x1_ASAP7_75t_R _16280_ (.A1(_00317_),
    .A2(_09000_),
    .B1(_09009_),
    .B2(_08438_),
    .Y(_09011_));
 OA21x2_ASAP7_75t_R _16281_ (.A1(_08733_),
    .A2(_09008_),
    .B(_09011_),
    .Y(_01461_));
 AOI22x1_ASAP7_75t_R _16282_ (.A1(_00284_),
    .A2(_09000_),
    .B1(_09009_),
    .B2(_08459_),
    .Y(_09012_));
 OA21x2_ASAP7_75t_R _16283_ (.A1(_08735_),
    .A2(_09008_),
    .B(_09012_),
    .Y(_01462_));
 AOI22x1_ASAP7_75t_R _16284_ (.A1(_00251_),
    .A2(_09000_),
    .B1(_09009_),
    .B2(_08477_),
    .Y(_09013_));
 OA21x2_ASAP7_75t_R _16285_ (.A1(_08737_),
    .A2(_09008_),
    .B(_09013_),
    .Y(_01463_));
 AOI22x1_ASAP7_75t_R _16286_ (.A1(_00217_),
    .A2(_09000_),
    .B1(_09009_),
    .B2(_08495_),
    .Y(_09014_));
 OA21x2_ASAP7_75t_R _16287_ (.A1(_08739_),
    .A2(_09008_),
    .B(_09014_),
    .Y(_01464_));
 AOI22x1_ASAP7_75t_R _16288_ (.A1(_00184_),
    .A2(_09000_),
    .B1(_09009_),
    .B2(_08512_),
    .Y(_09015_));
 OA21x2_ASAP7_75t_R _16289_ (.A1(_08741_),
    .A2(_09008_),
    .B(_09015_),
    .Y(_01465_));
 INVx1_ASAP7_75t_R _16290_ (.A(_00150_),
    .Y(_09016_));
 OA222x2_ASAP7_75t_R _16291_ (.A1(_09016_),
    .A2(_08984_),
    .B1(_08985_),
    .B2(_08744_),
    .C1(_08987_),
    .C2(_08518_),
    .Y(_01466_));
 AOI22x1_ASAP7_75t_R _16292_ (.A1(_00117_),
    .A2(_09006_),
    .B1(_09009_),
    .B2(_08546_),
    .Y(_09017_));
 OA21x2_ASAP7_75t_R _16293_ (.A1(_08745_),
    .A2(_09008_),
    .B(_09017_),
    .Y(_01467_));
 NOR2x1_ASAP7_75t_R _16294_ (.A(_01015_),
    .B(_08984_),
    .Y(_09018_));
 AO21x1_ASAP7_75t_R _16295_ (.A1(_08747_),
    .A2(_08984_),
    .B(_09018_),
    .Y(_01468_));
 BUFx4f_ASAP7_75t_R _16296_ (.A(_08989_),
    .Y(_09019_));
 AND3x1_ASAP7_75t_R _16297_ (.A(_08824_),
    .B(_08788_),
    .C(_09019_),
    .Y(_09020_));
 NOR2x1_ASAP7_75t_R _16298_ (.A(_00083_),
    .B(_08984_),
    .Y(_09021_));
 AO221x1_ASAP7_75t_R _16299_ (.A1(_08565_),
    .A2(_08984_),
    .B1(_09020_),
    .B2(_08752_),
    .C(_09021_),
    .Y(_01469_));
 AND2x2_ASAP7_75t_R _16300_ (.A(_00051_),
    .B(_09006_),
    .Y(_09022_));
 AOI221x1_ASAP7_75t_R _16301_ (.A1(_08591_),
    .A2(_09020_),
    .B1(_08993_),
    .B2(_08754_),
    .C(_09022_),
    .Y(_01470_));
 AOI22x1_ASAP7_75t_R _16302_ (.A1(_00982_),
    .A2(_09006_),
    .B1(_09009_),
    .B2(_08604_),
    .Y(_09023_));
 OA21x2_ASAP7_75t_R _16303_ (.A1(_08756_),
    .A2(_09008_),
    .B(_09023_),
    .Y(_01471_));
 NAND2x1_ASAP7_75t_R _16304_ (.A(_00949_),
    .B(_09006_),
    .Y(_09024_));
 OA221x2_ASAP7_75t_R _16305_ (.A1(_08758_),
    .A2(_08991_),
    .B1(_08985_),
    .B2(_08619_),
    .C(_09024_),
    .Y(_01472_));
 NAND2x1_ASAP7_75t_R _16306_ (.A(_00915_),
    .B(_09006_),
    .Y(_09025_));
 OA221x2_ASAP7_75t_R _16307_ (.A1(_08631_),
    .A2(_08991_),
    .B1(_08985_),
    .B2(_08760_),
    .C(_09025_),
    .Y(_01473_));
 AOI22x1_ASAP7_75t_R _16308_ (.A1(_00882_),
    .A2(_09006_),
    .B1(_09009_),
    .B2(_08644_),
    .Y(_09026_));
 OA21x2_ASAP7_75t_R _16309_ (.A1(_08762_),
    .A2(_09008_),
    .B(_09026_),
    .Y(_01474_));
 NAND2x1_ASAP7_75t_R _16310_ (.A(_00848_),
    .B(_08990_),
    .Y(_09027_));
 OA21x2_ASAP7_75t_R _16311_ (.A1(_08765_),
    .A2(_09006_),
    .B(_09027_),
    .Y(_09028_));
 OA21x2_ASAP7_75t_R _16312_ (.A1(_08764_),
    .A2(_09008_),
    .B(_09028_),
    .Y(_01475_));
 AOI22x1_ASAP7_75t_R _16313_ (.A1(_00815_),
    .A2(_09006_),
    .B1(_09009_),
    .B2(_08670_),
    .Y(_09029_));
 OA21x2_ASAP7_75t_R _16314_ (.A1(_08768_),
    .A2(_08985_),
    .B(_09029_),
    .Y(_01476_));
 NAND2x1_ASAP7_75t_R _16315_ (.A(_00781_),
    .B(_08990_),
    .Y(_09030_));
 OA21x2_ASAP7_75t_R _16316_ (.A1(_08771_),
    .A2(_09006_),
    .B(_09030_),
    .Y(_09031_));
 OA21x2_ASAP7_75t_R _16317_ (.A1(_08770_),
    .A2(_08985_),
    .B(_09031_),
    .Y(_01477_));
 AND2x6_ASAP7_75t_R _16318_ (.A(_08838_),
    .B(_08983_),
    .Y(_09032_));
 NAND2x2_ASAP7_75t_R _16319_ (.A(_08687_),
    .B(_09032_),
    .Y(_09033_));
 BUFx4f_ASAP7_75t_R _16320_ (.A(_09033_),
    .Y(_09034_));
 NAND2x2_ASAP7_75t_R _16321_ (.A(_08937_),
    .B(_09032_),
    .Y(_09035_));
 OA22x2_ASAP7_75t_R _16322_ (.A1(_03102_),
    .A2(_09032_),
    .B1(_09035_),
    .B2(_08793_),
    .Y(_09036_));
 OA21x2_ASAP7_75t_R _16323_ (.A1(_08093_),
    .A2(_09034_),
    .B(_09036_),
    .Y(_01478_));
 NAND2x2_ASAP7_75t_R _16324_ (.A(_08873_),
    .B(_08989_),
    .Y(_09037_));
 BUFx10_ASAP7_75t_R _16325_ (.A(_09037_),
    .Y(_09038_));
 AND3x2_ASAP7_75t_R _16326_ (.A(_08798_),
    .B(_08873_),
    .C(_08989_),
    .Y(_09039_));
 BUFx6f_ASAP7_75t_R _16327_ (.A(_09039_),
    .Y(_09040_));
 AOI22x1_ASAP7_75t_R _16328_ (.A1(_00749_),
    .A2(_09038_),
    .B1(_09040_),
    .B2(_08156_),
    .Y(_09041_));
 OA21x2_ASAP7_75t_R _16329_ (.A1(_08699_),
    .A2(_09034_),
    .B(_09041_),
    .Y(_01479_));
 AOI22x1_ASAP7_75t_R _16330_ (.A1(_00716_),
    .A2(_09038_),
    .B1(_09040_),
    .B2(_08185_),
    .Y(_09042_));
 OA21x2_ASAP7_75t_R _16331_ (.A1(_08705_),
    .A2(_09034_),
    .B(_09042_),
    .Y(_01480_));
 OA222x2_ASAP7_75t_R _16332_ (.A1(_05745_),
    .A2(_09032_),
    .B1(_09033_),
    .B2(_08707_),
    .C1(_09035_),
    .C2(_08191_),
    .Y(_01481_));
 INVx1_ASAP7_75t_R _16333_ (.A(_00650_),
    .Y(_09043_));
 OA222x2_ASAP7_75t_R _16334_ (.A1(_09043_),
    .A2(_09032_),
    .B1(_09033_),
    .B2(_08709_),
    .C1(_09035_),
    .C2(_08211_),
    .Y(_01482_));
 AOI22x1_ASAP7_75t_R _16335_ (.A1(_00617_),
    .A2(_09038_),
    .B1(_09040_),
    .B2(_08243_),
    .Y(_09044_));
 OA21x2_ASAP7_75t_R _16336_ (.A1(_08710_),
    .A2(_09034_),
    .B(_09044_),
    .Y(_01483_));
 AOI22x1_ASAP7_75t_R _16337_ (.A1(_00583_),
    .A2(_09038_),
    .B1(_09040_),
    .B2(_08259_),
    .Y(_09045_));
 OA21x2_ASAP7_75t_R _16338_ (.A1(_08712_),
    .A2(_09034_),
    .B(_09045_),
    .Y(_01484_));
 AOI22x1_ASAP7_75t_R _16339_ (.A1(_00550_),
    .A2(_09038_),
    .B1(_09040_),
    .B2(_08287_),
    .Y(_09046_));
 OA21x2_ASAP7_75t_R _16340_ (.A1(_08714_),
    .A2(_09034_),
    .B(_09046_),
    .Y(_01485_));
 AOI22x1_ASAP7_75t_R _16341_ (.A1(_00517_),
    .A2(_09038_),
    .B1(_09040_),
    .B2(_08308_),
    .Y(_09047_));
 OA21x2_ASAP7_75t_R _16342_ (.A1(_08716_),
    .A2(_09034_),
    .B(_09047_),
    .Y(_01486_));
 BUFx12_ASAP7_75t_R _16343_ (.A(_09037_),
    .Y(_09048_));
 AOI22x1_ASAP7_75t_R _16344_ (.A1(_00484_),
    .A2(_09048_),
    .B1(_09040_),
    .B2(_08327_),
    .Y(_09049_));
 OA21x2_ASAP7_75t_R _16345_ (.A1(_08719_),
    .A2(_09034_),
    .B(_09049_),
    .Y(_01487_));
 AOI22x1_ASAP7_75t_R _16346_ (.A1(_00451_),
    .A2(_09048_),
    .B1(_09040_),
    .B2(_08348_),
    .Y(_09050_));
 OA21x2_ASAP7_75t_R _16347_ (.A1(_08721_),
    .A2(_09034_),
    .B(_09050_),
    .Y(_01488_));
 BUFx10_ASAP7_75t_R _16348_ (.A(_08873_),
    .Y(_09051_));
 AO21x1_ASAP7_75t_R _16349_ (.A1(_09051_),
    .A2(_09019_),
    .B(_06771_),
    .Y(_09052_));
 OA21x2_ASAP7_75t_R _16350_ (.A1(_08723_),
    .A2(_09038_),
    .B(_09052_),
    .Y(_01489_));
 AOI22x1_ASAP7_75t_R _16351_ (.A1(_00418_),
    .A2(_09048_),
    .B1(_09040_),
    .B2(_08382_),
    .Y(_09053_));
 OA21x2_ASAP7_75t_R _16352_ (.A1(_08725_),
    .A2(_09034_),
    .B(_09053_),
    .Y(_01490_));
 AO21x1_ASAP7_75t_R _16353_ (.A1(_09051_),
    .A2(_09019_),
    .B(_04798_),
    .Y(_09054_));
 OA221x2_ASAP7_75t_R _16354_ (.A1(_08401_),
    .A2(_09038_),
    .B1(_09033_),
    .B2(_08727_),
    .C(_09054_),
    .Y(_01491_));
 BUFx4f_ASAP7_75t_R _16355_ (.A(_09033_),
    .Y(_09055_));
 BUFx6f_ASAP7_75t_R _16356_ (.A(_09039_),
    .Y(_09056_));
 AOI22x1_ASAP7_75t_R _16357_ (.A1(_00352_),
    .A2(_09048_),
    .B1(_09056_),
    .B2(_08420_),
    .Y(_09057_));
 OA21x2_ASAP7_75t_R _16358_ (.A1(_08729_),
    .A2(_09055_),
    .B(_09057_),
    .Y(_01492_));
 AOI22x1_ASAP7_75t_R _16359_ (.A1(_00318_),
    .A2(_09048_),
    .B1(_09056_),
    .B2(_08438_),
    .Y(_09058_));
 OA21x2_ASAP7_75t_R _16360_ (.A1(_08733_),
    .A2(_09055_),
    .B(_09058_),
    .Y(_01493_));
 AOI22x1_ASAP7_75t_R _16361_ (.A1(_00285_),
    .A2(_09048_),
    .B1(_09056_),
    .B2(_08459_),
    .Y(_09059_));
 OA21x2_ASAP7_75t_R _16362_ (.A1(_08735_),
    .A2(_09055_),
    .B(_09059_),
    .Y(_01494_));
 AOI22x1_ASAP7_75t_R _16363_ (.A1(_00252_),
    .A2(_09048_),
    .B1(_09056_),
    .B2(_08477_),
    .Y(_09060_));
 OA21x2_ASAP7_75t_R _16364_ (.A1(_08737_),
    .A2(_09055_),
    .B(_09060_),
    .Y(_01495_));
 AOI22x1_ASAP7_75t_R _16365_ (.A1(_00218_),
    .A2(_09048_),
    .B1(_09056_),
    .B2(_08495_),
    .Y(_09061_));
 OA21x2_ASAP7_75t_R _16366_ (.A1(_08739_),
    .A2(_09055_),
    .B(_09061_),
    .Y(_01496_));
 AOI22x1_ASAP7_75t_R _16367_ (.A1(_00185_),
    .A2(_09048_),
    .B1(_09056_),
    .B2(_08512_),
    .Y(_09062_));
 OA21x2_ASAP7_75t_R _16368_ (.A1(_08741_),
    .A2(_09055_),
    .B(_09062_),
    .Y(_01497_));
 INVx1_ASAP7_75t_R _16369_ (.A(_00151_),
    .Y(_09063_));
 OA222x2_ASAP7_75t_R _16370_ (.A1(_09063_),
    .A2(_09032_),
    .B1(_09033_),
    .B2(_08744_),
    .C1(_09035_),
    .C2(_08518_),
    .Y(_01498_));
 AOI22x1_ASAP7_75t_R _16371_ (.A1(_00118_),
    .A2(_09048_),
    .B1(_09056_),
    .B2(_08546_),
    .Y(_09064_));
 OA21x2_ASAP7_75t_R _16372_ (.A1(_08745_),
    .A2(_09055_),
    .B(_09064_),
    .Y(_01499_));
 NOR2x1_ASAP7_75t_R _16373_ (.A(_01016_),
    .B(_09032_),
    .Y(_09065_));
 AO21x1_ASAP7_75t_R _16374_ (.A1(_08747_),
    .A2(_09032_),
    .B(_09065_),
    .Y(_01500_));
 AND3x1_ASAP7_75t_R _16375_ (.A(_08824_),
    .B(_09051_),
    .C(_09019_),
    .Y(_09066_));
 NOR2x1_ASAP7_75t_R _16376_ (.A(_00084_),
    .B(_09032_),
    .Y(_09067_));
 AO221x1_ASAP7_75t_R _16377_ (.A1(_08565_),
    .A2(_09032_),
    .B1(_09066_),
    .B2(_08752_),
    .C(_09067_),
    .Y(_01501_));
 AND2x2_ASAP7_75t_R _16378_ (.A(_00052_),
    .B(_09037_),
    .Y(_09068_));
 AOI221x1_ASAP7_75t_R _16379_ (.A1(_08591_),
    .A2(_09066_),
    .B1(_09040_),
    .B2(_08754_),
    .C(_09068_),
    .Y(_01502_));
 AOI22x1_ASAP7_75t_R _16380_ (.A1(_00983_),
    .A2(_09037_),
    .B1(_09056_),
    .B2(_08604_),
    .Y(_09069_));
 OA21x2_ASAP7_75t_R _16381_ (.A1(_08756_),
    .A2(_09055_),
    .B(_09069_),
    .Y(_01503_));
 NAND2x1_ASAP7_75t_R _16382_ (.A(_00950_),
    .B(_09037_),
    .Y(_09070_));
 OA221x2_ASAP7_75t_R _16383_ (.A1(_08758_),
    .A2(_09038_),
    .B1(_09033_),
    .B2(_08619_),
    .C(_09070_),
    .Y(_01504_));
 AO21x1_ASAP7_75t_R _16384_ (.A1(_09051_),
    .A2(_09019_),
    .B(_06393_),
    .Y(_09071_));
 OA221x2_ASAP7_75t_R _16385_ (.A1(_08631_),
    .A2(_09038_),
    .B1(_09033_),
    .B2(_08760_),
    .C(_09071_),
    .Y(_01505_));
 AOI22x1_ASAP7_75t_R _16386_ (.A1(_00883_),
    .A2(_09037_),
    .B1(_09056_),
    .B2(_08644_),
    .Y(_09072_));
 OA21x2_ASAP7_75t_R _16387_ (.A1(_08762_),
    .A2(_09055_),
    .B(_09072_),
    .Y(_01506_));
 AO21x1_ASAP7_75t_R _16388_ (.A1(_08873_),
    .A2(_08989_),
    .B(_06219_),
    .Y(_09073_));
 OA21x2_ASAP7_75t_R _16389_ (.A1(_08765_),
    .A2(_09037_),
    .B(_09073_),
    .Y(_09074_));
 OA21x2_ASAP7_75t_R _16390_ (.A1(_08764_),
    .A2(_09055_),
    .B(_09074_),
    .Y(_01507_));
 AOI22x1_ASAP7_75t_R _16391_ (.A1(_00816_),
    .A2(_09037_),
    .B1(_09056_),
    .B2(_08670_),
    .Y(_09075_));
 OA21x2_ASAP7_75t_R _16392_ (.A1(_08768_),
    .A2(_09033_),
    .B(_09075_),
    .Y(_01508_));
 NAND2x1_ASAP7_75t_R _16393_ (.A(_00782_),
    .B(_09037_),
    .Y(_09076_));
 OA21x2_ASAP7_75t_R _16394_ (.A1(_08771_),
    .A2(_09037_),
    .B(_09076_),
    .Y(_09077_));
 OA21x2_ASAP7_75t_R _16395_ (.A1(_08770_),
    .A2(_09033_),
    .B(_09077_),
    .Y(_01509_));
 AND2x6_ASAP7_75t_R _16396_ (.A(_08098_),
    .B(_08983_),
    .Y(_09078_));
 NAND2x2_ASAP7_75t_R _16397_ (.A(_08687_),
    .B(_09078_),
    .Y(_09079_));
 BUFx4f_ASAP7_75t_R _16398_ (.A(_09079_),
    .Y(_09080_));
 NAND2x2_ASAP7_75t_R _16399_ (.A(_08115_),
    .B(_09078_),
    .Y(_09081_));
 NAND2x2_ASAP7_75t_R _16400_ (.A(_08117_),
    .B(_08983_),
    .Y(_09082_));
 NAND2x1_ASAP7_75t_R _16401_ (.A(_00018_),
    .B(_09082_),
    .Y(_09083_));
 OA21x2_ASAP7_75t_R _16402_ (.A1(_08111_),
    .A2(_09081_),
    .B(_09083_),
    .Y(_09084_));
 OA21x2_ASAP7_75t_R _16403_ (.A1(_08093_),
    .A2(_09080_),
    .B(_09084_),
    .Y(_01510_));
 BUFx10_ASAP7_75t_R _16404_ (.A(_09082_),
    .Y(_09085_));
 AND3x2_ASAP7_75t_R _16405_ (.A(_08117_),
    .B(_08701_),
    .C(_08989_),
    .Y(_09086_));
 BUFx10_ASAP7_75t_R _16406_ (.A(_09086_),
    .Y(_09087_));
 AOI22x1_ASAP7_75t_R _16407_ (.A1(_00750_),
    .A2(_09085_),
    .B1(_09087_),
    .B2(_08156_),
    .Y(_09088_));
 OA21x2_ASAP7_75t_R _16408_ (.A1(_08699_),
    .A2(_09080_),
    .B(_09088_),
    .Y(_01511_));
 AOI22x1_ASAP7_75t_R _16409_ (.A1(_00717_),
    .A2(_09085_),
    .B1(_09087_),
    .B2(_08185_),
    .Y(_09089_));
 OA21x2_ASAP7_75t_R _16410_ (.A1(_08705_),
    .A2(_09080_),
    .B(_09089_),
    .Y(_01512_));
 OA222x2_ASAP7_75t_R _16411_ (.A1(_05749_),
    .A2(_09078_),
    .B1(_09079_),
    .B2(_08707_),
    .C1(_09081_),
    .C2(_08191_),
    .Y(_01513_));
 OA222x2_ASAP7_75t_R _16412_ (.A1(_05625_),
    .A2(_09078_),
    .B1(_09079_),
    .B2(_08709_),
    .C1(_09081_),
    .C2(_08211_),
    .Y(_01514_));
 AOI22x1_ASAP7_75t_R _16413_ (.A1(_00618_),
    .A2(_09085_),
    .B1(_09087_),
    .B2(_08243_),
    .Y(_09090_));
 OA21x2_ASAP7_75t_R _16414_ (.A1(_08710_),
    .A2(_09080_),
    .B(_09090_),
    .Y(_01515_));
 AOI22x1_ASAP7_75t_R _16415_ (.A1(_00584_),
    .A2(_09085_),
    .B1(_09087_),
    .B2(_08259_),
    .Y(_09091_));
 OA21x2_ASAP7_75t_R _16416_ (.A1(_08712_),
    .A2(_09080_),
    .B(_09091_),
    .Y(_01516_));
 AOI22x1_ASAP7_75t_R _16417_ (.A1(_00551_),
    .A2(_09085_),
    .B1(_09087_),
    .B2(_08287_),
    .Y(_09092_));
 OA21x2_ASAP7_75t_R _16418_ (.A1(_08714_),
    .A2(_09080_),
    .B(_09092_),
    .Y(_01517_));
 BUFx12_ASAP7_75t_R _16419_ (.A(_09082_),
    .Y(_09093_));
 AOI22x1_ASAP7_75t_R _16420_ (.A1(_00518_),
    .A2(_09093_),
    .B1(_09087_),
    .B2(_08308_),
    .Y(_09094_));
 OA21x2_ASAP7_75t_R _16421_ (.A1(_08716_),
    .A2(_09080_),
    .B(_09094_),
    .Y(_01518_));
 AOI22x1_ASAP7_75t_R _16422_ (.A1(_00485_),
    .A2(_09093_),
    .B1(_09087_),
    .B2(_08327_),
    .Y(_09095_));
 OA21x2_ASAP7_75t_R _16423_ (.A1(_08719_),
    .A2(_09080_),
    .B(_09095_),
    .Y(_01519_));
 AOI22x1_ASAP7_75t_R _16424_ (.A1(_00452_),
    .A2(_09093_),
    .B1(_09087_),
    .B2(_08348_),
    .Y(_09096_));
 OA21x2_ASAP7_75t_R _16425_ (.A1(_08721_),
    .A2(_09080_),
    .B(_09096_),
    .Y(_01520_));
 NAND2x1_ASAP7_75t_R _16426_ (.A(_01050_),
    .B(_09085_),
    .Y(_09097_));
 OA21x2_ASAP7_75t_R _16427_ (.A1(_08723_),
    .A2(_09085_),
    .B(_09097_),
    .Y(_01521_));
 AOI22x1_ASAP7_75t_R _16428_ (.A1(_00419_),
    .A2(_09093_),
    .B1(_09087_),
    .B2(_08382_),
    .Y(_09098_));
 OA21x2_ASAP7_75t_R _16429_ (.A1(_08725_),
    .A2(_09080_),
    .B(_09098_),
    .Y(_01522_));
 BUFx6f_ASAP7_75t_R _16430_ (.A(_09082_),
    .Y(_09099_));
 NAND2x1_ASAP7_75t_R _16431_ (.A(_00386_),
    .B(_09099_),
    .Y(_09100_));
 OA221x2_ASAP7_75t_R _16432_ (.A1(_08401_),
    .A2(_09085_),
    .B1(_09079_),
    .B2(_08727_),
    .C(_09100_),
    .Y(_01523_));
 BUFx6f_ASAP7_75t_R _16433_ (.A(_09079_),
    .Y(_09101_));
 BUFx10_ASAP7_75t_R _16434_ (.A(_09086_),
    .Y(_09102_));
 AOI22x1_ASAP7_75t_R _16435_ (.A1(_00353_),
    .A2(_09093_),
    .B1(_09102_),
    .B2(_08420_),
    .Y(_09103_));
 OA21x2_ASAP7_75t_R _16436_ (.A1(_08729_),
    .A2(_09101_),
    .B(_09103_),
    .Y(_01524_));
 AOI22x1_ASAP7_75t_R _16437_ (.A1(_00319_),
    .A2(_09093_),
    .B1(_09102_),
    .B2(_08438_),
    .Y(_09104_));
 OA21x2_ASAP7_75t_R _16438_ (.A1(_08733_),
    .A2(_09101_),
    .B(_09104_),
    .Y(_01525_));
 AOI22x1_ASAP7_75t_R _16439_ (.A1(_00286_),
    .A2(_09093_),
    .B1(_09102_),
    .B2(_08459_),
    .Y(_09105_));
 OA21x2_ASAP7_75t_R _16440_ (.A1(_08735_),
    .A2(_09101_),
    .B(_09105_),
    .Y(_01526_));
 AOI22x1_ASAP7_75t_R _16441_ (.A1(_00253_),
    .A2(_09093_),
    .B1(_09102_),
    .B2(_08477_),
    .Y(_09106_));
 OA21x2_ASAP7_75t_R _16442_ (.A1(_08737_),
    .A2(_09101_),
    .B(_09106_),
    .Y(_01527_));
 AOI22x1_ASAP7_75t_R _16443_ (.A1(_00219_),
    .A2(_09093_),
    .B1(_09102_),
    .B2(_08495_),
    .Y(_09107_));
 OA21x2_ASAP7_75t_R _16444_ (.A1(_08739_),
    .A2(_09101_),
    .B(_09107_),
    .Y(_01528_));
 AOI22x1_ASAP7_75t_R _16445_ (.A1(_00186_),
    .A2(_09093_),
    .B1(_09102_),
    .B2(_08512_),
    .Y(_09108_));
 OA21x2_ASAP7_75t_R _16446_ (.A1(_08741_),
    .A2(_09101_),
    .B(_09108_),
    .Y(_01529_));
 OA222x2_ASAP7_75t_R _16447_ (.A1(_03966_),
    .A2(_09078_),
    .B1(_09079_),
    .B2(_08744_),
    .C1(_09081_),
    .C2(_08518_),
    .Y(_01530_));
 AOI22x1_ASAP7_75t_R _16448_ (.A1(_00119_),
    .A2(_09099_),
    .B1(_09102_),
    .B2(_08546_),
    .Y(_09109_));
 OA21x2_ASAP7_75t_R _16449_ (.A1(_08745_),
    .A2(_09101_),
    .B(_09109_),
    .Y(_01531_));
 NOR2x1_ASAP7_75t_R _16450_ (.A(_01017_),
    .B(_09078_),
    .Y(_09110_));
 AO21x1_ASAP7_75t_R _16451_ (.A1(_08747_),
    .A2(_09078_),
    .B(_09110_),
    .Y(_01532_));
 AND3x1_ASAP7_75t_R _16452_ (.A(_08145_),
    .B(_08577_),
    .C(_09019_),
    .Y(_09111_));
 NOR2x1_ASAP7_75t_R _16453_ (.A(_00085_),
    .B(_09078_),
    .Y(_09112_));
 AO221x1_ASAP7_75t_R _16454_ (.A1(_08565_),
    .A2(_09078_),
    .B1(_09111_),
    .B2(_08752_),
    .C(_09112_),
    .Y(_01533_));
 AND2x2_ASAP7_75t_R _16455_ (.A(_00053_),
    .B(_09099_),
    .Y(_09113_));
 AOI221x1_ASAP7_75t_R _16456_ (.A1(_08591_),
    .A2(_09111_),
    .B1(_09087_),
    .B2(_08754_),
    .C(_09113_),
    .Y(_01534_));
 AOI22x1_ASAP7_75t_R _16457_ (.A1(_00984_),
    .A2(_09099_),
    .B1(_09102_),
    .B2(_08604_),
    .Y(_09114_));
 OA21x2_ASAP7_75t_R _16458_ (.A1(_08756_),
    .A2(_09101_),
    .B(_09114_),
    .Y(_01535_));
 NAND2x1_ASAP7_75t_R _16459_ (.A(_00951_),
    .B(_09099_),
    .Y(_09115_));
 OA221x2_ASAP7_75t_R _16460_ (.A1(_08758_),
    .A2(_09085_),
    .B1(_09079_),
    .B2(_08619_),
    .C(_09115_),
    .Y(_01536_));
 NAND2x1_ASAP7_75t_R _16461_ (.A(_00917_),
    .B(_09099_),
    .Y(_09116_));
 OA221x2_ASAP7_75t_R _16462_ (.A1(_08631_),
    .A2(_09085_),
    .B1(_09079_),
    .B2(_08760_),
    .C(_09116_),
    .Y(_01537_));
 AOI22x1_ASAP7_75t_R _16463_ (.A1(_00884_),
    .A2(_09099_),
    .B1(_09102_),
    .B2(_08644_),
    .Y(_09117_));
 OA21x2_ASAP7_75t_R _16464_ (.A1(_08762_),
    .A2(_09101_),
    .B(_09117_),
    .Y(_01538_));
 NAND2x1_ASAP7_75t_R _16465_ (.A(_00850_),
    .B(_09082_),
    .Y(_09118_));
 OA21x2_ASAP7_75t_R _16466_ (.A1(_08765_),
    .A2(_09099_),
    .B(_09118_),
    .Y(_09119_));
 OA21x2_ASAP7_75t_R _16467_ (.A1(_08764_),
    .A2(_09101_),
    .B(_09119_),
    .Y(_01539_));
 AOI22x1_ASAP7_75t_R _16468_ (.A1(_00817_),
    .A2(_09099_),
    .B1(_09102_),
    .B2(_08670_),
    .Y(_09120_));
 OA21x2_ASAP7_75t_R _16469_ (.A1(_08768_),
    .A2(_09079_),
    .B(_09120_),
    .Y(_01540_));
 NAND2x1_ASAP7_75t_R _16470_ (.A(_00783_),
    .B(_09082_),
    .Y(_09121_));
 OA21x2_ASAP7_75t_R _16471_ (.A1(_08771_),
    .A2(_09099_),
    .B(_09121_),
    .Y(_09122_));
 OA21x2_ASAP7_75t_R _16472_ (.A1(_08770_),
    .A2(_09079_),
    .B(_09122_),
    .Y(_01541_));
 AND2x6_ASAP7_75t_R _16473_ (.A(_08689_),
    .B(_08983_),
    .Y(_09123_));
 NAND2x2_ASAP7_75t_R _16474_ (.A(_08687_),
    .B(_09123_),
    .Y(_09124_));
 BUFx4f_ASAP7_75t_R _16475_ (.A(_09124_),
    .Y(_09125_));
 NAND2x2_ASAP7_75t_R _16476_ (.A(_08937_),
    .B(_09123_),
    .Y(_09126_));
 OA22x2_ASAP7_75t_R _16477_ (.A1(_03101_),
    .A2(_09123_),
    .B1(_09126_),
    .B2(_08793_),
    .Y(_09127_));
 OA21x2_ASAP7_75t_R _16478_ (.A1(_08093_),
    .A2(_09125_),
    .B(_09127_),
    .Y(_01542_));
 NAND2x2_ASAP7_75t_R _16479_ (.A(_08749_),
    .B(_08989_),
    .Y(_09128_));
 BUFx12_ASAP7_75t_R _16480_ (.A(_09128_),
    .Y(_09129_));
 AND3x2_ASAP7_75t_R _16481_ (.A(_08798_),
    .B(_08749_),
    .C(_08989_),
    .Y(_09130_));
 BUFx6f_ASAP7_75t_R _16482_ (.A(_09130_),
    .Y(_09131_));
 AOI22x1_ASAP7_75t_R _16483_ (.A1(_00751_),
    .A2(_09129_),
    .B1(_09131_),
    .B2(_08156_),
    .Y(_09132_));
 OA21x2_ASAP7_75t_R _16484_ (.A1(_08699_),
    .A2(_09125_),
    .B(_09132_),
    .Y(_01543_));
 AOI22x1_ASAP7_75t_R _16485_ (.A1(_00718_),
    .A2(_09129_),
    .B1(_09131_),
    .B2(_08185_),
    .Y(_09133_));
 OA21x2_ASAP7_75t_R _16486_ (.A1(_08705_),
    .A2(_09125_),
    .B(_09133_),
    .Y(_01544_));
 OA222x2_ASAP7_75t_R _16487_ (.A1(_05750_),
    .A2(_09123_),
    .B1(_09124_),
    .B2(_08707_),
    .C1(_09126_),
    .C2(_08191_),
    .Y(_01545_));
 OA222x2_ASAP7_75t_R _16488_ (.A1(_05626_),
    .A2(_09123_),
    .B1(_09124_),
    .B2(_08709_),
    .C1(_09126_),
    .C2(_08211_),
    .Y(_01546_));
 AOI22x1_ASAP7_75t_R _16489_ (.A1(_00619_),
    .A2(_09129_),
    .B1(_09131_),
    .B2(_08243_),
    .Y(_09134_));
 OA21x2_ASAP7_75t_R _16490_ (.A1(_08710_),
    .A2(_09125_),
    .B(_09134_),
    .Y(_01547_));
 AOI22x1_ASAP7_75t_R _16491_ (.A1(_00585_),
    .A2(_09129_),
    .B1(_09131_),
    .B2(_08259_),
    .Y(_09135_));
 OA21x2_ASAP7_75t_R _16492_ (.A1(_08712_),
    .A2(_09125_),
    .B(_09135_),
    .Y(_01548_));
 AOI22x1_ASAP7_75t_R _16493_ (.A1(_00552_),
    .A2(_09129_),
    .B1(_09131_),
    .B2(_08287_),
    .Y(_09136_));
 OA21x2_ASAP7_75t_R _16494_ (.A1(_08714_),
    .A2(_09125_),
    .B(_09136_),
    .Y(_01549_));
 AOI22x1_ASAP7_75t_R _16495_ (.A1(_00519_),
    .A2(_09129_),
    .B1(_09131_),
    .B2(_08308_),
    .Y(_09137_));
 OA21x2_ASAP7_75t_R _16496_ (.A1(_08716_),
    .A2(_09125_),
    .B(_09137_),
    .Y(_01550_));
 BUFx12_ASAP7_75t_R _16497_ (.A(_09128_),
    .Y(_09138_));
 AOI22x1_ASAP7_75t_R _16498_ (.A1(_00486_),
    .A2(_09138_),
    .B1(_09131_),
    .B2(_08327_),
    .Y(_09139_));
 OA21x2_ASAP7_75t_R _16499_ (.A1(_08719_),
    .A2(_09125_),
    .B(_09139_),
    .Y(_01551_));
 AOI22x1_ASAP7_75t_R _16500_ (.A1(_00453_),
    .A2(_09138_),
    .B1(_09131_),
    .B2(_08348_),
    .Y(_09140_));
 OA21x2_ASAP7_75t_R _16501_ (.A1(_08721_),
    .A2(_09125_),
    .B(_09140_),
    .Y(_01552_));
 BUFx6f_ASAP7_75t_R _16502_ (.A(_08749_),
    .Y(_09141_));
 AO21x1_ASAP7_75t_R _16503_ (.A1(_09141_),
    .A2(_09019_),
    .B(_06776_),
    .Y(_09142_));
 OA21x2_ASAP7_75t_R _16504_ (.A1(_08723_),
    .A2(_09129_),
    .B(_09142_),
    .Y(_01553_));
 AOI22x1_ASAP7_75t_R _16505_ (.A1(_00420_),
    .A2(_09138_),
    .B1(_09131_),
    .B2(_08382_),
    .Y(_09143_));
 OA21x2_ASAP7_75t_R _16506_ (.A1(_08725_),
    .A2(_09125_),
    .B(_09143_),
    .Y(_01554_));
 AO21x1_ASAP7_75t_R _16507_ (.A1(_09141_),
    .A2(_09019_),
    .B(_04803_),
    .Y(_09144_));
 OA221x2_ASAP7_75t_R _16508_ (.A1(_08401_),
    .A2(_09129_),
    .B1(_09124_),
    .B2(_08727_),
    .C(_09144_),
    .Y(_01555_));
 BUFx4f_ASAP7_75t_R _16509_ (.A(_09124_),
    .Y(_09145_));
 BUFx10_ASAP7_75t_R _16510_ (.A(_09130_),
    .Y(_09146_));
 AOI22x1_ASAP7_75t_R _16511_ (.A1(_00354_),
    .A2(_09138_),
    .B1(_09146_),
    .B2(_08420_),
    .Y(_09147_));
 OA21x2_ASAP7_75t_R _16512_ (.A1(_08729_),
    .A2(_09145_),
    .B(_09147_),
    .Y(_01556_));
 AOI22x1_ASAP7_75t_R _16513_ (.A1(_00320_),
    .A2(_09138_),
    .B1(_09146_),
    .B2(_08438_),
    .Y(_09148_));
 OA21x2_ASAP7_75t_R _16514_ (.A1(_08733_),
    .A2(_09145_),
    .B(_09148_),
    .Y(_01557_));
 AOI22x1_ASAP7_75t_R _16515_ (.A1(_00287_),
    .A2(_09138_),
    .B1(_09146_),
    .B2(_08459_),
    .Y(_09149_));
 OA21x2_ASAP7_75t_R _16516_ (.A1(_08735_),
    .A2(_09145_),
    .B(_09149_),
    .Y(_01558_));
 AOI22x1_ASAP7_75t_R _16517_ (.A1(_00254_),
    .A2(_09138_),
    .B1(_09146_),
    .B2(_08477_),
    .Y(_09150_));
 OA21x2_ASAP7_75t_R _16518_ (.A1(_08737_),
    .A2(_09145_),
    .B(_09150_),
    .Y(_01559_));
 AOI22x1_ASAP7_75t_R _16519_ (.A1(_00220_),
    .A2(_09138_),
    .B1(_09146_),
    .B2(_08495_),
    .Y(_09151_));
 OA21x2_ASAP7_75t_R _16520_ (.A1(_08739_),
    .A2(_09145_),
    .B(_09151_),
    .Y(_01560_));
 AOI22x1_ASAP7_75t_R _16521_ (.A1(_00187_),
    .A2(_09138_),
    .B1(_09146_),
    .B2(_08512_),
    .Y(_09152_));
 OA21x2_ASAP7_75t_R _16522_ (.A1(_08741_),
    .A2(_09145_),
    .B(_09152_),
    .Y(_01561_));
 OA222x2_ASAP7_75t_R _16523_ (.A1(_03967_),
    .A2(_09123_),
    .B1(_09124_),
    .B2(_08744_),
    .C1(_09126_),
    .C2(_08518_),
    .Y(_01562_));
 AOI22x1_ASAP7_75t_R _16524_ (.A1(_00120_),
    .A2(_09138_),
    .B1(_09146_),
    .B2(_08546_),
    .Y(_09153_));
 OA21x2_ASAP7_75t_R _16525_ (.A1(_08745_),
    .A2(_09145_),
    .B(_09153_),
    .Y(_01563_));
 NOR2x1_ASAP7_75t_R _16526_ (.A(_01018_),
    .B(_09123_),
    .Y(_09154_));
 AO21x1_ASAP7_75t_R _16527_ (.A1(_08747_),
    .A2(_09123_),
    .B(_09154_),
    .Y(_01564_));
 AND3x1_ASAP7_75t_R _16528_ (.A(_08824_),
    .B(_08750_),
    .C(_08989_),
    .Y(_09155_));
 NOR2x1_ASAP7_75t_R _16529_ (.A(_00086_),
    .B(_09123_),
    .Y(_09156_));
 AO221x1_ASAP7_75t_R _16530_ (.A1(_08565_),
    .A2(_09123_),
    .B1(_09155_),
    .B2(_08752_),
    .C(_09156_),
    .Y(_01565_));
 AND2x2_ASAP7_75t_R _16531_ (.A(_00054_),
    .B(_09128_),
    .Y(_09157_));
 AOI221x1_ASAP7_75t_R _16532_ (.A1(_08591_),
    .A2(_09155_),
    .B1(_09131_),
    .B2(_08754_),
    .C(_09157_),
    .Y(_01566_));
 AOI22x1_ASAP7_75t_R _16533_ (.A1(_00985_),
    .A2(_09128_),
    .B1(_09146_),
    .B2(_08604_),
    .Y(_09158_));
 OA21x2_ASAP7_75t_R _16534_ (.A1(_08756_),
    .A2(_09145_),
    .B(_09158_),
    .Y(_01567_));
 AO21x1_ASAP7_75t_R _16535_ (.A1(_09141_),
    .A2(_09019_),
    .B(_06500_),
    .Y(_09159_));
 OA221x2_ASAP7_75t_R _16536_ (.A1(_08758_),
    .A2(_09129_),
    .B1(_09124_),
    .B2(_08619_),
    .C(_09159_),
    .Y(_01568_));
 AO21x1_ASAP7_75t_R _16537_ (.A1(_09141_),
    .A2(_09019_),
    .B(_06400_),
    .Y(_09160_));
 OA221x2_ASAP7_75t_R _16538_ (.A1(_08631_),
    .A2(_09129_),
    .B1(_09124_),
    .B2(_08760_),
    .C(_09160_),
    .Y(_01569_));
 AOI22x1_ASAP7_75t_R _16539_ (.A1(_00885_),
    .A2(_09128_),
    .B1(_09146_),
    .B2(_08644_),
    .Y(_09161_));
 OA21x2_ASAP7_75t_R _16540_ (.A1(_08762_),
    .A2(_09145_),
    .B(_09161_),
    .Y(_01570_));
 NAND2x1_ASAP7_75t_R _16541_ (.A(_00851_),
    .B(_09128_),
    .Y(_09162_));
 OA21x2_ASAP7_75t_R _16542_ (.A1(_08765_),
    .A2(_09128_),
    .B(_09162_),
    .Y(_09163_));
 OA21x2_ASAP7_75t_R _16543_ (.A1(_08764_),
    .A2(_09145_),
    .B(_09163_),
    .Y(_01571_));
 AOI22x1_ASAP7_75t_R _16544_ (.A1(_00818_),
    .A2(_09128_),
    .B1(_09146_),
    .B2(_08670_),
    .Y(_09164_));
 OA21x2_ASAP7_75t_R _16545_ (.A1(_08768_),
    .A2(_09124_),
    .B(_09164_),
    .Y(_01572_));
 NAND2x1_ASAP7_75t_R _16546_ (.A(_00784_),
    .B(_09128_),
    .Y(_09165_));
 OA21x2_ASAP7_75t_R _16547_ (.A1(_08771_),
    .A2(_09128_),
    .B(_09165_),
    .Y(_09166_));
 OA21x2_ASAP7_75t_R _16548_ (.A1(_08770_),
    .A2(_09124_),
    .B(_09166_),
    .Y(_01573_));
 BUFx6f_ASAP7_75t_R _16549_ (.A(_08092_),
    .Y(_09167_));
 AND2x6_ASAP7_75t_R _16550_ (.A(_08777_),
    .B(_08838_),
    .Y(_09168_));
 NAND2x2_ASAP7_75t_R _16551_ (.A(_08687_),
    .B(_09168_),
    .Y(_09169_));
 BUFx6f_ASAP7_75t_R _16552_ (.A(_09169_),
    .Y(_09170_));
 NAND2x2_ASAP7_75t_R _16553_ (.A(_08937_),
    .B(_09168_),
    .Y(_09171_));
 OA22x2_ASAP7_75t_R _16554_ (.A1(_03084_),
    .A2(_09168_),
    .B1(_09171_),
    .B2(_08793_),
    .Y(_09172_));
 OA21x2_ASAP7_75t_R _16555_ (.A1(_09167_),
    .A2(_09170_),
    .B(_09172_),
    .Y(_01574_));
 NAND2x2_ASAP7_75t_R _16556_ (.A(_08777_),
    .B(_08838_),
    .Y(_09173_));
 BUFx12_ASAP7_75t_R _16557_ (.A(_09173_),
    .Y(_09174_));
 BUFx6f_ASAP7_75t_R _16558_ (.A(_08777_),
    .Y(_09175_));
 AND3x2_ASAP7_75t_R _16559_ (.A(_08798_),
    .B(_09175_),
    .C(_08847_),
    .Y(_09176_));
 BUFx10_ASAP7_75t_R _16560_ (.A(_09176_),
    .Y(_09177_));
 BUFx10_ASAP7_75t_R _16561_ (.A(_08155_),
    .Y(_09178_));
 AOI22x1_ASAP7_75t_R _16562_ (.A1(_00733_),
    .A2(_09174_),
    .B1(_09177_),
    .B2(_09178_),
    .Y(_09179_));
 OA21x2_ASAP7_75t_R _16563_ (.A1(_08699_),
    .A2(_09170_),
    .B(_09179_),
    .Y(_01575_));
 BUFx10_ASAP7_75t_R _16564_ (.A(_08184_),
    .Y(_09180_));
 AOI22x1_ASAP7_75t_R _16565_ (.A1(_00700_),
    .A2(_09174_),
    .B1(_09177_),
    .B2(_09180_),
    .Y(_09181_));
 OA21x2_ASAP7_75t_R _16566_ (.A1(_08705_),
    .A2(_09170_),
    .B(_09181_),
    .Y(_01576_));
 BUFx6f_ASAP7_75t_R _16567_ (.A(_08190_),
    .Y(_09182_));
 OA222x2_ASAP7_75t_R _16568_ (.A1(_05725_),
    .A2(_09168_),
    .B1(_09169_),
    .B2(_08707_),
    .C1(_09171_),
    .C2(_09182_),
    .Y(_01577_));
 INVx1_ASAP7_75t_R _16569_ (.A(_00634_),
    .Y(_09183_));
 BUFx6f_ASAP7_75t_R _16570_ (.A(_08210_),
    .Y(_09184_));
 OA222x2_ASAP7_75t_R _16571_ (.A1(_09183_),
    .A2(_09168_),
    .B1(_09169_),
    .B2(_08709_),
    .C1(_09171_),
    .C2(_09184_),
    .Y(_01578_));
 BUFx10_ASAP7_75t_R _16572_ (.A(_08242_),
    .Y(_09185_));
 AOI22x1_ASAP7_75t_R _16573_ (.A1(_00601_),
    .A2(_09174_),
    .B1(_09177_),
    .B2(_09185_),
    .Y(_09186_));
 OA21x2_ASAP7_75t_R _16574_ (.A1(_08710_),
    .A2(_09170_),
    .B(_09186_),
    .Y(_01579_));
 BUFx10_ASAP7_75t_R _16575_ (.A(_08258_),
    .Y(_09187_));
 AOI22x1_ASAP7_75t_R _16576_ (.A1(_00567_),
    .A2(_09174_),
    .B1(_09177_),
    .B2(_09187_),
    .Y(_09188_));
 OA21x2_ASAP7_75t_R _16577_ (.A1(_08712_),
    .A2(_09170_),
    .B(_09188_),
    .Y(_01580_));
 BUFx10_ASAP7_75t_R _16578_ (.A(_08286_),
    .Y(_09189_));
 AOI22x1_ASAP7_75t_R _16579_ (.A1(_00534_),
    .A2(_09174_),
    .B1(_09177_),
    .B2(_09189_),
    .Y(_09190_));
 OA21x2_ASAP7_75t_R _16580_ (.A1(_08714_),
    .A2(_09170_),
    .B(_09190_),
    .Y(_01581_));
 BUFx12_ASAP7_75t_R _16581_ (.A(_09173_),
    .Y(_09191_));
 BUFx12f_ASAP7_75t_R _16582_ (.A(_08307_),
    .Y(_09192_));
 AOI22x1_ASAP7_75t_R _16583_ (.A1(_00501_),
    .A2(_09191_),
    .B1(_09177_),
    .B2(_09192_),
    .Y(_09193_));
 OA21x2_ASAP7_75t_R _16584_ (.A1(_08716_),
    .A2(_09170_),
    .B(_09193_),
    .Y(_01582_));
 BUFx10_ASAP7_75t_R _16585_ (.A(_08326_),
    .Y(_09194_));
 AOI22x1_ASAP7_75t_R _16586_ (.A1(_00468_),
    .A2(_09191_),
    .B1(_09177_),
    .B2(_09194_),
    .Y(_09195_));
 OA21x2_ASAP7_75t_R _16587_ (.A1(_08719_),
    .A2(_09170_),
    .B(_09195_),
    .Y(_01583_));
 BUFx12_ASAP7_75t_R _16588_ (.A(_08347_),
    .Y(_09196_));
 AOI22x1_ASAP7_75t_R _16589_ (.A1(_00435_),
    .A2(_09191_),
    .B1(_09177_),
    .B2(_09196_),
    .Y(_09197_));
 OA21x2_ASAP7_75t_R _16590_ (.A1(_08721_),
    .A2(_09170_),
    .B(_09197_),
    .Y(_01584_));
 NAND2x1_ASAP7_75t_R _16591_ (.A(_01033_),
    .B(_09174_),
    .Y(_09198_));
 OA21x2_ASAP7_75t_R _16592_ (.A1(_08723_),
    .A2(_09174_),
    .B(_09198_),
    .Y(_01585_));
 BUFx12_ASAP7_75t_R _16593_ (.A(_08381_),
    .Y(_09199_));
 AOI22x1_ASAP7_75t_R _16594_ (.A1(_00402_),
    .A2(_09191_),
    .B1(_09177_),
    .B2(_09199_),
    .Y(_09200_));
 OA21x2_ASAP7_75t_R _16595_ (.A1(_08725_),
    .A2(_09170_),
    .B(_09200_),
    .Y(_01586_));
 BUFx10_ASAP7_75t_R _16596_ (.A(_08400_),
    .Y(_09201_));
 BUFx6f_ASAP7_75t_R _16597_ (.A(_09173_),
    .Y(_09202_));
 NAND2x1_ASAP7_75t_R _16598_ (.A(_00369_),
    .B(_09202_),
    .Y(_09203_));
 OA221x2_ASAP7_75t_R _16599_ (.A1(_09201_),
    .A2(_09174_),
    .B1(_09169_),
    .B2(_08727_),
    .C(_09203_),
    .Y(_01587_));
 BUFx4f_ASAP7_75t_R _16600_ (.A(_09169_),
    .Y(_09204_));
 BUFx6f_ASAP7_75t_R _16601_ (.A(_09176_),
    .Y(_09205_));
 BUFx10_ASAP7_75t_R _16602_ (.A(_08419_),
    .Y(_09206_));
 AOI22x1_ASAP7_75t_R _16603_ (.A1(_00336_),
    .A2(_09191_),
    .B1(_09205_),
    .B2(_09206_),
    .Y(_09207_));
 OA21x2_ASAP7_75t_R _16604_ (.A1(_08729_),
    .A2(_09204_),
    .B(_09207_),
    .Y(_01588_));
 BUFx12_ASAP7_75t_R _16605_ (.A(_08437_),
    .Y(_09208_));
 AOI22x1_ASAP7_75t_R _16606_ (.A1(_00302_),
    .A2(_09191_),
    .B1(_09205_),
    .B2(_09208_),
    .Y(_09209_));
 OA21x2_ASAP7_75t_R _16607_ (.A1(_08733_),
    .A2(_09204_),
    .B(_09209_),
    .Y(_01589_));
 BUFx12_ASAP7_75t_R _16608_ (.A(_08458_),
    .Y(_09210_));
 AOI22x1_ASAP7_75t_R _16609_ (.A1(_00269_),
    .A2(_09191_),
    .B1(_09205_),
    .B2(_09210_),
    .Y(_09211_));
 OA21x2_ASAP7_75t_R _16610_ (.A1(_08735_),
    .A2(_09204_),
    .B(_09211_),
    .Y(_01590_));
 BUFx10_ASAP7_75t_R _16611_ (.A(_08476_),
    .Y(_09212_));
 AOI22x1_ASAP7_75t_R _16612_ (.A1(_00236_),
    .A2(_09191_),
    .B1(_09205_),
    .B2(_09212_),
    .Y(_09213_));
 OA21x2_ASAP7_75t_R _16613_ (.A1(_08737_),
    .A2(_09204_),
    .B(_09213_),
    .Y(_01591_));
 BUFx10_ASAP7_75t_R _16614_ (.A(_08494_),
    .Y(_09214_));
 AOI22x1_ASAP7_75t_R _16615_ (.A1(_00202_),
    .A2(_09191_),
    .B1(_09205_),
    .B2(_09214_),
    .Y(_09215_));
 OA21x2_ASAP7_75t_R _16616_ (.A1(_08739_),
    .A2(_09204_),
    .B(_09215_),
    .Y(_01592_));
 BUFx10_ASAP7_75t_R _16617_ (.A(_08511_),
    .Y(_09216_));
 AOI22x1_ASAP7_75t_R _16618_ (.A1(_00169_),
    .A2(_09191_),
    .B1(_09205_),
    .B2(_09216_),
    .Y(_09217_));
 OA21x2_ASAP7_75t_R _16619_ (.A1(_08741_),
    .A2(_09204_),
    .B(_09217_),
    .Y(_01593_));
 INVx1_ASAP7_75t_R _16620_ (.A(_00135_),
    .Y(_09218_));
 BUFx6f_ASAP7_75t_R _16621_ (.A(_08517_),
    .Y(_09219_));
 OA222x2_ASAP7_75t_R _16622_ (.A1(_09218_),
    .A2(_09168_),
    .B1(_09169_),
    .B2(_08744_),
    .C1(_09171_),
    .C2(_09219_),
    .Y(_01594_));
 BUFx10_ASAP7_75t_R _16623_ (.A(_08545_),
    .Y(_09220_));
 AOI22x1_ASAP7_75t_R _16624_ (.A1(_00102_),
    .A2(_09202_),
    .B1(_09205_),
    .B2(_09220_),
    .Y(_09221_));
 OA21x2_ASAP7_75t_R _16625_ (.A1(_08745_),
    .A2(_09204_),
    .B(_09221_),
    .Y(_01595_));
 NOR2x1_ASAP7_75t_R _16626_ (.A(_01000_),
    .B(_09168_),
    .Y(_09222_));
 AO21x1_ASAP7_75t_R _16627_ (.A1(_08747_),
    .A2(_09168_),
    .B(_09222_),
    .Y(_01596_));
 BUFx6f_ASAP7_75t_R _16628_ (.A(_08564_),
    .Y(_09223_));
 AND3x1_ASAP7_75t_R _16629_ (.A(_08824_),
    .B(_09175_),
    .C(_08873_),
    .Y(_09224_));
 NOR2x1_ASAP7_75t_R _16630_ (.A(_00068_),
    .B(_09168_),
    .Y(_09225_));
 AO221x1_ASAP7_75t_R _16631_ (.A1(_09223_),
    .A2(_09168_),
    .B1(_09224_),
    .B2(_08752_),
    .C(_09225_),
    .Y(_01597_));
 BUFx6f_ASAP7_75t_R _16632_ (.A(_08590_),
    .Y(_09226_));
 AND2x2_ASAP7_75t_R _16633_ (.A(_00036_),
    .B(_09202_),
    .Y(_09227_));
 AOI221x1_ASAP7_75t_R _16634_ (.A1(_09226_),
    .A2(_09224_),
    .B1(_09177_),
    .B2(_08754_),
    .C(_09227_),
    .Y(_01598_));
 BUFx12f_ASAP7_75t_R _16635_ (.A(_08603_),
    .Y(_09228_));
 AOI22x1_ASAP7_75t_R _16636_ (.A1(_00967_),
    .A2(_09202_),
    .B1(_09205_),
    .B2(_09228_),
    .Y(_09229_));
 OA21x2_ASAP7_75t_R _16637_ (.A1(_08756_),
    .A2(_09204_),
    .B(_09229_),
    .Y(_01599_));
 BUFx10_ASAP7_75t_R _16638_ (.A(_08618_),
    .Y(_09230_));
 AO21x1_ASAP7_75t_R _16639_ (.A1(_09175_),
    .A2(_09051_),
    .B(_06478_),
    .Y(_09231_));
 OA221x2_ASAP7_75t_R _16640_ (.A1(_08758_),
    .A2(_09174_),
    .B1(_09169_),
    .B2(_09230_),
    .C(_09231_),
    .Y(_01600_));
 BUFx10_ASAP7_75t_R _16641_ (.A(_08630_),
    .Y(_09232_));
 NAND2x1_ASAP7_75t_R _16642_ (.A(_00900_),
    .B(_09202_),
    .Y(_09233_));
 OA221x2_ASAP7_75t_R _16643_ (.A1(_09232_),
    .A2(_09174_),
    .B1(_09169_),
    .B2(_08760_),
    .C(_09233_),
    .Y(_01601_));
 BUFx12f_ASAP7_75t_R _16644_ (.A(_08643_),
    .Y(_09234_));
 AOI22x1_ASAP7_75t_R _16645_ (.A1(_00867_),
    .A2(_09202_),
    .B1(_09205_),
    .B2(_09234_),
    .Y(_09235_));
 OA21x2_ASAP7_75t_R _16646_ (.A1(_08762_),
    .A2(_09204_),
    .B(_09235_),
    .Y(_01602_));
 NAND2x1_ASAP7_75t_R _16647_ (.A(_00833_),
    .B(_09202_),
    .Y(_09236_));
 OA21x2_ASAP7_75t_R _16648_ (.A1(_08765_),
    .A2(_09202_),
    .B(_09236_),
    .Y(_09237_));
 OA21x2_ASAP7_75t_R _16649_ (.A1(_08764_),
    .A2(_09204_),
    .B(_09237_),
    .Y(_01603_));
 BUFx10_ASAP7_75t_R _16650_ (.A(_08669_),
    .Y(_09238_));
 AOI22x1_ASAP7_75t_R _16651_ (.A1(_00800_),
    .A2(_09202_),
    .B1(_09205_),
    .B2(_09238_),
    .Y(_09239_));
 OA21x2_ASAP7_75t_R _16652_ (.A1(_08768_),
    .A2(_09169_),
    .B(_09239_),
    .Y(_01604_));
 NAND2x1_ASAP7_75t_R _16653_ (.A(_00766_),
    .B(_09173_),
    .Y(_09240_));
 OA21x2_ASAP7_75t_R _16654_ (.A1(_08771_),
    .A2(_09202_),
    .B(_09240_),
    .Y(_09241_));
 OA21x2_ASAP7_75t_R _16655_ (.A1(_08770_),
    .A2(_09169_),
    .B(_09241_),
    .Y(_01605_));
 OR4x2_ASAP7_75t_R _16656_ (.A(_03713_),
    .B(_08099_),
    .C(net2),
    .D(_08100_),
    .Y(_09242_));
 OR3x1_ASAP7_75t_R _16657_ (.A(_08113_),
    .B(_08778_),
    .C(_09242_),
    .Y(_09243_));
 BUFx6f_ASAP7_75t_R _16658_ (.A(_09243_),
    .Y(_09244_));
 BUFx6f_ASAP7_75t_R _16659_ (.A(_09244_),
    .Y(_09245_));
 OR3x4_ASAP7_75t_R _16660_ (.A(_08106_),
    .B(_08778_),
    .C(_09242_),
    .Y(_09246_));
 CKINVDCx6p67_ASAP7_75t_R _16661_ (.A(_09242_),
    .Y(_09247_));
 NAND2x2_ASAP7_75t_R _16662_ (.A(_08787_),
    .B(_09247_),
    .Y(_09248_));
 NAND2x1_ASAP7_75t_R _16663_ (.A(_00020_),
    .B(_09248_),
    .Y(_09249_));
 OA21x2_ASAP7_75t_R _16664_ (.A1(_08111_),
    .A2(_09246_),
    .B(_09249_),
    .Y(_09250_));
 OA21x2_ASAP7_75t_R _16665_ (.A1(_09167_),
    .A2(_09245_),
    .B(_09250_),
    .Y(_01606_));
 BUFx4f_ASAP7_75t_R _16666_ (.A(_08143_),
    .Y(_09251_));
 BUFx12f_ASAP7_75t_R _16667_ (.A(_09248_),
    .Y(_09252_));
 BUFx4f_ASAP7_75t_R _16668_ (.A(_09247_),
    .Y(_09253_));
 AND3x2_ASAP7_75t_R _16669_ (.A(_08798_),
    .B(_08795_),
    .C(_09253_),
    .Y(_09254_));
 BUFx12f_ASAP7_75t_R _16670_ (.A(_09254_),
    .Y(_09255_));
 AOI22x1_ASAP7_75t_R _16671_ (.A1(_00752_),
    .A2(_09252_),
    .B1(_09255_),
    .B2(_09178_),
    .Y(_09256_));
 OA21x2_ASAP7_75t_R _16672_ (.A1(_09251_),
    .A2(_09245_),
    .B(_09256_),
    .Y(_01607_));
 BUFx4f_ASAP7_75t_R _16673_ (.A(_08178_),
    .Y(_09257_));
 AOI22x1_ASAP7_75t_R _16674_ (.A1(_00719_),
    .A2(_09252_),
    .B1(_09255_),
    .B2(_09180_),
    .Y(_09258_));
 OA21x2_ASAP7_75t_R _16675_ (.A1(_09257_),
    .A2(_09245_),
    .B(_09258_),
    .Y(_01608_));
 AND2x6_ASAP7_75t_R _16676_ (.A(_08788_),
    .B(_09253_),
    .Y(_09259_));
 BUFx6f_ASAP7_75t_R _16677_ (.A(_08206_),
    .Y(_09260_));
 OA222x2_ASAP7_75t_R _16678_ (.A1(_05694_),
    .A2(_09259_),
    .B1(_09244_),
    .B2(_09260_),
    .C1(_09246_),
    .C2(_09182_),
    .Y(_01609_));
 BUFx6f_ASAP7_75t_R _16679_ (.A(_08224_),
    .Y(_09261_));
 OA222x2_ASAP7_75t_R _16680_ (.A1(_05631_),
    .A2(_09259_),
    .B1(_09244_),
    .B2(_09261_),
    .C1(_09246_),
    .C2(_09184_),
    .Y(_01610_));
 BUFx4f_ASAP7_75t_R _16681_ (.A(_08240_),
    .Y(_09262_));
 AOI22x1_ASAP7_75t_R _16682_ (.A1(_00620_),
    .A2(_09252_),
    .B1(_09255_),
    .B2(_09185_),
    .Y(_09263_));
 OA21x2_ASAP7_75t_R _16683_ (.A1(_09262_),
    .A2(_09245_),
    .B(_09263_),
    .Y(_01611_));
 BUFx4f_ASAP7_75t_R _16684_ (.A(_08256_),
    .Y(_09264_));
 AOI22x1_ASAP7_75t_R _16685_ (.A1(_00586_),
    .A2(_09252_),
    .B1(_09255_),
    .B2(_09187_),
    .Y(_09265_));
 OA21x2_ASAP7_75t_R _16686_ (.A1(_09264_),
    .A2(_09245_),
    .B(_09265_),
    .Y(_01612_));
 BUFx4f_ASAP7_75t_R _16687_ (.A(_08279_),
    .Y(_09266_));
 AOI22x1_ASAP7_75t_R _16688_ (.A1(_00553_),
    .A2(_09252_),
    .B1(_09255_),
    .B2(_09189_),
    .Y(_09267_));
 OA21x2_ASAP7_75t_R _16689_ (.A1(_09266_),
    .A2(_09245_),
    .B(_09267_),
    .Y(_01613_));
 BUFx4f_ASAP7_75t_R _16690_ (.A(_08301_),
    .Y(_09268_));
 BUFx16f_ASAP7_75t_R _16691_ (.A(_09248_),
    .Y(_09269_));
 AOI22x1_ASAP7_75t_R _16692_ (.A1(_00520_),
    .A2(_09269_),
    .B1(_09255_),
    .B2(_09192_),
    .Y(_09270_));
 OA21x2_ASAP7_75t_R _16693_ (.A1(_09268_),
    .A2(_09245_),
    .B(_09270_),
    .Y(_01614_));
 BUFx4f_ASAP7_75t_R _16694_ (.A(_08323_),
    .Y(_09271_));
 AOI22x1_ASAP7_75t_R _16695_ (.A1(_00487_),
    .A2(_09269_),
    .B1(_09255_),
    .B2(_09194_),
    .Y(_09272_));
 OA21x2_ASAP7_75t_R _16696_ (.A1(_09271_),
    .A2(_09245_),
    .B(_09272_),
    .Y(_01615_));
 BUFx4f_ASAP7_75t_R _16697_ (.A(_08344_),
    .Y(_09273_));
 AOI22x1_ASAP7_75t_R _16698_ (.A1(_00454_),
    .A2(_09269_),
    .B1(_09255_),
    .B2(_09196_),
    .Y(_09274_));
 OA21x2_ASAP7_75t_R _16699_ (.A1(_09273_),
    .A2(_09245_),
    .B(_09274_),
    .Y(_01616_));
 BUFx6f_ASAP7_75t_R _16700_ (.A(_08364_),
    .Y(_09275_));
 NAND2x1_ASAP7_75t_R _16701_ (.A(_01052_),
    .B(_09252_),
    .Y(_09276_));
 OA21x2_ASAP7_75t_R _16702_ (.A1(_09275_),
    .A2(_09252_),
    .B(_09276_),
    .Y(_01617_));
 BUFx4f_ASAP7_75t_R _16703_ (.A(_08378_),
    .Y(_09277_));
 AOI22x1_ASAP7_75t_R _16704_ (.A1(_00421_),
    .A2(_09269_),
    .B1(_09255_),
    .B2(_09199_),
    .Y(_09278_));
 OA21x2_ASAP7_75t_R _16705_ (.A1(_09277_),
    .A2(_09245_),
    .B(_09278_),
    .Y(_01618_));
 BUFx6f_ASAP7_75t_R _16706_ (.A(_08396_),
    .Y(_09279_));
 BUFx10_ASAP7_75t_R _16707_ (.A(_09248_),
    .Y(_09280_));
 NAND2x1_ASAP7_75t_R _16708_ (.A(_00388_),
    .B(_09280_),
    .Y(_09281_));
 OA221x2_ASAP7_75t_R _16709_ (.A1(_09201_),
    .A2(_09252_),
    .B1(_09244_),
    .B2(_09279_),
    .C(_09281_),
    .Y(_01619_));
 BUFx4f_ASAP7_75t_R _16710_ (.A(_08415_),
    .Y(_09282_));
 BUFx6f_ASAP7_75t_R _16711_ (.A(_09244_),
    .Y(_09283_));
 BUFx12_ASAP7_75t_R _16712_ (.A(_09254_),
    .Y(_09284_));
 AOI22x1_ASAP7_75t_R _16713_ (.A1(_00355_),
    .A2(_09269_),
    .B1(_09284_),
    .B2(_09206_),
    .Y(_09285_));
 OA21x2_ASAP7_75t_R _16714_ (.A1(_09282_),
    .A2(_09283_),
    .B(_09285_),
    .Y(_01620_));
 BUFx4f_ASAP7_75t_R _16715_ (.A(_08434_),
    .Y(_09286_));
 AOI22x1_ASAP7_75t_R _16716_ (.A1(_00321_),
    .A2(_09269_),
    .B1(_09284_),
    .B2(_09208_),
    .Y(_09287_));
 OA21x2_ASAP7_75t_R _16717_ (.A1(_09286_),
    .A2(_09283_),
    .B(_09287_),
    .Y(_01621_));
 BUFx6f_ASAP7_75t_R _16718_ (.A(_08455_),
    .Y(_09288_));
 AOI22x1_ASAP7_75t_R _16719_ (.A1(_00288_),
    .A2(_09269_),
    .B1(_09284_),
    .B2(_09210_),
    .Y(_09289_));
 OA21x2_ASAP7_75t_R _16720_ (.A1(_09288_),
    .A2(_09283_),
    .B(_09289_),
    .Y(_01622_));
 BUFx6f_ASAP7_75t_R _16721_ (.A(_08472_),
    .Y(_09290_));
 AOI22x1_ASAP7_75t_R _16722_ (.A1(_00255_),
    .A2(_09269_),
    .B1(_09284_),
    .B2(_09212_),
    .Y(_09291_));
 OA21x2_ASAP7_75t_R _16723_ (.A1(_09290_),
    .A2(_09283_),
    .B(_09291_),
    .Y(_01623_));
 BUFx6f_ASAP7_75t_R _16724_ (.A(_08491_),
    .Y(_09292_));
 AOI22x1_ASAP7_75t_R _16725_ (.A1(_00221_),
    .A2(_09269_),
    .B1(_09284_),
    .B2(_09214_),
    .Y(_09293_));
 OA21x2_ASAP7_75t_R _16726_ (.A1(_09292_),
    .A2(_09283_),
    .B(_09293_),
    .Y(_01624_));
 BUFx6f_ASAP7_75t_R _16727_ (.A(_08508_),
    .Y(_09294_));
 AOI22x1_ASAP7_75t_R _16728_ (.A1(_00188_),
    .A2(_09269_),
    .B1(_09284_),
    .B2(_09216_),
    .Y(_09295_));
 OA21x2_ASAP7_75t_R _16729_ (.A1(_09294_),
    .A2(_09283_),
    .B(_09295_),
    .Y(_01625_));
 BUFx6f_ASAP7_75t_R _16730_ (.A(_08531_),
    .Y(_09296_));
 OA222x2_ASAP7_75t_R _16731_ (.A1(_03974_),
    .A2(_09259_),
    .B1(_09244_),
    .B2(_09296_),
    .C1(_09246_),
    .C2(_09219_),
    .Y(_01626_));
 BUFx6f_ASAP7_75t_R _16732_ (.A(_08542_),
    .Y(_09297_));
 AOI22x1_ASAP7_75t_R _16733_ (.A1(_00121_),
    .A2(_09280_),
    .B1(_09284_),
    .B2(_09220_),
    .Y(_09298_));
 OA21x2_ASAP7_75t_R _16734_ (.A1(_09297_),
    .A2(_09283_),
    .B(_09298_),
    .Y(_01627_));
 BUFx3_ASAP7_75t_R _16735_ (.A(_08560_),
    .Y(_09299_));
 NOR2x1_ASAP7_75t_R _16736_ (.A(_01019_),
    .B(_09259_),
    .Y(_09300_));
 AO21x1_ASAP7_75t_R _16737_ (.A1(_09299_),
    .A2(_09259_),
    .B(_09300_),
    .Y(_01628_));
 AND3x1_ASAP7_75t_R _16738_ (.A(_08824_),
    .B(_08788_),
    .C(_09253_),
    .Y(_09301_));
 BUFx4f_ASAP7_75t_R _16739_ (.A(_08576_),
    .Y(_09302_));
 NOR2x1_ASAP7_75t_R _16740_ (.A(_00087_),
    .B(_09259_),
    .Y(_09303_));
 AO221x1_ASAP7_75t_R _16741_ (.A1(_09223_),
    .A2(_09259_),
    .B1(_09301_),
    .B2(_09302_),
    .C(_09303_),
    .Y(_01629_));
 BUFx6f_ASAP7_75t_R _16742_ (.A(_08594_),
    .Y(_09304_));
 AND2x2_ASAP7_75t_R _16743_ (.A(_00055_),
    .B(_09280_),
    .Y(_09305_));
 AOI221x1_ASAP7_75t_R _16744_ (.A1(_09226_),
    .A2(_09301_),
    .B1(_09255_),
    .B2(_09304_),
    .C(_09305_),
    .Y(_01630_));
 BUFx10_ASAP7_75t_R _16745_ (.A(_08601_),
    .Y(_09306_));
 AOI22x1_ASAP7_75t_R _16746_ (.A1(_00986_),
    .A2(_09280_),
    .B1(_09284_),
    .B2(_09228_),
    .Y(_09307_));
 OA21x2_ASAP7_75t_R _16747_ (.A1(_09306_),
    .A2(_09283_),
    .B(_09307_),
    .Y(_01631_));
 BUFx6f_ASAP7_75t_R _16748_ (.A(_08609_),
    .Y(_09308_));
 NAND2x1_ASAP7_75t_R _16749_ (.A(_00953_),
    .B(_09280_),
    .Y(_09309_));
 OA221x2_ASAP7_75t_R _16750_ (.A1(_09308_),
    .A2(_09252_),
    .B1(_09244_),
    .B2(_09230_),
    .C(_09309_),
    .Y(_01632_));
 BUFx6f_ASAP7_75t_R _16751_ (.A(_08628_),
    .Y(_09310_));
 NAND2x1_ASAP7_75t_R _16752_ (.A(_00919_),
    .B(_09280_),
    .Y(_09311_));
 OA221x2_ASAP7_75t_R _16753_ (.A1(_09232_),
    .A2(_09252_),
    .B1(_09244_),
    .B2(_09310_),
    .C(_09311_),
    .Y(_01633_));
 BUFx10_ASAP7_75t_R _16754_ (.A(_08641_),
    .Y(_09312_));
 AOI22x1_ASAP7_75t_R _16755_ (.A1(_00886_),
    .A2(_09280_),
    .B1(_09284_),
    .B2(_09234_),
    .Y(_09313_));
 OA21x2_ASAP7_75t_R _16756_ (.A1(_09312_),
    .A2(_09283_),
    .B(_09313_),
    .Y(_01634_));
 BUFx6f_ASAP7_75t_R _16757_ (.A(_08654_),
    .Y(_09314_));
 BUFx6f_ASAP7_75t_R _16758_ (.A(_08656_),
    .Y(_09315_));
 NAND2x1_ASAP7_75t_R _16759_ (.A(_00852_),
    .B(_09248_),
    .Y(_09316_));
 OA21x2_ASAP7_75t_R _16760_ (.A1(_09315_),
    .A2(_09280_),
    .B(_09316_),
    .Y(_09317_));
 OA21x2_ASAP7_75t_R _16761_ (.A1(_09314_),
    .A2(_09283_),
    .B(_09317_),
    .Y(_01635_));
 BUFx4f_ASAP7_75t_R _16762_ (.A(_08667_),
    .Y(_09318_));
 AOI22x1_ASAP7_75t_R _16763_ (.A1(_00819_),
    .A2(_09280_),
    .B1(_09284_),
    .B2(_09238_),
    .Y(_09319_));
 OA21x2_ASAP7_75t_R _16764_ (.A1(_09318_),
    .A2(_09244_),
    .B(_09319_),
    .Y(_01636_));
 BUFx6f_ASAP7_75t_R _16765_ (.A(_08680_),
    .Y(_09320_));
 BUFx6f_ASAP7_75t_R _16766_ (.A(_08684_),
    .Y(_09321_));
 NAND2x1_ASAP7_75t_R _16767_ (.A(_00785_),
    .B(_09248_),
    .Y(_09322_));
 OA21x2_ASAP7_75t_R _16768_ (.A1(_09321_),
    .A2(_09280_),
    .B(_09322_),
    .Y(_09323_));
 OA21x2_ASAP7_75t_R _16769_ (.A1(_09320_),
    .A2(_09244_),
    .B(_09323_),
    .Y(_01637_));
 BUFx16f_ASAP7_75t_R _16770_ (.A(_08105_),
    .Y(_09324_));
 AND2x6_ASAP7_75t_R _16771_ (.A(_08837_),
    .B(_09247_),
    .Y(_09325_));
 NAND2x2_ASAP7_75t_R _16772_ (.A(_09324_),
    .B(_09325_),
    .Y(_09326_));
 BUFx6f_ASAP7_75t_R _16773_ (.A(_09326_),
    .Y(_09327_));
 INVx1_ASAP7_75t_R _16774_ (.A(_00021_),
    .Y(_09328_));
 NAND2x2_ASAP7_75t_R _16775_ (.A(_08937_),
    .B(_09325_),
    .Y(_09329_));
 BUFx6f_ASAP7_75t_R _16776_ (.A(_08110_),
    .Y(_09330_));
 OA22x2_ASAP7_75t_R _16777_ (.A1(_09328_),
    .A2(_09325_),
    .B1(_09329_),
    .B2(_09330_),
    .Y(_09331_));
 OA21x2_ASAP7_75t_R _16778_ (.A1(_09167_),
    .A2(_09327_),
    .B(_09331_),
    .Y(_01638_));
 NAND2x2_ASAP7_75t_R _16779_ (.A(_08847_),
    .B(_09253_),
    .Y(_09332_));
 BUFx12f_ASAP7_75t_R _16780_ (.A(_09332_),
    .Y(_09333_));
 AND3x2_ASAP7_75t_R _16781_ (.A(_08798_),
    .B(_08847_),
    .C(_09253_),
    .Y(_09334_));
 BUFx12f_ASAP7_75t_R _16782_ (.A(_09334_),
    .Y(_09335_));
 AOI22x1_ASAP7_75t_R _16783_ (.A1(_00753_),
    .A2(_09333_),
    .B1(_09335_),
    .B2(_09178_),
    .Y(_09336_));
 OA21x2_ASAP7_75t_R _16784_ (.A1(_09251_),
    .A2(_09327_),
    .B(_09336_),
    .Y(_01639_));
 AOI22x1_ASAP7_75t_R _16785_ (.A1(_00720_),
    .A2(_09333_),
    .B1(_09335_),
    .B2(_09180_),
    .Y(_09337_));
 OA21x2_ASAP7_75t_R _16786_ (.A1(_09257_),
    .A2(_09327_),
    .B(_09337_),
    .Y(_01640_));
 OA222x2_ASAP7_75t_R _16787_ (.A1(_05692_),
    .A2(_09325_),
    .B1(_09326_),
    .B2(_09260_),
    .C1(_09329_),
    .C2(_09182_),
    .Y(_01641_));
 OA222x2_ASAP7_75t_R _16788_ (.A1(_05632_),
    .A2(_09325_),
    .B1(_09326_),
    .B2(_09261_),
    .C1(_09329_),
    .C2(_09184_),
    .Y(_01642_));
 AOI22x1_ASAP7_75t_R _16789_ (.A1(_00621_),
    .A2(_09333_),
    .B1(_09335_),
    .B2(_09185_),
    .Y(_09338_));
 OA21x2_ASAP7_75t_R _16790_ (.A1(_09262_),
    .A2(_09327_),
    .B(_09338_),
    .Y(_01643_));
 AOI22x1_ASAP7_75t_R _16791_ (.A1(_00587_),
    .A2(_09333_),
    .B1(_09335_),
    .B2(_09187_),
    .Y(_09339_));
 OA21x2_ASAP7_75t_R _16792_ (.A1(_09264_),
    .A2(_09327_),
    .B(_09339_),
    .Y(_01644_));
 AOI22x1_ASAP7_75t_R _16793_ (.A1(_00554_),
    .A2(_09333_),
    .B1(_09335_),
    .B2(_09189_),
    .Y(_09340_));
 OA21x2_ASAP7_75t_R _16794_ (.A1(_09266_),
    .A2(_09327_),
    .B(_09340_),
    .Y(_01645_));
 BUFx16f_ASAP7_75t_R _16795_ (.A(_09332_),
    .Y(_09341_));
 AOI22x1_ASAP7_75t_R _16796_ (.A1(_00521_),
    .A2(_09341_),
    .B1(_09335_),
    .B2(_09192_),
    .Y(_09342_));
 OA21x2_ASAP7_75t_R _16797_ (.A1(_09268_),
    .A2(_09327_),
    .B(_09342_),
    .Y(_01646_));
 AOI22x1_ASAP7_75t_R _16798_ (.A1(_00488_),
    .A2(_09341_),
    .B1(_09335_),
    .B2(_09194_),
    .Y(_09343_));
 OA21x2_ASAP7_75t_R _16799_ (.A1(_09271_),
    .A2(_09327_),
    .B(_09343_),
    .Y(_01647_));
 AOI22x1_ASAP7_75t_R _16800_ (.A1(_00455_),
    .A2(_09341_),
    .B1(_09335_),
    .B2(_09196_),
    .Y(_09344_));
 OA21x2_ASAP7_75t_R _16801_ (.A1(_09273_),
    .A2(_09327_),
    .B(_09344_),
    .Y(_01648_));
 NAND2x1_ASAP7_75t_R _16802_ (.A(_01053_),
    .B(_09333_),
    .Y(_09345_));
 OA21x2_ASAP7_75t_R _16803_ (.A1(_09275_),
    .A2(_09333_),
    .B(_09345_),
    .Y(_01649_));
 AOI22x1_ASAP7_75t_R _16804_ (.A1(_00422_),
    .A2(_09341_),
    .B1(_09335_),
    .B2(_09199_),
    .Y(_09346_));
 OA21x2_ASAP7_75t_R _16805_ (.A1(_09277_),
    .A2(_09327_),
    .B(_09346_),
    .Y(_01650_));
 BUFx10_ASAP7_75t_R _16806_ (.A(_09332_),
    .Y(_09347_));
 NAND2x1_ASAP7_75t_R _16807_ (.A(_00389_),
    .B(_09347_),
    .Y(_09348_));
 OA221x2_ASAP7_75t_R _16808_ (.A1(_09201_),
    .A2(_09333_),
    .B1(_09326_),
    .B2(_09279_),
    .C(_09348_),
    .Y(_01651_));
 BUFx4f_ASAP7_75t_R _16809_ (.A(_09326_),
    .Y(_09349_));
 BUFx10_ASAP7_75t_R _16810_ (.A(_09334_),
    .Y(_09350_));
 AOI22x1_ASAP7_75t_R _16811_ (.A1(_00356_),
    .A2(_09341_),
    .B1(_09350_),
    .B2(_09206_),
    .Y(_09351_));
 OA21x2_ASAP7_75t_R _16812_ (.A1(_09282_),
    .A2(_09349_),
    .B(_09351_),
    .Y(_01652_));
 AOI22x1_ASAP7_75t_R _16813_ (.A1(_00322_),
    .A2(_09341_),
    .B1(_09350_),
    .B2(_09208_),
    .Y(_09352_));
 OA21x2_ASAP7_75t_R _16814_ (.A1(_09286_),
    .A2(_09349_),
    .B(_09352_),
    .Y(_01653_));
 AOI22x1_ASAP7_75t_R _16815_ (.A1(_00289_),
    .A2(_09341_),
    .B1(_09350_),
    .B2(_09210_),
    .Y(_09353_));
 OA21x2_ASAP7_75t_R _16816_ (.A1(_09288_),
    .A2(_09349_),
    .B(_09353_),
    .Y(_01654_));
 AOI22x1_ASAP7_75t_R _16817_ (.A1(_00256_),
    .A2(_09341_),
    .B1(_09350_),
    .B2(_09212_),
    .Y(_09354_));
 OA21x2_ASAP7_75t_R _16818_ (.A1(_09290_),
    .A2(_09349_),
    .B(_09354_),
    .Y(_01655_));
 AOI22x1_ASAP7_75t_R _16819_ (.A1(_00222_),
    .A2(_09341_),
    .B1(_09350_),
    .B2(_09214_),
    .Y(_09355_));
 OA21x2_ASAP7_75t_R _16820_ (.A1(_09292_),
    .A2(_09349_),
    .B(_09355_),
    .Y(_01656_));
 AOI22x1_ASAP7_75t_R _16821_ (.A1(_00189_),
    .A2(_09341_),
    .B1(_09350_),
    .B2(_09216_),
    .Y(_09356_));
 OA21x2_ASAP7_75t_R _16822_ (.A1(_09294_),
    .A2(_09349_),
    .B(_09356_),
    .Y(_01657_));
 OA222x2_ASAP7_75t_R _16823_ (.A1(_03977_),
    .A2(_09325_),
    .B1(_09326_),
    .B2(_09296_),
    .C1(_09329_),
    .C2(_09219_),
    .Y(_01658_));
 AOI22x1_ASAP7_75t_R _16824_ (.A1(_00122_),
    .A2(_09347_),
    .B1(_09350_),
    .B2(_09220_),
    .Y(_09357_));
 OA21x2_ASAP7_75t_R _16825_ (.A1(_09297_),
    .A2(_09349_),
    .B(_09357_),
    .Y(_01659_));
 NOR2x1_ASAP7_75t_R _16826_ (.A(_01020_),
    .B(_09325_),
    .Y(_09358_));
 AO21x1_ASAP7_75t_R _16827_ (.A1(_09299_),
    .A2(_09325_),
    .B(_09358_),
    .Y(_01660_));
 AND3x1_ASAP7_75t_R _16828_ (.A(_08824_),
    .B(_09051_),
    .C(_09253_),
    .Y(_09359_));
 NOR2x1_ASAP7_75t_R _16829_ (.A(_00088_),
    .B(_09325_),
    .Y(_09360_));
 AO221x1_ASAP7_75t_R _16830_ (.A1(_09223_),
    .A2(_09325_),
    .B1(_09359_),
    .B2(_09302_),
    .C(_09360_),
    .Y(_01661_));
 AND2x2_ASAP7_75t_R _16831_ (.A(_00056_),
    .B(_09347_),
    .Y(_09361_));
 AOI221x1_ASAP7_75t_R _16832_ (.A1(_09226_),
    .A2(_09359_),
    .B1(_09335_),
    .B2(_09304_),
    .C(_09361_),
    .Y(_01662_));
 AOI22x1_ASAP7_75t_R _16833_ (.A1(_00987_),
    .A2(_09347_),
    .B1(_09350_),
    .B2(_09228_),
    .Y(_09362_));
 OA21x2_ASAP7_75t_R _16834_ (.A1(_09306_),
    .A2(_09349_),
    .B(_09362_),
    .Y(_01663_));
 NAND2x1_ASAP7_75t_R _16835_ (.A(_00954_),
    .B(_09347_),
    .Y(_09363_));
 OA221x2_ASAP7_75t_R _16836_ (.A1(_09308_),
    .A2(_09333_),
    .B1(_09326_),
    .B2(_09230_),
    .C(_09363_),
    .Y(_01664_));
 NAND2x1_ASAP7_75t_R _16837_ (.A(_00920_),
    .B(_09347_),
    .Y(_09364_));
 OA221x2_ASAP7_75t_R _16838_ (.A1(_09232_),
    .A2(_09333_),
    .B1(_09326_),
    .B2(_09310_),
    .C(_09364_),
    .Y(_01665_));
 AOI22x1_ASAP7_75t_R _16839_ (.A1(_00887_),
    .A2(_09347_),
    .B1(_09350_),
    .B2(_09234_),
    .Y(_09365_));
 OA21x2_ASAP7_75t_R _16840_ (.A1(_09312_),
    .A2(_09349_),
    .B(_09365_),
    .Y(_01666_));
 NAND2x1_ASAP7_75t_R _16841_ (.A(_00853_),
    .B(_09332_),
    .Y(_09366_));
 OA21x2_ASAP7_75t_R _16842_ (.A1(_09315_),
    .A2(_09347_),
    .B(_09366_),
    .Y(_09367_));
 OA21x2_ASAP7_75t_R _16843_ (.A1(_09314_),
    .A2(_09349_),
    .B(_09367_),
    .Y(_01667_));
 AOI22x1_ASAP7_75t_R _16844_ (.A1(_00820_),
    .A2(_09347_),
    .B1(_09350_),
    .B2(_09238_),
    .Y(_09368_));
 OA21x2_ASAP7_75t_R _16845_ (.A1(_09318_),
    .A2(_09326_),
    .B(_09368_),
    .Y(_01668_));
 NAND2x1_ASAP7_75t_R _16846_ (.A(_00786_),
    .B(_09332_),
    .Y(_09369_));
 OA21x2_ASAP7_75t_R _16847_ (.A1(_09321_),
    .A2(_09347_),
    .B(_09369_),
    .Y(_09370_));
 OA21x2_ASAP7_75t_R _16848_ (.A1(_09320_),
    .A2(_09326_),
    .B(_09370_),
    .Y(_01669_));
 AND2x6_ASAP7_75t_R _16849_ (.A(_08098_),
    .B(_09247_),
    .Y(_09371_));
 NAND2x2_ASAP7_75t_R _16850_ (.A(_09324_),
    .B(_09371_),
    .Y(_09372_));
 BUFx10_ASAP7_75t_R _16851_ (.A(_09372_),
    .Y(_09373_));
 NAND2x2_ASAP7_75t_R _16852_ (.A(_08115_),
    .B(_09371_),
    .Y(_09374_));
 NAND2x2_ASAP7_75t_R _16853_ (.A(_08117_),
    .B(_09247_),
    .Y(_09375_));
 NAND2x1_ASAP7_75t_R _16854_ (.A(_00022_),
    .B(_09375_),
    .Y(_09376_));
 OA21x2_ASAP7_75t_R _16855_ (.A1(_08111_),
    .A2(_09374_),
    .B(_09376_),
    .Y(_09377_));
 OA21x2_ASAP7_75t_R _16856_ (.A1(_09167_),
    .A2(_09373_),
    .B(_09377_),
    .Y(_01670_));
 BUFx12f_ASAP7_75t_R _16857_ (.A(_09375_),
    .Y(_09378_));
 AND3x2_ASAP7_75t_R _16858_ (.A(_08117_),
    .B(_08701_),
    .C(_09253_),
    .Y(_09379_));
 BUFx12f_ASAP7_75t_R _16859_ (.A(_09379_),
    .Y(_09380_));
 AOI22x1_ASAP7_75t_R _16860_ (.A1(_00754_),
    .A2(_09378_),
    .B1(_09380_),
    .B2(_09178_),
    .Y(_09381_));
 OA21x2_ASAP7_75t_R _16861_ (.A1(_09251_),
    .A2(_09373_),
    .B(_09381_),
    .Y(_01671_));
 AOI22x1_ASAP7_75t_R _16862_ (.A1(_00721_),
    .A2(_09378_),
    .B1(_09380_),
    .B2(_09180_),
    .Y(_09382_));
 OA21x2_ASAP7_75t_R _16863_ (.A1(_09257_),
    .A2(_09373_),
    .B(_09382_),
    .Y(_01672_));
 OA222x2_ASAP7_75t_R _16864_ (.A1(_05688_),
    .A2(_09371_),
    .B1(_09372_),
    .B2(_09260_),
    .C1(_09374_),
    .C2(_09182_),
    .Y(_01673_));
 INVx1_ASAP7_75t_R _16865_ (.A(_00655_),
    .Y(_09383_));
 OA222x2_ASAP7_75t_R _16866_ (.A1(_09383_),
    .A2(_09371_),
    .B1(_09372_),
    .B2(_09261_),
    .C1(_09374_),
    .C2(_09184_),
    .Y(_01674_));
 AOI22x1_ASAP7_75t_R _16867_ (.A1(_00622_),
    .A2(_09378_),
    .B1(_09380_),
    .B2(_09185_),
    .Y(_09384_));
 OA21x2_ASAP7_75t_R _16868_ (.A1(_09262_),
    .A2(_09373_),
    .B(_09384_),
    .Y(_01675_));
 AOI22x1_ASAP7_75t_R _16869_ (.A1(_00588_),
    .A2(_09378_),
    .B1(_09380_),
    .B2(_09187_),
    .Y(_09385_));
 OA21x2_ASAP7_75t_R _16870_ (.A1(_09264_),
    .A2(_09373_),
    .B(_09385_),
    .Y(_01676_));
 AOI22x1_ASAP7_75t_R _16871_ (.A1(_00555_),
    .A2(_09378_),
    .B1(_09380_),
    .B2(_09189_),
    .Y(_09386_));
 OA21x2_ASAP7_75t_R _16872_ (.A1(_09266_),
    .A2(_09373_),
    .B(_09386_),
    .Y(_01677_));
 BUFx16f_ASAP7_75t_R _16873_ (.A(_09375_),
    .Y(_09387_));
 AOI22x1_ASAP7_75t_R _16874_ (.A1(_00522_),
    .A2(_09387_),
    .B1(_09380_),
    .B2(_09192_),
    .Y(_09388_));
 OA21x2_ASAP7_75t_R _16875_ (.A1(_09268_),
    .A2(_09373_),
    .B(_09388_),
    .Y(_01678_));
 AOI22x1_ASAP7_75t_R _16876_ (.A1(_00489_),
    .A2(_09387_),
    .B1(_09380_),
    .B2(_09194_),
    .Y(_09389_));
 OA21x2_ASAP7_75t_R _16877_ (.A1(_09271_),
    .A2(_09373_),
    .B(_09389_),
    .Y(_01679_));
 AOI22x1_ASAP7_75t_R _16878_ (.A1(_00456_),
    .A2(_09387_),
    .B1(_09380_),
    .B2(_09196_),
    .Y(_09390_));
 OA21x2_ASAP7_75t_R _16879_ (.A1(_09273_),
    .A2(_09373_),
    .B(_09390_),
    .Y(_01680_));
 NAND2x1_ASAP7_75t_R _16880_ (.A(_01054_),
    .B(_09378_),
    .Y(_09391_));
 OA21x2_ASAP7_75t_R _16881_ (.A1(_09275_),
    .A2(_09378_),
    .B(_09391_),
    .Y(_01681_));
 AOI22x1_ASAP7_75t_R _16882_ (.A1(_00423_),
    .A2(_09387_),
    .B1(_09380_),
    .B2(_09199_),
    .Y(_09392_));
 OA21x2_ASAP7_75t_R _16883_ (.A1(_09277_),
    .A2(_09373_),
    .B(_09392_),
    .Y(_01682_));
 BUFx10_ASAP7_75t_R _16884_ (.A(_09375_),
    .Y(_09393_));
 NAND2x1_ASAP7_75t_R _16885_ (.A(_00390_),
    .B(_09393_),
    .Y(_09394_));
 OA221x2_ASAP7_75t_R _16886_ (.A1(_09201_),
    .A2(_09378_),
    .B1(_09372_),
    .B2(_09279_),
    .C(_09394_),
    .Y(_01683_));
 BUFx4f_ASAP7_75t_R _16887_ (.A(_09372_),
    .Y(_09395_));
 BUFx10_ASAP7_75t_R _16888_ (.A(_09379_),
    .Y(_09396_));
 AOI22x1_ASAP7_75t_R _16889_ (.A1(_00357_),
    .A2(_09387_),
    .B1(_09396_),
    .B2(_09206_),
    .Y(_09397_));
 OA21x2_ASAP7_75t_R _16890_ (.A1(_09282_),
    .A2(_09395_),
    .B(_09397_),
    .Y(_01684_));
 AOI22x1_ASAP7_75t_R _16891_ (.A1(_00323_),
    .A2(_09387_),
    .B1(_09396_),
    .B2(_09208_),
    .Y(_09398_));
 OA21x2_ASAP7_75t_R _16892_ (.A1(_09286_),
    .A2(_09395_),
    .B(_09398_),
    .Y(_01685_));
 AOI22x1_ASAP7_75t_R _16893_ (.A1(_00290_),
    .A2(_09387_),
    .B1(_09396_),
    .B2(_09210_),
    .Y(_09399_));
 OA21x2_ASAP7_75t_R _16894_ (.A1(_09288_),
    .A2(_09395_),
    .B(_09399_),
    .Y(_01686_));
 AOI22x1_ASAP7_75t_R _16895_ (.A1(_00257_),
    .A2(_09387_),
    .B1(_09396_),
    .B2(_09212_),
    .Y(_09400_));
 OA21x2_ASAP7_75t_R _16896_ (.A1(_09290_),
    .A2(_09395_),
    .B(_09400_),
    .Y(_01687_));
 AOI22x1_ASAP7_75t_R _16897_ (.A1(_00223_),
    .A2(_09387_),
    .B1(_09396_),
    .B2(_09214_),
    .Y(_09401_));
 OA21x2_ASAP7_75t_R _16898_ (.A1(_09292_),
    .A2(_09395_),
    .B(_09401_),
    .Y(_01688_));
 AOI22x1_ASAP7_75t_R _16899_ (.A1(_00190_),
    .A2(_09387_),
    .B1(_09396_),
    .B2(_09216_),
    .Y(_09402_));
 OA21x2_ASAP7_75t_R _16900_ (.A1(_09294_),
    .A2(_09395_),
    .B(_09402_),
    .Y(_01689_));
 INVx1_ASAP7_75t_R _16901_ (.A(_00156_),
    .Y(_09403_));
 OA222x2_ASAP7_75t_R _16902_ (.A1(_09403_),
    .A2(_09371_),
    .B1(_09372_),
    .B2(_09296_),
    .C1(_09374_),
    .C2(_09219_),
    .Y(_01690_));
 AOI22x1_ASAP7_75t_R _16903_ (.A1(_00123_),
    .A2(_09393_),
    .B1(_09396_),
    .B2(_09220_),
    .Y(_09404_));
 OA21x2_ASAP7_75t_R _16904_ (.A1(_09297_),
    .A2(_09395_),
    .B(_09404_),
    .Y(_01691_));
 NOR2x1_ASAP7_75t_R _16905_ (.A(_01021_),
    .B(_09371_),
    .Y(_09405_));
 AO21x1_ASAP7_75t_R _16906_ (.A1(_09299_),
    .A2(_09371_),
    .B(_09405_),
    .Y(_01692_));
 AND3x2_ASAP7_75t_R _16907_ (.A(_08145_),
    .B(_08577_),
    .C(_09253_),
    .Y(_09406_));
 NOR2x1_ASAP7_75t_R _16908_ (.A(_00089_),
    .B(_09371_),
    .Y(_09407_));
 AO221x1_ASAP7_75t_R _16909_ (.A1(_09223_),
    .A2(_09371_),
    .B1(_09406_),
    .B2(_09302_),
    .C(_09407_),
    .Y(_01693_));
 AND2x2_ASAP7_75t_R _16910_ (.A(_00057_),
    .B(_09393_),
    .Y(_09408_));
 AOI221x1_ASAP7_75t_R _16911_ (.A1(_09226_),
    .A2(_09406_),
    .B1(_09380_),
    .B2(_09304_),
    .C(_09408_),
    .Y(_01694_));
 AOI22x1_ASAP7_75t_R _16912_ (.A1(_00988_),
    .A2(_09393_),
    .B1(_09396_),
    .B2(_09228_),
    .Y(_09409_));
 OA21x2_ASAP7_75t_R _16913_ (.A1(_09306_),
    .A2(_09395_),
    .B(_09409_),
    .Y(_01695_));
 NAND2x1_ASAP7_75t_R _16914_ (.A(_00955_),
    .B(_09393_),
    .Y(_09410_));
 OA221x2_ASAP7_75t_R _16915_ (.A1(_09308_),
    .A2(_09378_),
    .B1(_09372_),
    .B2(_09230_),
    .C(_09410_),
    .Y(_01696_));
 NAND2x1_ASAP7_75t_R _16916_ (.A(_00921_),
    .B(_09393_),
    .Y(_09411_));
 OA221x2_ASAP7_75t_R _16917_ (.A1(_09232_),
    .A2(_09378_),
    .B1(_09372_),
    .B2(_09310_),
    .C(_09411_),
    .Y(_01697_));
 AOI22x1_ASAP7_75t_R _16918_ (.A1(_00888_),
    .A2(_09393_),
    .B1(_09396_),
    .B2(_09234_),
    .Y(_09412_));
 OA21x2_ASAP7_75t_R _16919_ (.A1(_09312_),
    .A2(_09395_),
    .B(_09412_),
    .Y(_01698_));
 NAND2x1_ASAP7_75t_R _16920_ (.A(_00854_),
    .B(_09375_),
    .Y(_09413_));
 OA21x2_ASAP7_75t_R _16921_ (.A1(_09315_),
    .A2(_09393_),
    .B(_09413_),
    .Y(_09414_));
 OA21x2_ASAP7_75t_R _16922_ (.A1(_09314_),
    .A2(_09395_),
    .B(_09414_),
    .Y(_01699_));
 AOI22x1_ASAP7_75t_R _16923_ (.A1(_00821_),
    .A2(_09393_),
    .B1(_09396_),
    .B2(_09238_),
    .Y(_09415_));
 OA21x2_ASAP7_75t_R _16924_ (.A1(_09318_),
    .A2(_09372_),
    .B(_09415_),
    .Y(_01700_));
 NAND2x1_ASAP7_75t_R _16925_ (.A(_00787_),
    .B(_09375_),
    .Y(_09416_));
 OA21x2_ASAP7_75t_R _16926_ (.A1(_09321_),
    .A2(_09393_),
    .B(_09416_),
    .Y(_09417_));
 OA21x2_ASAP7_75t_R _16927_ (.A1(_09320_),
    .A2(_09372_),
    .B(_09417_),
    .Y(_01701_));
 AND2x6_ASAP7_75t_R _16928_ (.A(_08689_),
    .B(_09247_),
    .Y(_09418_));
 NAND2x2_ASAP7_75t_R _16929_ (.A(_09324_),
    .B(_09418_),
    .Y(_09419_));
 BUFx10_ASAP7_75t_R _16930_ (.A(_09419_),
    .Y(_09420_));
 NAND2x2_ASAP7_75t_R _16931_ (.A(_08937_),
    .B(_09418_),
    .Y(_09421_));
 OA22x2_ASAP7_75t_R _16932_ (.A1(_03030_),
    .A2(_09418_),
    .B1(_09421_),
    .B2(_09330_),
    .Y(_09422_));
 OA21x2_ASAP7_75t_R _16933_ (.A1(_09167_),
    .A2(_09420_),
    .B(_09422_),
    .Y(_01702_));
 NAND2x2_ASAP7_75t_R _16934_ (.A(_08694_),
    .B(_09247_),
    .Y(_09423_));
 BUFx12f_ASAP7_75t_R _16935_ (.A(_09423_),
    .Y(_09424_));
 BUFx4f_ASAP7_75t_R _16936_ (.A(_08113_),
    .Y(_09425_));
 AND3x2_ASAP7_75t_R _16937_ (.A(_09425_),
    .B(_08749_),
    .C(_09253_),
    .Y(_09426_));
 BUFx12f_ASAP7_75t_R _16938_ (.A(_09426_),
    .Y(_09427_));
 AOI22x1_ASAP7_75t_R _16939_ (.A1(_00755_),
    .A2(_09424_),
    .B1(_09427_),
    .B2(_09178_),
    .Y(_09428_));
 OA21x2_ASAP7_75t_R _16940_ (.A1(_09251_),
    .A2(_09420_),
    .B(_09428_),
    .Y(_01703_));
 AOI22x1_ASAP7_75t_R _16941_ (.A1(_00722_),
    .A2(_09424_),
    .B1(_09427_),
    .B2(_09180_),
    .Y(_09429_));
 OA21x2_ASAP7_75t_R _16942_ (.A1(_09257_),
    .A2(_09420_),
    .B(_09429_),
    .Y(_01704_));
 INVx1_ASAP7_75t_R _16943_ (.A(_00689_),
    .Y(_09430_));
 OA222x2_ASAP7_75t_R _16944_ (.A1(_09430_),
    .A2(_09418_),
    .B1(_09419_),
    .B2(_09260_),
    .C1(_09421_),
    .C2(_09182_),
    .Y(_01705_));
 INVx1_ASAP7_75t_R _16945_ (.A(_00656_),
    .Y(_09431_));
 OA222x2_ASAP7_75t_R _16946_ (.A1(_09431_),
    .A2(_09418_),
    .B1(_09419_),
    .B2(_09261_),
    .C1(_09421_),
    .C2(_09184_),
    .Y(_01706_));
 AOI22x1_ASAP7_75t_R _16947_ (.A1(_00623_),
    .A2(_09424_),
    .B1(_09427_),
    .B2(_09185_),
    .Y(_09432_));
 OA21x2_ASAP7_75t_R _16948_ (.A1(_09262_),
    .A2(_09420_),
    .B(_09432_),
    .Y(_01707_));
 AOI22x1_ASAP7_75t_R _16949_ (.A1(_00589_),
    .A2(_09424_),
    .B1(_09427_),
    .B2(_09187_),
    .Y(_09433_));
 OA21x2_ASAP7_75t_R _16950_ (.A1(_09264_),
    .A2(_09420_),
    .B(_09433_),
    .Y(_01708_));
 AOI22x1_ASAP7_75t_R _16951_ (.A1(_00556_),
    .A2(_09424_),
    .B1(_09427_),
    .B2(_09189_),
    .Y(_09434_));
 OA21x2_ASAP7_75t_R _16952_ (.A1(_09266_),
    .A2(_09420_),
    .B(_09434_),
    .Y(_01709_));
 BUFx16f_ASAP7_75t_R _16953_ (.A(_09423_),
    .Y(_09435_));
 AOI22x1_ASAP7_75t_R _16954_ (.A1(_00523_),
    .A2(_09435_),
    .B1(_09427_),
    .B2(_09192_),
    .Y(_09436_));
 OA21x2_ASAP7_75t_R _16955_ (.A1(_09268_),
    .A2(_09420_),
    .B(_09436_),
    .Y(_01710_));
 AOI22x1_ASAP7_75t_R _16956_ (.A1(_00490_),
    .A2(_09435_),
    .B1(_09427_),
    .B2(_09194_),
    .Y(_09437_));
 OA21x2_ASAP7_75t_R _16957_ (.A1(_09271_),
    .A2(_09420_),
    .B(_09437_),
    .Y(_01711_));
 AOI22x1_ASAP7_75t_R _16958_ (.A1(_00457_),
    .A2(_09435_),
    .B1(_09427_),
    .B2(_09196_),
    .Y(_09438_));
 OA21x2_ASAP7_75t_R _16959_ (.A1(_09273_),
    .A2(_09420_),
    .B(_09438_),
    .Y(_01712_));
 NAND2x1_ASAP7_75t_R _16960_ (.A(_01055_),
    .B(_09424_),
    .Y(_09439_));
 OA21x2_ASAP7_75t_R _16961_ (.A1(_09275_),
    .A2(_09424_),
    .B(_09439_),
    .Y(_01713_));
 AOI22x1_ASAP7_75t_R _16962_ (.A1(_00424_),
    .A2(_09435_),
    .B1(_09427_),
    .B2(_09199_),
    .Y(_09440_));
 OA21x2_ASAP7_75t_R _16963_ (.A1(_09277_),
    .A2(_09420_),
    .B(_09440_),
    .Y(_01714_));
 BUFx12_ASAP7_75t_R _16964_ (.A(_09423_),
    .Y(_09441_));
 NAND2x1_ASAP7_75t_R _16965_ (.A(_00391_),
    .B(_09441_),
    .Y(_09442_));
 OA221x2_ASAP7_75t_R _16966_ (.A1(_09201_),
    .A2(_09424_),
    .B1(_09419_),
    .B2(_09279_),
    .C(_09442_),
    .Y(_01715_));
 BUFx6f_ASAP7_75t_R _16967_ (.A(_09419_),
    .Y(_09443_));
 BUFx12_ASAP7_75t_R _16968_ (.A(_09426_),
    .Y(_09444_));
 AOI22x1_ASAP7_75t_R _16969_ (.A1(_00358_),
    .A2(_09435_),
    .B1(_09444_),
    .B2(_09206_),
    .Y(_09445_));
 OA21x2_ASAP7_75t_R _16970_ (.A1(_09282_),
    .A2(_09443_),
    .B(_09445_),
    .Y(_01716_));
 AOI22x1_ASAP7_75t_R _16971_ (.A1(_00324_),
    .A2(_09435_),
    .B1(_09444_),
    .B2(_09208_),
    .Y(_09446_));
 OA21x2_ASAP7_75t_R _16972_ (.A1(_09286_),
    .A2(_09443_),
    .B(_09446_),
    .Y(_01717_));
 AOI22x1_ASAP7_75t_R _16973_ (.A1(_00291_),
    .A2(_09435_),
    .B1(_09444_),
    .B2(_09210_),
    .Y(_09447_));
 OA21x2_ASAP7_75t_R _16974_ (.A1(_09288_),
    .A2(_09443_),
    .B(_09447_),
    .Y(_01718_));
 AOI22x1_ASAP7_75t_R _16975_ (.A1(_00258_),
    .A2(_09435_),
    .B1(_09444_),
    .B2(_09212_),
    .Y(_09448_));
 OA21x2_ASAP7_75t_R _16976_ (.A1(_09290_),
    .A2(_09443_),
    .B(_09448_),
    .Y(_01719_));
 AOI22x1_ASAP7_75t_R _16977_ (.A1(_00224_),
    .A2(_09435_),
    .B1(_09444_),
    .B2(_09214_),
    .Y(_09449_));
 OA21x2_ASAP7_75t_R _16978_ (.A1(_09292_),
    .A2(_09443_),
    .B(_09449_),
    .Y(_01720_));
 AOI22x1_ASAP7_75t_R _16979_ (.A1(_00191_),
    .A2(_09435_),
    .B1(_09444_),
    .B2(_09216_),
    .Y(_09450_));
 OA21x2_ASAP7_75t_R _16980_ (.A1(_09294_),
    .A2(_09443_),
    .B(_09450_),
    .Y(_01721_));
 INVx1_ASAP7_75t_R _16981_ (.A(_00157_),
    .Y(_09451_));
 OA222x2_ASAP7_75t_R _16982_ (.A1(_09451_),
    .A2(_09418_),
    .B1(_09419_),
    .B2(_09296_),
    .C1(_09421_),
    .C2(_09219_),
    .Y(_01722_));
 AOI22x1_ASAP7_75t_R _16983_ (.A1(_00124_),
    .A2(_09441_),
    .B1(_09444_),
    .B2(_09220_),
    .Y(_09452_));
 OA21x2_ASAP7_75t_R _16984_ (.A1(_09297_),
    .A2(_09443_),
    .B(_09452_),
    .Y(_01723_));
 NOR2x1_ASAP7_75t_R _16985_ (.A(_01022_),
    .B(_09418_),
    .Y(_09453_));
 AO21x1_ASAP7_75t_R _16986_ (.A1(_09299_),
    .A2(_09418_),
    .B(_09453_),
    .Y(_01724_));
 AND3x2_ASAP7_75t_R _16987_ (.A(_08824_),
    .B(_08750_),
    .C(_09253_),
    .Y(_09454_));
 NOR2x1_ASAP7_75t_R _16988_ (.A(_00090_),
    .B(_09418_),
    .Y(_09455_));
 AO221x1_ASAP7_75t_R _16989_ (.A1(_09223_),
    .A2(_09418_),
    .B1(_09454_),
    .B2(_09302_),
    .C(_09455_),
    .Y(_01725_));
 AND2x2_ASAP7_75t_R _16990_ (.A(_00058_),
    .B(_09441_),
    .Y(_09456_));
 AOI221x1_ASAP7_75t_R _16991_ (.A1(_09226_),
    .A2(_09454_),
    .B1(_09427_),
    .B2(_09304_),
    .C(_09456_),
    .Y(_01726_));
 AOI22x1_ASAP7_75t_R _16992_ (.A1(_00989_),
    .A2(_09441_),
    .B1(_09444_),
    .B2(_09228_),
    .Y(_09457_));
 OA21x2_ASAP7_75t_R _16993_ (.A1(_09306_),
    .A2(_09443_),
    .B(_09457_),
    .Y(_01727_));
 NAND2x1_ASAP7_75t_R _16994_ (.A(_00956_),
    .B(_09441_),
    .Y(_09458_));
 OA221x2_ASAP7_75t_R _16995_ (.A1(_09308_),
    .A2(_09424_),
    .B1(_09419_),
    .B2(_09230_),
    .C(_09458_),
    .Y(_01728_));
 NAND2x1_ASAP7_75t_R _16996_ (.A(_00922_),
    .B(_09441_),
    .Y(_09459_));
 OA221x2_ASAP7_75t_R _16997_ (.A1(_09232_),
    .A2(_09424_),
    .B1(_09419_),
    .B2(_09310_),
    .C(_09459_),
    .Y(_01729_));
 AOI22x1_ASAP7_75t_R _16998_ (.A1(_00889_),
    .A2(_09441_),
    .B1(_09444_),
    .B2(_09234_),
    .Y(_09460_));
 OA21x2_ASAP7_75t_R _16999_ (.A1(_09312_),
    .A2(_09443_),
    .B(_09460_),
    .Y(_01730_));
 NAND2x1_ASAP7_75t_R _17000_ (.A(_00855_),
    .B(_09423_),
    .Y(_09461_));
 OA21x2_ASAP7_75t_R _17001_ (.A1(_09315_),
    .A2(_09441_),
    .B(_09461_),
    .Y(_09462_));
 OA21x2_ASAP7_75t_R _17002_ (.A1(_09314_),
    .A2(_09443_),
    .B(_09462_),
    .Y(_01731_));
 AOI22x1_ASAP7_75t_R _17003_ (.A1(_00822_),
    .A2(_09441_),
    .B1(_09444_),
    .B2(_09238_),
    .Y(_09463_));
 OA21x2_ASAP7_75t_R _17004_ (.A1(_09318_),
    .A2(_09419_),
    .B(_09463_),
    .Y(_01732_));
 NAND2x1_ASAP7_75t_R _17005_ (.A(_00788_),
    .B(_09423_),
    .Y(_09464_));
 OA21x2_ASAP7_75t_R _17006_ (.A1(_09321_),
    .A2(_09441_),
    .B(_09464_),
    .Y(_09465_));
 OA21x2_ASAP7_75t_R _17007_ (.A1(_09320_),
    .A2(_09419_),
    .B(_09465_),
    .Y(_01733_));
 AND4x2_ASAP7_75t_R _17008_ (.A(_03025_),
    .B(net5),
    .C(net2),
    .D(_08100_),
    .Y(_09466_));
 AND2x6_ASAP7_75t_R _17009_ (.A(_08787_),
    .B(_09466_),
    .Y(_09467_));
 NAND2x2_ASAP7_75t_R _17010_ (.A(_09324_),
    .B(_09467_),
    .Y(_09468_));
 BUFx10_ASAP7_75t_R _17011_ (.A(_09468_),
    .Y(_09469_));
 NAND2x2_ASAP7_75t_R _17012_ (.A(_08114_),
    .B(_09467_),
    .Y(_09470_));
 OA22x2_ASAP7_75t_R _17013_ (.A1(_03168_),
    .A2(_09467_),
    .B1(_09470_),
    .B2(_09330_),
    .Y(_09471_));
 OA21x2_ASAP7_75t_R _17014_ (.A1(_09167_),
    .A2(_09469_),
    .B(_09471_),
    .Y(_01734_));
 BUFx12_ASAP7_75t_R _17015_ (.A(_09466_),
    .Y(_09472_));
 NAND2x2_ASAP7_75t_R _17016_ (.A(_08787_),
    .B(_09472_),
    .Y(_09473_));
 BUFx12f_ASAP7_75t_R _17017_ (.A(_09473_),
    .Y(_09474_));
 AND3x2_ASAP7_75t_R _17018_ (.A(_09425_),
    .B(_08795_),
    .C(_09472_),
    .Y(_09475_));
 BUFx12_ASAP7_75t_R _17019_ (.A(_09475_),
    .Y(_09476_));
 AOI22x1_ASAP7_75t_R _17020_ (.A1(_00756_),
    .A2(_09474_),
    .B1(_09476_),
    .B2(_09178_),
    .Y(_09477_));
 OA21x2_ASAP7_75t_R _17021_ (.A1(_09251_),
    .A2(_09469_),
    .B(_09477_),
    .Y(_01735_));
 AOI22x1_ASAP7_75t_R _17022_ (.A1(_00723_),
    .A2(_09474_),
    .B1(_09476_),
    .B2(_09180_),
    .Y(_09478_));
 OA21x2_ASAP7_75t_R _17023_ (.A1(_09257_),
    .A2(_09469_),
    .B(_09478_),
    .Y(_01736_));
 INVx1_ASAP7_75t_R _17024_ (.A(_00690_),
    .Y(_09479_));
 OA222x2_ASAP7_75t_R _17025_ (.A1(_09479_),
    .A2(_09467_),
    .B1(_09468_),
    .B2(_09260_),
    .C1(_09470_),
    .C2(_09182_),
    .Y(_01737_));
 INVx1_ASAP7_75t_R _17026_ (.A(_00657_),
    .Y(_09480_));
 OA222x2_ASAP7_75t_R _17027_ (.A1(_09480_),
    .A2(_09467_),
    .B1(_09468_),
    .B2(_09261_),
    .C1(_09470_),
    .C2(_09184_),
    .Y(_01738_));
 AOI22x1_ASAP7_75t_R _17028_ (.A1(_00624_),
    .A2(_09474_),
    .B1(_09476_),
    .B2(_09185_),
    .Y(_09481_));
 OA21x2_ASAP7_75t_R _17029_ (.A1(_09262_),
    .A2(_09469_),
    .B(_09481_),
    .Y(_01739_));
 AOI22x1_ASAP7_75t_R _17030_ (.A1(_00590_),
    .A2(_09474_),
    .B1(_09476_),
    .B2(_09187_),
    .Y(_09482_));
 OA21x2_ASAP7_75t_R _17031_ (.A1(_09264_),
    .A2(_09469_),
    .B(_09482_),
    .Y(_01740_));
 AOI22x1_ASAP7_75t_R _17032_ (.A1(_00557_),
    .A2(_09474_),
    .B1(_09476_),
    .B2(_09189_),
    .Y(_09483_));
 OA21x2_ASAP7_75t_R _17033_ (.A1(_09266_),
    .A2(_09469_),
    .B(_09483_),
    .Y(_01741_));
 BUFx12f_ASAP7_75t_R _17034_ (.A(_09473_),
    .Y(_09484_));
 AOI22x1_ASAP7_75t_R _17035_ (.A1(_00524_),
    .A2(_09484_),
    .B1(_09476_),
    .B2(_09192_),
    .Y(_09485_));
 OA21x2_ASAP7_75t_R _17036_ (.A1(_09268_),
    .A2(_09469_),
    .B(_09485_),
    .Y(_01742_));
 AOI22x1_ASAP7_75t_R _17037_ (.A1(_00491_),
    .A2(_09484_),
    .B1(_09476_),
    .B2(_09194_),
    .Y(_09486_));
 OA21x2_ASAP7_75t_R _17038_ (.A1(_09271_),
    .A2(_09469_),
    .B(_09486_),
    .Y(_01743_));
 AOI22x1_ASAP7_75t_R _17039_ (.A1(_00458_),
    .A2(_09484_),
    .B1(_09476_),
    .B2(_09196_),
    .Y(_09487_));
 OA21x2_ASAP7_75t_R _17040_ (.A1(_09273_),
    .A2(_09469_),
    .B(_09487_),
    .Y(_01744_));
 NAND2x1_ASAP7_75t_R _17041_ (.A(_01056_),
    .B(_09474_),
    .Y(_09488_));
 OA21x2_ASAP7_75t_R _17042_ (.A1(_09275_),
    .A2(_09474_),
    .B(_09488_),
    .Y(_01745_));
 AOI22x1_ASAP7_75t_R _17043_ (.A1(_00425_),
    .A2(_09484_),
    .B1(_09476_),
    .B2(_09199_),
    .Y(_09489_));
 OA21x2_ASAP7_75t_R _17044_ (.A1(_09277_),
    .A2(_09469_),
    .B(_09489_),
    .Y(_01746_));
 BUFx10_ASAP7_75t_R _17045_ (.A(_09473_),
    .Y(_09490_));
 NAND2x1_ASAP7_75t_R _17046_ (.A(_00392_),
    .B(_09490_),
    .Y(_09491_));
 OA221x2_ASAP7_75t_R _17047_ (.A1(_09201_),
    .A2(_09474_),
    .B1(_09468_),
    .B2(_09279_),
    .C(_09491_),
    .Y(_01747_));
 BUFx4f_ASAP7_75t_R _17048_ (.A(_09468_),
    .Y(_09492_));
 BUFx10_ASAP7_75t_R _17049_ (.A(_09475_),
    .Y(_09493_));
 AOI22x1_ASAP7_75t_R _17050_ (.A1(_00359_),
    .A2(_09484_),
    .B1(_09493_),
    .B2(_09206_),
    .Y(_09494_));
 OA21x2_ASAP7_75t_R _17051_ (.A1(_09282_),
    .A2(_09492_),
    .B(_09494_),
    .Y(_01748_));
 AOI22x1_ASAP7_75t_R _17052_ (.A1(_00325_),
    .A2(_09484_),
    .B1(_09493_),
    .B2(_09208_),
    .Y(_09495_));
 OA21x2_ASAP7_75t_R _17053_ (.A1(_09286_),
    .A2(_09492_),
    .B(_09495_),
    .Y(_01749_));
 AOI22x1_ASAP7_75t_R _17054_ (.A1(_00292_),
    .A2(_09484_),
    .B1(_09493_),
    .B2(_09210_),
    .Y(_09496_));
 OA21x2_ASAP7_75t_R _17055_ (.A1(_09288_),
    .A2(_09492_),
    .B(_09496_),
    .Y(_01750_));
 AOI22x1_ASAP7_75t_R _17056_ (.A1(_00259_),
    .A2(_09484_),
    .B1(_09493_),
    .B2(_09212_),
    .Y(_09497_));
 OA21x2_ASAP7_75t_R _17057_ (.A1(_09290_),
    .A2(_09492_),
    .B(_09497_),
    .Y(_01751_));
 AOI22x1_ASAP7_75t_R _17058_ (.A1(_00225_),
    .A2(_09484_),
    .B1(_09493_),
    .B2(_09214_),
    .Y(_09498_));
 OA21x2_ASAP7_75t_R _17059_ (.A1(_09292_),
    .A2(_09492_),
    .B(_09498_),
    .Y(_01752_));
 AOI22x1_ASAP7_75t_R _17060_ (.A1(_00192_),
    .A2(_09484_),
    .B1(_09493_),
    .B2(_09216_),
    .Y(_09499_));
 OA21x2_ASAP7_75t_R _17061_ (.A1(_09294_),
    .A2(_09492_),
    .B(_09499_),
    .Y(_01753_));
 INVx1_ASAP7_75t_R _17062_ (.A(_00158_),
    .Y(_09500_));
 OA222x2_ASAP7_75t_R _17063_ (.A1(_09500_),
    .A2(_09467_),
    .B1(_09468_),
    .B2(_09296_),
    .C1(_09470_),
    .C2(_09219_),
    .Y(_01754_));
 AOI22x1_ASAP7_75t_R _17064_ (.A1(_00125_),
    .A2(_09490_),
    .B1(_09493_),
    .B2(_09220_),
    .Y(_09501_));
 OA21x2_ASAP7_75t_R _17065_ (.A1(_09297_),
    .A2(_09492_),
    .B(_09501_),
    .Y(_01755_));
 NOR2x1_ASAP7_75t_R _17066_ (.A(_01023_),
    .B(_09467_),
    .Y(_09502_));
 AO21x1_ASAP7_75t_R _17067_ (.A1(_09299_),
    .A2(_09467_),
    .B(_09502_),
    .Y(_01756_));
 BUFx4f_ASAP7_75t_R _17068_ (.A(_08687_),
    .Y(_09503_));
 BUFx6f_ASAP7_75t_R _17069_ (.A(_09472_),
    .Y(_09504_));
 AND3x1_ASAP7_75t_R _17070_ (.A(_09503_),
    .B(_08788_),
    .C(_09504_),
    .Y(_09505_));
 NOR2x1_ASAP7_75t_R _17071_ (.A(_00091_),
    .B(_09467_),
    .Y(_09506_));
 AO221x1_ASAP7_75t_R _17072_ (.A1(_09223_),
    .A2(_09467_),
    .B1(_09505_),
    .B2(_09302_),
    .C(_09506_),
    .Y(_01757_));
 AND2x2_ASAP7_75t_R _17073_ (.A(_00059_),
    .B(_09490_),
    .Y(_09507_));
 AOI221x1_ASAP7_75t_R _17074_ (.A1(_09226_),
    .A2(_09505_),
    .B1(_09476_),
    .B2(_09304_),
    .C(_09507_),
    .Y(_01758_));
 AOI22x1_ASAP7_75t_R _17075_ (.A1(_00990_),
    .A2(_09490_),
    .B1(_09493_),
    .B2(_09228_),
    .Y(_09508_));
 OA21x2_ASAP7_75t_R _17076_ (.A1(_09306_),
    .A2(_09492_),
    .B(_09508_),
    .Y(_01759_));
 NAND2x1_ASAP7_75t_R _17077_ (.A(_00957_),
    .B(_09490_),
    .Y(_09509_));
 OA221x2_ASAP7_75t_R _17078_ (.A1(_09308_),
    .A2(_09474_),
    .B1(_09468_),
    .B2(_09230_),
    .C(_09509_),
    .Y(_01760_));
 NAND2x1_ASAP7_75t_R _17079_ (.A(_00923_),
    .B(_09490_),
    .Y(_09510_));
 OA221x2_ASAP7_75t_R _17080_ (.A1(_09232_),
    .A2(_09474_),
    .B1(_09468_),
    .B2(_09310_),
    .C(_09510_),
    .Y(_01761_));
 AOI22x1_ASAP7_75t_R _17081_ (.A1(_00890_),
    .A2(_09490_),
    .B1(_09493_),
    .B2(_09234_),
    .Y(_09511_));
 OA21x2_ASAP7_75t_R _17082_ (.A1(_09312_),
    .A2(_09492_),
    .B(_09511_),
    .Y(_01762_));
 NAND2x1_ASAP7_75t_R _17083_ (.A(_00856_),
    .B(_09473_),
    .Y(_09512_));
 OA21x2_ASAP7_75t_R _17084_ (.A1(_09315_),
    .A2(_09490_),
    .B(_09512_),
    .Y(_09513_));
 OA21x2_ASAP7_75t_R _17085_ (.A1(_09314_),
    .A2(_09492_),
    .B(_09513_),
    .Y(_01763_));
 AOI22x1_ASAP7_75t_R _17086_ (.A1(_00823_),
    .A2(_09490_),
    .B1(_09493_),
    .B2(_09238_),
    .Y(_09514_));
 OA21x2_ASAP7_75t_R _17087_ (.A1(_09318_),
    .A2(_09468_),
    .B(_09514_),
    .Y(_01764_));
 NAND2x1_ASAP7_75t_R _17088_ (.A(_00789_),
    .B(_09473_),
    .Y(_09515_));
 OA21x2_ASAP7_75t_R _17089_ (.A1(_09321_),
    .A2(_09490_),
    .B(_09515_),
    .Y(_09516_));
 OA21x2_ASAP7_75t_R _17090_ (.A1(_09320_),
    .A2(_09468_),
    .B(_09516_),
    .Y(_01765_));
 AND2x6_ASAP7_75t_R _17091_ (.A(_08837_),
    .B(_09466_),
    .Y(_09517_));
 NAND2x2_ASAP7_75t_R _17092_ (.A(_09324_),
    .B(_09517_),
    .Y(_09518_));
 BUFx12_ASAP7_75t_R _17093_ (.A(_09518_),
    .Y(_09519_));
 NAND2x2_ASAP7_75t_R _17094_ (.A(_08114_),
    .B(_09517_),
    .Y(_09520_));
 OA22x2_ASAP7_75t_R _17095_ (.A1(_03165_),
    .A2(_09517_),
    .B1(_09520_),
    .B2(_09330_),
    .Y(_09521_));
 OA21x2_ASAP7_75t_R _17096_ (.A1(_09167_),
    .A2(_09519_),
    .B(_09521_),
    .Y(_01766_));
 NAND2x2_ASAP7_75t_R _17097_ (.A(_08847_),
    .B(_09472_),
    .Y(_09522_));
 BUFx16f_ASAP7_75t_R _17098_ (.A(_09522_),
    .Y(_09523_));
 AND3x2_ASAP7_75t_R _17099_ (.A(_09425_),
    .B(_08847_),
    .C(_09472_),
    .Y(_09524_));
 BUFx12_ASAP7_75t_R _17100_ (.A(_09524_),
    .Y(_09525_));
 AOI22x1_ASAP7_75t_R _17101_ (.A1(_00757_),
    .A2(_09523_),
    .B1(_09525_),
    .B2(_09178_),
    .Y(_09526_));
 OA21x2_ASAP7_75t_R _17102_ (.A1(_09251_),
    .A2(_09519_),
    .B(_09526_),
    .Y(_01767_));
 AOI22x1_ASAP7_75t_R _17103_ (.A1(_00724_),
    .A2(_09523_),
    .B1(_09525_),
    .B2(_09180_),
    .Y(_09527_));
 OA21x2_ASAP7_75t_R _17104_ (.A1(_09257_),
    .A2(_09519_),
    .B(_09527_),
    .Y(_01768_));
 OA222x2_ASAP7_75t_R _17105_ (.A1(_05756_),
    .A2(_09517_),
    .B1(_09518_),
    .B2(_09260_),
    .C1(_09520_),
    .C2(_09182_),
    .Y(_01769_));
 OA222x2_ASAP7_75t_R _17106_ (.A1(_05616_),
    .A2(_09517_),
    .B1(_09518_),
    .B2(_09261_),
    .C1(_09520_),
    .C2(_09184_),
    .Y(_01770_));
 AOI22x1_ASAP7_75t_R _17107_ (.A1(_00625_),
    .A2(_09523_),
    .B1(_09525_),
    .B2(_09185_),
    .Y(_09528_));
 OA21x2_ASAP7_75t_R _17108_ (.A1(_09262_),
    .A2(_09519_),
    .B(_09528_),
    .Y(_01771_));
 AOI22x1_ASAP7_75t_R _17109_ (.A1(_00591_),
    .A2(_09523_),
    .B1(_09525_),
    .B2(_09187_),
    .Y(_09529_));
 OA21x2_ASAP7_75t_R _17110_ (.A1(_09264_),
    .A2(_09519_),
    .B(_09529_),
    .Y(_01772_));
 AOI22x1_ASAP7_75t_R _17111_ (.A1(_00558_),
    .A2(_09523_),
    .B1(_09525_),
    .B2(_09189_),
    .Y(_09530_));
 OA21x2_ASAP7_75t_R _17112_ (.A1(_09266_),
    .A2(_09519_),
    .B(_09530_),
    .Y(_01773_));
 AOI22x1_ASAP7_75t_R _17113_ (.A1(_00525_),
    .A2(_09523_),
    .B1(_09525_),
    .B2(_09192_),
    .Y(_09531_));
 OA21x2_ASAP7_75t_R _17114_ (.A1(_09268_),
    .A2(_09519_),
    .B(_09531_),
    .Y(_01774_));
 BUFx12f_ASAP7_75t_R _17115_ (.A(_09522_),
    .Y(_09532_));
 AOI22x1_ASAP7_75t_R _17116_ (.A1(_00492_),
    .A2(_09532_),
    .B1(_09525_),
    .B2(_09194_),
    .Y(_09533_));
 OA21x2_ASAP7_75t_R _17117_ (.A1(_09271_),
    .A2(_09519_),
    .B(_09533_),
    .Y(_01775_));
 AOI22x1_ASAP7_75t_R _17118_ (.A1(_00459_),
    .A2(_09532_),
    .B1(_09525_),
    .B2(_09196_),
    .Y(_09534_));
 OA21x2_ASAP7_75t_R _17119_ (.A1(_09273_),
    .A2(_09519_),
    .B(_09534_),
    .Y(_01776_));
 AO21x1_ASAP7_75t_R _17120_ (.A1(_09051_),
    .A2(_09504_),
    .B(_06784_),
    .Y(_09535_));
 OA21x2_ASAP7_75t_R _17121_ (.A1(_09275_),
    .A2(_09523_),
    .B(_09535_),
    .Y(_01777_));
 AOI22x1_ASAP7_75t_R _17122_ (.A1(_00426_),
    .A2(_09532_),
    .B1(_09525_),
    .B2(_09199_),
    .Y(_09536_));
 OA21x2_ASAP7_75t_R _17123_ (.A1(_09277_),
    .A2(_09519_),
    .B(_09536_),
    .Y(_01778_));
 AO21x1_ASAP7_75t_R _17124_ (.A1(_09051_),
    .A2(_09504_),
    .B(_04820_),
    .Y(_09537_));
 OA221x2_ASAP7_75t_R _17125_ (.A1(_09201_),
    .A2(_09523_),
    .B1(_09518_),
    .B2(_09279_),
    .C(_09537_),
    .Y(_01779_));
 BUFx4f_ASAP7_75t_R _17126_ (.A(_09518_),
    .Y(_09538_));
 BUFx6f_ASAP7_75t_R _17127_ (.A(_09524_),
    .Y(_09539_));
 AOI22x1_ASAP7_75t_R _17128_ (.A1(_00360_),
    .A2(_09532_),
    .B1(_09539_),
    .B2(_09206_),
    .Y(_09540_));
 OA21x2_ASAP7_75t_R _17129_ (.A1(_09282_),
    .A2(_09538_),
    .B(_09540_),
    .Y(_01780_));
 AOI22x1_ASAP7_75t_R _17130_ (.A1(_00326_),
    .A2(_09532_),
    .B1(_09539_),
    .B2(_09208_),
    .Y(_09541_));
 OA21x2_ASAP7_75t_R _17131_ (.A1(_09286_),
    .A2(_09538_),
    .B(_09541_),
    .Y(_01781_));
 AOI22x1_ASAP7_75t_R _17132_ (.A1(_00293_),
    .A2(_09532_),
    .B1(_09539_),
    .B2(_09210_),
    .Y(_09542_));
 OA21x2_ASAP7_75t_R _17133_ (.A1(_09288_),
    .A2(_09538_),
    .B(_09542_),
    .Y(_01782_));
 AOI22x1_ASAP7_75t_R _17134_ (.A1(_00260_),
    .A2(_09532_),
    .B1(_09539_),
    .B2(_09212_),
    .Y(_09543_));
 OA21x2_ASAP7_75t_R _17135_ (.A1(_09290_),
    .A2(_09538_),
    .B(_09543_),
    .Y(_01783_));
 AOI22x1_ASAP7_75t_R _17136_ (.A1(_00226_),
    .A2(_09532_),
    .B1(_09539_),
    .B2(_09214_),
    .Y(_09544_));
 OA21x2_ASAP7_75t_R _17137_ (.A1(_09292_),
    .A2(_09538_),
    .B(_09544_),
    .Y(_01784_));
 AOI22x1_ASAP7_75t_R _17138_ (.A1(_00193_),
    .A2(_09532_),
    .B1(_09539_),
    .B2(_09216_),
    .Y(_09545_));
 OA21x2_ASAP7_75t_R _17139_ (.A1(_09294_),
    .A2(_09538_),
    .B(_09545_),
    .Y(_01785_));
 INVx1_ASAP7_75t_R _17140_ (.A(_00159_),
    .Y(_09546_));
 OA222x2_ASAP7_75t_R _17141_ (.A1(_09546_),
    .A2(_09517_),
    .B1(_09518_),
    .B2(_09296_),
    .C1(_09520_),
    .C2(_09219_),
    .Y(_01786_));
 AOI22x1_ASAP7_75t_R _17142_ (.A1(_00126_),
    .A2(_09532_),
    .B1(_09539_),
    .B2(_09220_),
    .Y(_09547_));
 OA21x2_ASAP7_75t_R _17143_ (.A1(_09297_),
    .A2(_09538_),
    .B(_09547_),
    .Y(_01787_));
 NOR2x1_ASAP7_75t_R _17144_ (.A(_01024_),
    .B(_09517_),
    .Y(_02246_));
 AO21x1_ASAP7_75t_R _17145_ (.A1(_09299_),
    .A2(_09517_),
    .B(_02246_),
    .Y(_01788_));
 AND3x1_ASAP7_75t_R _17146_ (.A(_09503_),
    .B(_09051_),
    .C(_09504_),
    .Y(_02247_));
 NOR2x1_ASAP7_75t_R _17147_ (.A(_00092_),
    .B(_09517_),
    .Y(_02248_));
 AO221x1_ASAP7_75t_R _17148_ (.A1(_09223_),
    .A2(_09517_),
    .B1(_02247_),
    .B2(_09302_),
    .C(_02248_),
    .Y(_01789_));
 BUFx10_ASAP7_75t_R _17149_ (.A(_09522_),
    .Y(_02249_));
 AND2x2_ASAP7_75t_R _17150_ (.A(_00060_),
    .B(_02249_),
    .Y(_02250_));
 AOI221x1_ASAP7_75t_R _17151_ (.A1(_09226_),
    .A2(_02247_),
    .B1(_09525_),
    .B2(_09304_),
    .C(_02250_),
    .Y(_01790_));
 AOI22x1_ASAP7_75t_R _17152_ (.A1(_00991_),
    .A2(_02249_),
    .B1(_09539_),
    .B2(_09228_),
    .Y(_02251_));
 OA21x2_ASAP7_75t_R _17153_ (.A1(_09306_),
    .A2(_09538_),
    .B(_02251_),
    .Y(_01791_));
 NAND2x1_ASAP7_75t_R _17154_ (.A(_00958_),
    .B(_02249_),
    .Y(_02252_));
 OA221x2_ASAP7_75t_R _17155_ (.A1(_09308_),
    .A2(_09523_),
    .B1(_09518_),
    .B2(_09230_),
    .C(_02252_),
    .Y(_01792_));
 NAND2x1_ASAP7_75t_R _17156_ (.A(_00924_),
    .B(_02249_),
    .Y(_02253_));
 OA221x2_ASAP7_75t_R _17157_ (.A1(_09232_),
    .A2(_09523_),
    .B1(_09518_),
    .B2(_09310_),
    .C(_02253_),
    .Y(_01793_));
 AOI22x1_ASAP7_75t_R _17158_ (.A1(_00891_),
    .A2(_02249_),
    .B1(_09539_),
    .B2(_09234_),
    .Y(_02254_));
 OA21x2_ASAP7_75t_R _17159_ (.A1(_09312_),
    .A2(_09538_),
    .B(_02254_),
    .Y(_01794_));
 NAND2x1_ASAP7_75t_R _17160_ (.A(_00857_),
    .B(_02249_),
    .Y(_02255_));
 OA21x2_ASAP7_75t_R _17161_ (.A1(_09315_),
    .A2(_02249_),
    .B(_02255_),
    .Y(_02256_));
 OA21x2_ASAP7_75t_R _17162_ (.A1(_09314_),
    .A2(_09538_),
    .B(_02256_),
    .Y(_01795_));
 AOI22x1_ASAP7_75t_R _17163_ (.A1(_00824_),
    .A2(_02249_),
    .B1(_09539_),
    .B2(_09238_),
    .Y(_02257_));
 OA21x2_ASAP7_75t_R _17164_ (.A1(_09318_),
    .A2(_09518_),
    .B(_02257_),
    .Y(_01796_));
 NAND2x1_ASAP7_75t_R _17165_ (.A(_00790_),
    .B(_02249_),
    .Y(_02258_));
 OA21x2_ASAP7_75t_R _17166_ (.A1(_09321_),
    .A2(_02249_),
    .B(_02258_),
    .Y(_02259_));
 OA21x2_ASAP7_75t_R _17167_ (.A1(_09320_),
    .A2(_09518_),
    .B(_02259_),
    .Y(_01797_));
 AND2x6_ASAP7_75t_R _17168_ (.A(_08098_),
    .B(_09472_),
    .Y(_02260_));
 NAND2x2_ASAP7_75t_R _17169_ (.A(_09324_),
    .B(_02260_),
    .Y(_02261_));
 BUFx10_ASAP7_75t_R _17170_ (.A(_02261_),
    .Y(_02262_));
 NAND2x2_ASAP7_75t_R _17171_ (.A(_08115_),
    .B(_02260_),
    .Y(_02263_));
 NAND2x2_ASAP7_75t_R _17172_ (.A(_08098_),
    .B(_09472_),
    .Y(_02264_));
 NAND2x1_ASAP7_75t_R _17173_ (.A(_00026_),
    .B(_02264_),
    .Y(_02265_));
 OA21x2_ASAP7_75t_R _17174_ (.A1(_08111_),
    .A2(_02263_),
    .B(_02265_),
    .Y(_02266_));
 OA21x2_ASAP7_75t_R _17175_ (.A1(_09167_),
    .A2(_02262_),
    .B(_02266_),
    .Y(_01798_));
 BUFx12f_ASAP7_75t_R _17176_ (.A(_02264_),
    .Y(_02267_));
 AND3x2_ASAP7_75t_R _17177_ (.A(_08117_),
    .B(_08701_),
    .C(_09472_),
    .Y(_02268_));
 BUFx12_ASAP7_75t_R _17178_ (.A(_02268_),
    .Y(_02269_));
 AOI22x1_ASAP7_75t_R _17179_ (.A1(_00758_),
    .A2(_02267_),
    .B1(_02269_),
    .B2(_09178_),
    .Y(_02270_));
 OA21x2_ASAP7_75t_R _17180_ (.A1(_09251_),
    .A2(_02262_),
    .B(_02270_),
    .Y(_01799_));
 AOI22x1_ASAP7_75t_R _17181_ (.A1(_00725_),
    .A2(_02267_),
    .B1(_02269_),
    .B2(_09180_),
    .Y(_02271_));
 OA21x2_ASAP7_75t_R _17182_ (.A1(_09257_),
    .A2(_02262_),
    .B(_02271_),
    .Y(_01800_));
 OA222x2_ASAP7_75t_R _17183_ (.A1(_05761_),
    .A2(_02260_),
    .B1(_02261_),
    .B2(_09260_),
    .C1(_02263_),
    .C2(_09182_),
    .Y(_01801_));
 INVx1_ASAP7_75t_R _17184_ (.A(_00659_),
    .Y(_02272_));
 OA222x2_ASAP7_75t_R _17185_ (.A1(_02272_),
    .A2(_02260_),
    .B1(_02261_),
    .B2(_09261_),
    .C1(_02263_),
    .C2(_09184_),
    .Y(_01802_));
 AOI22x1_ASAP7_75t_R _17186_ (.A1(_00626_),
    .A2(_02267_),
    .B1(_02269_),
    .B2(_09185_),
    .Y(_02273_));
 OA21x2_ASAP7_75t_R _17187_ (.A1(_09262_),
    .A2(_02262_),
    .B(_02273_),
    .Y(_01803_));
 AOI22x1_ASAP7_75t_R _17188_ (.A1(_00592_),
    .A2(_02267_),
    .B1(_02269_),
    .B2(_09187_),
    .Y(_02274_));
 OA21x2_ASAP7_75t_R _17189_ (.A1(_09264_),
    .A2(_02262_),
    .B(_02274_),
    .Y(_01804_));
 AOI22x1_ASAP7_75t_R _17190_ (.A1(_00559_),
    .A2(_02267_),
    .B1(_02269_),
    .B2(_09189_),
    .Y(_02275_));
 OA21x2_ASAP7_75t_R _17191_ (.A1(_09266_),
    .A2(_02262_),
    .B(_02275_),
    .Y(_01805_));
 BUFx16f_ASAP7_75t_R _17192_ (.A(_02264_),
    .Y(_02276_));
 AOI22x1_ASAP7_75t_R _17193_ (.A1(_00526_),
    .A2(_02276_),
    .B1(_02269_),
    .B2(_09192_),
    .Y(_02277_));
 OA21x2_ASAP7_75t_R _17194_ (.A1(_09268_),
    .A2(_02262_),
    .B(_02277_),
    .Y(_01806_));
 AOI22x1_ASAP7_75t_R _17195_ (.A1(_00493_),
    .A2(_02276_),
    .B1(_02269_),
    .B2(_09194_),
    .Y(_02278_));
 OA21x2_ASAP7_75t_R _17196_ (.A1(_09271_),
    .A2(_02262_),
    .B(_02278_),
    .Y(_01807_));
 AOI22x1_ASAP7_75t_R _17197_ (.A1(_00460_),
    .A2(_02276_),
    .B1(_02269_),
    .B2(_09196_),
    .Y(_02279_));
 OA21x2_ASAP7_75t_R _17198_ (.A1(_09273_),
    .A2(_02262_),
    .B(_02279_),
    .Y(_01808_));
 NAND2x1_ASAP7_75t_R _17199_ (.A(_01058_),
    .B(_02267_),
    .Y(_02280_));
 OA21x2_ASAP7_75t_R _17200_ (.A1(_09275_),
    .A2(_02267_),
    .B(_02280_),
    .Y(_01809_));
 AOI22x1_ASAP7_75t_R _17201_ (.A1(_00427_),
    .A2(_02276_),
    .B1(_02269_),
    .B2(_09199_),
    .Y(_02281_));
 OA21x2_ASAP7_75t_R _17202_ (.A1(_09277_),
    .A2(_02262_),
    .B(_02281_),
    .Y(_01810_));
 BUFx10_ASAP7_75t_R _17203_ (.A(_02264_),
    .Y(_02282_));
 NAND2x1_ASAP7_75t_R _17204_ (.A(_00394_),
    .B(_02282_),
    .Y(_02283_));
 OA221x2_ASAP7_75t_R _17205_ (.A1(_09201_),
    .A2(_02267_),
    .B1(_02261_),
    .B2(_09279_),
    .C(_02283_),
    .Y(_01811_));
 BUFx4f_ASAP7_75t_R _17206_ (.A(_02261_),
    .Y(_02284_));
 BUFx6f_ASAP7_75t_R _17207_ (.A(_02268_),
    .Y(_02285_));
 AOI22x1_ASAP7_75t_R _17208_ (.A1(_00361_),
    .A2(_02276_),
    .B1(_02285_),
    .B2(_09206_),
    .Y(_02286_));
 OA21x2_ASAP7_75t_R _17209_ (.A1(_09282_),
    .A2(_02284_),
    .B(_02286_),
    .Y(_01812_));
 AOI22x1_ASAP7_75t_R _17210_ (.A1(_00327_),
    .A2(_02276_),
    .B1(_02285_),
    .B2(_09208_),
    .Y(_02287_));
 OA21x2_ASAP7_75t_R _17211_ (.A1(_09286_),
    .A2(_02284_),
    .B(_02287_),
    .Y(_01813_));
 AOI22x1_ASAP7_75t_R _17212_ (.A1(_00294_),
    .A2(_02276_),
    .B1(_02285_),
    .B2(_09210_),
    .Y(_02288_));
 OA21x2_ASAP7_75t_R _17213_ (.A1(_09288_),
    .A2(_02284_),
    .B(_02288_),
    .Y(_01814_));
 AOI22x1_ASAP7_75t_R _17214_ (.A1(_00261_),
    .A2(_02276_),
    .B1(_02285_),
    .B2(_09212_),
    .Y(_02289_));
 OA21x2_ASAP7_75t_R _17215_ (.A1(_09290_),
    .A2(_02284_),
    .B(_02289_),
    .Y(_01815_));
 AOI22x1_ASAP7_75t_R _17216_ (.A1(_00227_),
    .A2(_02276_),
    .B1(_02285_),
    .B2(_09214_),
    .Y(_02290_));
 OA21x2_ASAP7_75t_R _17217_ (.A1(_09292_),
    .A2(_02284_),
    .B(_02290_),
    .Y(_01816_));
 AOI22x1_ASAP7_75t_R _17218_ (.A1(_00194_),
    .A2(_02276_),
    .B1(_02285_),
    .B2(_09216_),
    .Y(_02291_));
 OA21x2_ASAP7_75t_R _17219_ (.A1(_09294_),
    .A2(_02284_),
    .B(_02291_),
    .Y(_01817_));
 INVx1_ASAP7_75t_R _17220_ (.A(_00160_),
    .Y(_02292_));
 OA222x2_ASAP7_75t_R _17221_ (.A1(_02292_),
    .A2(_02260_),
    .B1(_02261_),
    .B2(_09296_),
    .C1(_02263_),
    .C2(_09219_),
    .Y(_01818_));
 AOI22x1_ASAP7_75t_R _17222_ (.A1(_00127_),
    .A2(_02282_),
    .B1(_02285_),
    .B2(_09220_),
    .Y(_02293_));
 OA21x2_ASAP7_75t_R _17223_ (.A1(_09297_),
    .A2(_02284_),
    .B(_02293_),
    .Y(_01819_));
 NOR2x1_ASAP7_75t_R _17224_ (.A(_01025_),
    .B(_02260_),
    .Y(_02294_));
 AO21x1_ASAP7_75t_R _17225_ (.A1(_09299_),
    .A2(_02260_),
    .B(_02294_),
    .Y(_01820_));
 AND3x1_ASAP7_75t_R _17226_ (.A(_08145_),
    .B(_08577_),
    .C(_09504_),
    .Y(_02295_));
 NOR2x1_ASAP7_75t_R _17227_ (.A(_00093_),
    .B(_02260_),
    .Y(_02296_));
 AO221x1_ASAP7_75t_R _17228_ (.A1(_09223_),
    .A2(_02260_),
    .B1(_02295_),
    .B2(_09302_),
    .C(_02296_),
    .Y(_01821_));
 AND2x2_ASAP7_75t_R _17229_ (.A(_00061_),
    .B(_02282_),
    .Y(_02297_));
 AOI221x1_ASAP7_75t_R _17230_ (.A1(_09226_),
    .A2(_02295_),
    .B1(_02269_),
    .B2(_09304_),
    .C(_02297_),
    .Y(_01822_));
 AOI22x1_ASAP7_75t_R _17231_ (.A1(_00992_),
    .A2(_02282_),
    .B1(_02285_),
    .B2(_09228_),
    .Y(_02298_));
 OA21x2_ASAP7_75t_R _17232_ (.A1(_09306_),
    .A2(_02284_),
    .B(_02298_),
    .Y(_01823_));
 NAND2x1_ASAP7_75t_R _17233_ (.A(_00959_),
    .B(_02282_),
    .Y(_02299_));
 OA221x2_ASAP7_75t_R _17234_ (.A1(_09308_),
    .A2(_02267_),
    .B1(_02261_),
    .B2(_09230_),
    .C(_02299_),
    .Y(_01824_));
 NAND2x1_ASAP7_75t_R _17235_ (.A(_00925_),
    .B(_02282_),
    .Y(_02300_));
 OA221x2_ASAP7_75t_R _17236_ (.A1(_09232_),
    .A2(_02267_),
    .B1(_02261_),
    .B2(_09310_),
    .C(_02300_),
    .Y(_01825_));
 AOI22x1_ASAP7_75t_R _17237_ (.A1(_00892_),
    .A2(_02282_),
    .B1(_02285_),
    .B2(_09234_),
    .Y(_02301_));
 OA21x2_ASAP7_75t_R _17238_ (.A1(_09312_),
    .A2(_02284_),
    .B(_02301_),
    .Y(_01826_));
 NAND2x1_ASAP7_75t_R _17239_ (.A(_00858_),
    .B(_02264_),
    .Y(_02302_));
 OA21x2_ASAP7_75t_R _17240_ (.A1(_09315_),
    .A2(_02282_),
    .B(_02302_),
    .Y(_02303_));
 OA21x2_ASAP7_75t_R _17241_ (.A1(_09314_),
    .A2(_02284_),
    .B(_02303_),
    .Y(_01827_));
 AOI22x1_ASAP7_75t_R _17242_ (.A1(_00825_),
    .A2(_02282_),
    .B1(_02285_),
    .B2(_09238_),
    .Y(_02304_));
 OA21x2_ASAP7_75t_R _17243_ (.A1(_09318_),
    .A2(_02261_),
    .B(_02304_),
    .Y(_01828_));
 NAND2x1_ASAP7_75t_R _17244_ (.A(_00791_),
    .B(_02264_),
    .Y(_02305_));
 OA21x2_ASAP7_75t_R _17245_ (.A1(_09321_),
    .A2(_02282_),
    .B(_02305_),
    .Y(_02306_));
 OA21x2_ASAP7_75t_R _17246_ (.A1(_09320_),
    .A2(_02261_),
    .B(_02306_),
    .Y(_01829_));
 AND2x6_ASAP7_75t_R _17247_ (.A(_08689_),
    .B(_09466_),
    .Y(_02307_));
 NAND2x2_ASAP7_75t_R _17248_ (.A(_09324_),
    .B(_02307_),
    .Y(_02308_));
 BUFx12_ASAP7_75t_R _17249_ (.A(_02308_),
    .Y(_02309_));
 NAND2x2_ASAP7_75t_R _17250_ (.A(_08114_),
    .B(_02307_),
    .Y(_02310_));
 OA22x2_ASAP7_75t_R _17251_ (.A1(_03164_),
    .A2(_02307_),
    .B1(_02310_),
    .B2(_09330_),
    .Y(_02311_));
 OA21x2_ASAP7_75t_R _17252_ (.A1(_09167_),
    .A2(_02309_),
    .B(_02311_),
    .Y(_01830_));
 NAND2x2_ASAP7_75t_R _17253_ (.A(_08749_),
    .B(_09472_),
    .Y(_02312_));
 BUFx12f_ASAP7_75t_R _17254_ (.A(_02312_),
    .Y(_02313_));
 AND3x2_ASAP7_75t_R _17255_ (.A(_09425_),
    .B(_08749_),
    .C(_09472_),
    .Y(_02314_));
 BUFx12_ASAP7_75t_R _17256_ (.A(_02314_),
    .Y(_02315_));
 AOI22x1_ASAP7_75t_R _17257_ (.A1(_00759_),
    .A2(_02313_),
    .B1(_02315_),
    .B2(_09178_),
    .Y(_02316_));
 OA21x2_ASAP7_75t_R _17258_ (.A1(_09251_),
    .A2(_02309_),
    .B(_02316_),
    .Y(_01831_));
 AOI22x1_ASAP7_75t_R _17259_ (.A1(_00726_),
    .A2(_02313_),
    .B1(_02315_),
    .B2(_09180_),
    .Y(_02317_));
 OA21x2_ASAP7_75t_R _17260_ (.A1(_09257_),
    .A2(_02309_),
    .B(_02317_),
    .Y(_01832_));
 OA222x2_ASAP7_75t_R _17261_ (.A1(_05759_),
    .A2(_02307_),
    .B1(_02308_),
    .B2(_09260_),
    .C1(_02310_),
    .C2(_09182_),
    .Y(_01833_));
 INVx1_ASAP7_75t_R _17262_ (.A(_00660_),
    .Y(_02318_));
 OA222x2_ASAP7_75t_R _17263_ (.A1(_02318_),
    .A2(_02307_),
    .B1(_02308_),
    .B2(_09261_),
    .C1(_02310_),
    .C2(_09184_),
    .Y(_01834_));
 AOI22x1_ASAP7_75t_R _17264_ (.A1(_00627_),
    .A2(_02313_),
    .B1(_02315_),
    .B2(_09185_),
    .Y(_02319_));
 OA21x2_ASAP7_75t_R _17265_ (.A1(_09262_),
    .A2(_02309_),
    .B(_02319_),
    .Y(_01835_));
 AOI22x1_ASAP7_75t_R _17266_ (.A1(_00593_),
    .A2(_02313_),
    .B1(_02315_),
    .B2(_09187_),
    .Y(_02320_));
 OA21x2_ASAP7_75t_R _17267_ (.A1(_09264_),
    .A2(_02309_),
    .B(_02320_),
    .Y(_01836_));
 AOI22x1_ASAP7_75t_R _17268_ (.A1(_00560_),
    .A2(_02313_),
    .B1(_02315_),
    .B2(_09189_),
    .Y(_02321_));
 OA21x2_ASAP7_75t_R _17269_ (.A1(_09266_),
    .A2(_02309_),
    .B(_02321_),
    .Y(_01837_));
 AOI22x1_ASAP7_75t_R _17270_ (.A1(_00527_),
    .A2(_02313_),
    .B1(_02315_),
    .B2(_09192_),
    .Y(_02322_));
 OA21x2_ASAP7_75t_R _17271_ (.A1(_09268_),
    .A2(_02309_),
    .B(_02322_),
    .Y(_01838_));
 BUFx12f_ASAP7_75t_R _17272_ (.A(_02312_),
    .Y(_02323_));
 AOI22x1_ASAP7_75t_R _17273_ (.A1(_00494_),
    .A2(_02323_),
    .B1(_02315_),
    .B2(_09194_),
    .Y(_02324_));
 OA21x2_ASAP7_75t_R _17274_ (.A1(_09271_),
    .A2(_02309_),
    .B(_02324_),
    .Y(_01839_));
 AOI22x1_ASAP7_75t_R _17275_ (.A1(_00461_),
    .A2(_02323_),
    .B1(_02315_),
    .B2(_09196_),
    .Y(_02325_));
 OA21x2_ASAP7_75t_R _17276_ (.A1(_09273_),
    .A2(_02309_),
    .B(_02325_),
    .Y(_01840_));
 AO21x1_ASAP7_75t_R _17277_ (.A1(_09141_),
    .A2(_09504_),
    .B(_06787_),
    .Y(_02326_));
 OA21x2_ASAP7_75t_R _17278_ (.A1(_09275_),
    .A2(_02313_),
    .B(_02326_),
    .Y(_01841_));
 AOI22x1_ASAP7_75t_R _17279_ (.A1(_00428_),
    .A2(_02323_),
    .B1(_02315_),
    .B2(_09199_),
    .Y(_02327_));
 OA21x2_ASAP7_75t_R _17280_ (.A1(_09277_),
    .A2(_02309_),
    .B(_02327_),
    .Y(_01842_));
 AO21x1_ASAP7_75t_R _17281_ (.A1(_09141_),
    .A2(_09504_),
    .B(_04815_),
    .Y(_02328_));
 OA221x2_ASAP7_75t_R _17282_ (.A1(_09201_),
    .A2(_02313_),
    .B1(_02308_),
    .B2(_09279_),
    .C(_02328_),
    .Y(_01843_));
 BUFx6f_ASAP7_75t_R _17283_ (.A(_02308_),
    .Y(_02329_));
 BUFx10_ASAP7_75t_R _17284_ (.A(_02314_),
    .Y(_02330_));
 AOI22x1_ASAP7_75t_R _17285_ (.A1(_00362_),
    .A2(_02323_),
    .B1(_02330_),
    .B2(_09206_),
    .Y(_02331_));
 OA21x2_ASAP7_75t_R _17286_ (.A1(_09282_),
    .A2(_02329_),
    .B(_02331_),
    .Y(_01844_));
 AOI22x1_ASAP7_75t_R _17287_ (.A1(_00328_),
    .A2(_02323_),
    .B1(_02330_),
    .B2(_09208_),
    .Y(_02332_));
 OA21x2_ASAP7_75t_R _17288_ (.A1(_09286_),
    .A2(_02329_),
    .B(_02332_),
    .Y(_01845_));
 AOI22x1_ASAP7_75t_R _17289_ (.A1(_00295_),
    .A2(_02323_),
    .B1(_02330_),
    .B2(_09210_),
    .Y(_02333_));
 OA21x2_ASAP7_75t_R _17290_ (.A1(_09288_),
    .A2(_02329_),
    .B(_02333_),
    .Y(_01846_));
 AOI22x1_ASAP7_75t_R _17291_ (.A1(_00262_),
    .A2(_02323_),
    .B1(_02330_),
    .B2(_09212_),
    .Y(_02334_));
 OA21x2_ASAP7_75t_R _17292_ (.A1(_09290_),
    .A2(_02329_),
    .B(_02334_),
    .Y(_01847_));
 AOI22x1_ASAP7_75t_R _17293_ (.A1(_00228_),
    .A2(_02323_),
    .B1(_02330_),
    .B2(_09214_),
    .Y(_02335_));
 OA21x2_ASAP7_75t_R _17294_ (.A1(_09292_),
    .A2(_02329_),
    .B(_02335_),
    .Y(_01848_));
 AOI22x1_ASAP7_75t_R _17295_ (.A1(_00195_),
    .A2(_02323_),
    .B1(_02330_),
    .B2(_09216_),
    .Y(_02336_));
 OA21x2_ASAP7_75t_R _17296_ (.A1(_09294_),
    .A2(_02329_),
    .B(_02336_),
    .Y(_01849_));
 INVx1_ASAP7_75t_R _17297_ (.A(_00161_),
    .Y(_02337_));
 OA222x2_ASAP7_75t_R _17298_ (.A1(_02337_),
    .A2(_02307_),
    .B1(_02308_),
    .B2(_09296_),
    .C1(_02310_),
    .C2(_09219_),
    .Y(_01850_));
 AOI22x1_ASAP7_75t_R _17299_ (.A1(_00128_),
    .A2(_02323_),
    .B1(_02330_),
    .B2(_09220_),
    .Y(_02338_));
 OA21x2_ASAP7_75t_R _17300_ (.A1(_09297_),
    .A2(_02329_),
    .B(_02338_),
    .Y(_01851_));
 NOR2x1_ASAP7_75t_R _17301_ (.A(_01026_),
    .B(_02307_),
    .Y(_02339_));
 AO21x1_ASAP7_75t_R _17302_ (.A1(_09299_),
    .A2(_02307_),
    .B(_02339_),
    .Y(_01852_));
 AND3x1_ASAP7_75t_R _17303_ (.A(_09503_),
    .B(_08750_),
    .C(_09504_),
    .Y(_02340_));
 NOR2x1_ASAP7_75t_R _17304_ (.A(_00094_),
    .B(_02307_),
    .Y(_02341_));
 AO221x1_ASAP7_75t_R _17305_ (.A1(_09223_),
    .A2(_02307_),
    .B1(_02340_),
    .B2(_09302_),
    .C(_02341_),
    .Y(_01853_));
 AND2x2_ASAP7_75t_R _17306_ (.A(_00062_),
    .B(_02312_),
    .Y(_02342_));
 AOI221x1_ASAP7_75t_R _17307_ (.A1(_09226_),
    .A2(_02340_),
    .B1(_02315_),
    .B2(_09304_),
    .C(_02342_),
    .Y(_01854_));
 AOI22x1_ASAP7_75t_R _17308_ (.A1(_00993_),
    .A2(_02312_),
    .B1(_02330_),
    .B2(_09228_),
    .Y(_02343_));
 OA21x2_ASAP7_75t_R _17309_ (.A1(_09306_),
    .A2(_02329_),
    .B(_02343_),
    .Y(_01855_));
 AO21x1_ASAP7_75t_R _17310_ (.A1(_09141_),
    .A2(_09504_),
    .B(_06515_),
    .Y(_02344_));
 OA221x2_ASAP7_75t_R _17311_ (.A1(_09308_),
    .A2(_02313_),
    .B1(_02308_),
    .B2(_09230_),
    .C(_02344_),
    .Y(_01856_));
 NAND2x1_ASAP7_75t_R _17312_ (.A(_00926_),
    .B(_02312_),
    .Y(_02345_));
 OA221x2_ASAP7_75t_R _17313_ (.A1(_09232_),
    .A2(_02313_),
    .B1(_02308_),
    .B2(_09310_),
    .C(_02345_),
    .Y(_01857_));
 AOI22x1_ASAP7_75t_R _17314_ (.A1(_00893_),
    .A2(_02312_),
    .B1(_02330_),
    .B2(_09234_),
    .Y(_02346_));
 OA21x2_ASAP7_75t_R _17315_ (.A1(_09312_),
    .A2(_02329_),
    .B(_02346_),
    .Y(_01858_));
 AO21x1_ASAP7_75t_R _17316_ (.A1(_08750_),
    .A2(_09504_),
    .B(_06232_),
    .Y(_02347_));
 OA21x2_ASAP7_75t_R _17317_ (.A1(_09315_),
    .A2(_02312_),
    .B(_02347_),
    .Y(_02348_));
 OA21x2_ASAP7_75t_R _17318_ (.A1(_09314_),
    .A2(_02329_),
    .B(_02348_),
    .Y(_01859_));
 AOI22x1_ASAP7_75t_R _17319_ (.A1(_00826_),
    .A2(_02312_),
    .B1(_02330_),
    .B2(_09238_),
    .Y(_02349_));
 OA21x2_ASAP7_75t_R _17320_ (.A1(_09318_),
    .A2(_02308_),
    .B(_02349_),
    .Y(_01860_));
 NAND2x1_ASAP7_75t_R _17321_ (.A(_00792_),
    .B(_02312_),
    .Y(_02350_));
 OA21x2_ASAP7_75t_R _17322_ (.A1(_09321_),
    .A2(_02312_),
    .B(_02350_),
    .Y(_02351_));
 OA21x2_ASAP7_75t_R _17323_ (.A1(_09320_),
    .A2(_02308_),
    .B(_02351_),
    .Y(_01861_));
 AND4x2_ASAP7_75t_R _17324_ (.A(_03025_),
    .B(net5),
    .C(net2),
    .D(_06618_),
    .Y(_02352_));
 BUFx12f_ASAP7_75t_R _17325_ (.A(_02352_),
    .Y(_02353_));
 AND2x6_ASAP7_75t_R _17326_ (.A(_08787_),
    .B(_02353_),
    .Y(_02354_));
 NAND2x2_ASAP7_75t_R _17327_ (.A(_09324_),
    .B(_02354_),
    .Y(_02355_));
 BUFx6f_ASAP7_75t_R _17328_ (.A(_02355_),
    .Y(_02356_));
 NAND2x2_ASAP7_75t_R _17329_ (.A(_08115_),
    .B(_02354_),
    .Y(_02357_));
 NAND2x2_ASAP7_75t_R _17330_ (.A(_08787_),
    .B(_02353_),
    .Y(_02358_));
 NAND2x1_ASAP7_75t_R _17331_ (.A(_00028_),
    .B(_02358_),
    .Y(_02359_));
 OA21x2_ASAP7_75t_R _17332_ (.A1(_08111_),
    .A2(_02357_),
    .B(_02359_),
    .Y(_02360_));
 OA21x2_ASAP7_75t_R _17333_ (.A1(_09167_),
    .A2(_02356_),
    .B(_02360_),
    .Y(_01862_));
 BUFx12f_ASAP7_75t_R _17334_ (.A(_02358_),
    .Y(_02361_));
 BUFx6f_ASAP7_75t_R _17335_ (.A(_02353_),
    .Y(_02362_));
 AND3x2_ASAP7_75t_R _17336_ (.A(_09425_),
    .B(_08795_),
    .C(_02362_),
    .Y(_02363_));
 BUFx12_ASAP7_75t_R _17337_ (.A(_02363_),
    .Y(_02364_));
 AOI22x1_ASAP7_75t_R _17338_ (.A1(_00760_),
    .A2(_02361_),
    .B1(_02364_),
    .B2(_09178_),
    .Y(_02365_));
 OA21x2_ASAP7_75t_R _17339_ (.A1(_09251_),
    .A2(_02356_),
    .B(_02365_),
    .Y(_01863_));
 AOI22x1_ASAP7_75t_R _17340_ (.A1(_00727_),
    .A2(_02361_),
    .B1(_02364_),
    .B2(_09180_),
    .Y(_02366_));
 OA21x2_ASAP7_75t_R _17341_ (.A1(_09257_),
    .A2(_02356_),
    .B(_02366_),
    .Y(_01864_));
 OA222x2_ASAP7_75t_R _17342_ (.A1(_05770_),
    .A2(_02354_),
    .B1(_02355_),
    .B2(_09260_),
    .C1(_02357_),
    .C2(_09182_),
    .Y(_01865_));
 OA222x2_ASAP7_75t_R _17343_ (.A1(_05614_),
    .A2(_02354_),
    .B1(_02355_),
    .B2(_09261_),
    .C1(_02357_),
    .C2(_09184_),
    .Y(_01866_));
 AOI22x1_ASAP7_75t_R _17344_ (.A1(_00628_),
    .A2(_02361_),
    .B1(_02364_),
    .B2(_09185_),
    .Y(_02367_));
 OA21x2_ASAP7_75t_R _17345_ (.A1(_09262_),
    .A2(_02356_),
    .B(_02367_),
    .Y(_01867_));
 AOI22x1_ASAP7_75t_R _17346_ (.A1(_00594_),
    .A2(_02361_),
    .B1(_02364_),
    .B2(_09187_),
    .Y(_02368_));
 OA21x2_ASAP7_75t_R _17347_ (.A1(_09264_),
    .A2(_02356_),
    .B(_02368_),
    .Y(_01868_));
 AOI22x1_ASAP7_75t_R _17348_ (.A1(_00561_),
    .A2(_02361_),
    .B1(_02364_),
    .B2(_09189_),
    .Y(_02369_));
 OA21x2_ASAP7_75t_R _17349_ (.A1(_09266_),
    .A2(_02356_),
    .B(_02369_),
    .Y(_01869_));
 BUFx12f_ASAP7_75t_R _17350_ (.A(_02358_),
    .Y(_02370_));
 AOI22x1_ASAP7_75t_R _17351_ (.A1(_00528_),
    .A2(_02370_),
    .B1(_02364_),
    .B2(_09192_),
    .Y(_02371_));
 OA21x2_ASAP7_75t_R _17352_ (.A1(_09268_),
    .A2(_02356_),
    .B(_02371_),
    .Y(_01870_));
 AOI22x1_ASAP7_75t_R _17353_ (.A1(_00495_),
    .A2(_02370_),
    .B1(_02364_),
    .B2(_09194_),
    .Y(_02372_));
 OA21x2_ASAP7_75t_R _17354_ (.A1(_09271_),
    .A2(_02356_),
    .B(_02372_),
    .Y(_01871_));
 AOI22x1_ASAP7_75t_R _17355_ (.A1(_00462_),
    .A2(_02370_),
    .B1(_02364_),
    .B2(_09196_),
    .Y(_02373_));
 OA21x2_ASAP7_75t_R _17356_ (.A1(_09273_),
    .A2(_02356_),
    .B(_02373_),
    .Y(_01872_));
 NAND2x1_ASAP7_75t_R _17357_ (.A(_01060_),
    .B(_02361_),
    .Y(_02374_));
 OA21x2_ASAP7_75t_R _17358_ (.A1(_09275_),
    .A2(_02361_),
    .B(_02374_),
    .Y(_01873_));
 AOI22x1_ASAP7_75t_R _17359_ (.A1(_00429_),
    .A2(_02370_),
    .B1(_02364_),
    .B2(_09199_),
    .Y(_02375_));
 OA21x2_ASAP7_75t_R _17360_ (.A1(_09277_),
    .A2(_02356_),
    .B(_02375_),
    .Y(_01874_));
 BUFx10_ASAP7_75t_R _17361_ (.A(_02358_),
    .Y(_02376_));
 NAND2x1_ASAP7_75t_R _17362_ (.A(_00396_),
    .B(_02376_),
    .Y(_02377_));
 OA221x2_ASAP7_75t_R _17363_ (.A1(_09201_),
    .A2(_02361_),
    .B1(_02355_),
    .B2(_09279_),
    .C(_02377_),
    .Y(_01875_));
 BUFx4f_ASAP7_75t_R _17364_ (.A(_02355_),
    .Y(_02378_));
 BUFx6f_ASAP7_75t_R _17365_ (.A(_02363_),
    .Y(_02379_));
 AOI22x1_ASAP7_75t_R _17366_ (.A1(_00363_),
    .A2(_02370_),
    .B1(_02379_),
    .B2(_09206_),
    .Y(_02380_));
 OA21x2_ASAP7_75t_R _17367_ (.A1(_09282_),
    .A2(_02378_),
    .B(_02380_),
    .Y(_01876_));
 AOI22x1_ASAP7_75t_R _17368_ (.A1(_00329_),
    .A2(_02370_),
    .B1(_02379_),
    .B2(_09208_),
    .Y(_02381_));
 OA21x2_ASAP7_75t_R _17369_ (.A1(_09286_),
    .A2(_02378_),
    .B(_02381_),
    .Y(_01877_));
 AOI22x1_ASAP7_75t_R _17370_ (.A1(_00296_),
    .A2(_02370_),
    .B1(_02379_),
    .B2(_09210_),
    .Y(_02382_));
 OA21x2_ASAP7_75t_R _17371_ (.A1(_09288_),
    .A2(_02378_),
    .B(_02382_),
    .Y(_01878_));
 AOI22x1_ASAP7_75t_R _17372_ (.A1(_00263_),
    .A2(_02370_),
    .B1(_02379_),
    .B2(_09212_),
    .Y(_02383_));
 OA21x2_ASAP7_75t_R _17373_ (.A1(_09290_),
    .A2(_02378_),
    .B(_02383_),
    .Y(_01879_));
 AOI22x1_ASAP7_75t_R _17374_ (.A1(_00229_),
    .A2(_02370_),
    .B1(_02379_),
    .B2(_09214_),
    .Y(_02384_));
 OA21x2_ASAP7_75t_R _17375_ (.A1(_09292_),
    .A2(_02378_),
    .B(_02384_),
    .Y(_01880_));
 AOI22x1_ASAP7_75t_R _17376_ (.A1(_00196_),
    .A2(_02370_),
    .B1(_02379_),
    .B2(_09216_),
    .Y(_02385_));
 OA21x2_ASAP7_75t_R _17377_ (.A1(_09294_),
    .A2(_02378_),
    .B(_02385_),
    .Y(_01881_));
 OA222x2_ASAP7_75t_R _17378_ (.A1(_03995_),
    .A2(_02354_),
    .B1(_02355_),
    .B2(_09296_),
    .C1(_02357_),
    .C2(_09219_),
    .Y(_01882_));
 AOI22x1_ASAP7_75t_R _17379_ (.A1(_00129_),
    .A2(_02376_),
    .B1(_02379_),
    .B2(_09220_),
    .Y(_02386_));
 OA21x2_ASAP7_75t_R _17380_ (.A1(_09297_),
    .A2(_02378_),
    .B(_02386_),
    .Y(_01883_));
 NOR2x1_ASAP7_75t_R _17381_ (.A(_01027_),
    .B(_02354_),
    .Y(_02387_));
 AO21x1_ASAP7_75t_R _17382_ (.A1(_09299_),
    .A2(_02354_),
    .B(_02387_),
    .Y(_01884_));
 AND3x1_ASAP7_75t_R _17383_ (.A(_09503_),
    .B(_08788_),
    .C(_02362_),
    .Y(_02388_));
 NOR2x1_ASAP7_75t_R _17384_ (.A(_00095_),
    .B(_02354_),
    .Y(_02389_));
 AO221x1_ASAP7_75t_R _17385_ (.A1(_09223_),
    .A2(_02354_),
    .B1(_02388_),
    .B2(_09302_),
    .C(_02389_),
    .Y(_01885_));
 AND2x2_ASAP7_75t_R _17386_ (.A(_00063_),
    .B(_02376_),
    .Y(_02390_));
 AOI221x1_ASAP7_75t_R _17387_ (.A1(_09226_),
    .A2(_02388_),
    .B1(_02364_),
    .B2(_09304_),
    .C(_02390_),
    .Y(_01886_));
 AOI22x1_ASAP7_75t_R _17388_ (.A1(_00994_),
    .A2(_02376_),
    .B1(_02379_),
    .B2(_09228_),
    .Y(_02391_));
 OA21x2_ASAP7_75t_R _17389_ (.A1(_09306_),
    .A2(_02378_),
    .B(_02391_),
    .Y(_01887_));
 NAND2x1_ASAP7_75t_R _17390_ (.A(_00961_),
    .B(_02376_),
    .Y(_02392_));
 OA221x2_ASAP7_75t_R _17391_ (.A1(_09308_),
    .A2(_02361_),
    .B1(_02355_),
    .B2(_09230_),
    .C(_02392_),
    .Y(_01888_));
 NAND2x1_ASAP7_75t_R _17392_ (.A(_00927_),
    .B(_02376_),
    .Y(_02393_));
 OA221x2_ASAP7_75t_R _17393_ (.A1(_09232_),
    .A2(_02361_),
    .B1(_02355_),
    .B2(_09310_),
    .C(_02393_),
    .Y(_01889_));
 AOI22x1_ASAP7_75t_R _17394_ (.A1(_00894_),
    .A2(_02376_),
    .B1(_02379_),
    .B2(_09234_),
    .Y(_02394_));
 OA21x2_ASAP7_75t_R _17395_ (.A1(_09312_),
    .A2(_02378_),
    .B(_02394_),
    .Y(_01890_));
 NAND2x1_ASAP7_75t_R _17396_ (.A(_00860_),
    .B(_02358_),
    .Y(_02395_));
 OA21x2_ASAP7_75t_R _17397_ (.A1(_09315_),
    .A2(_02376_),
    .B(_02395_),
    .Y(_02396_));
 OA21x2_ASAP7_75t_R _17398_ (.A1(_09314_),
    .A2(_02378_),
    .B(_02396_),
    .Y(_01891_));
 AOI22x1_ASAP7_75t_R _17399_ (.A1(_00827_),
    .A2(_02376_),
    .B1(_02379_),
    .B2(_09238_),
    .Y(_02397_));
 OA21x2_ASAP7_75t_R _17400_ (.A1(_09318_),
    .A2(_02355_),
    .B(_02397_),
    .Y(_01892_));
 NAND2x1_ASAP7_75t_R _17401_ (.A(_00793_),
    .B(_02358_),
    .Y(_02398_));
 OA21x2_ASAP7_75t_R _17402_ (.A1(_09321_),
    .A2(_02376_),
    .B(_02398_),
    .Y(_02399_));
 OA21x2_ASAP7_75t_R _17403_ (.A1(_09320_),
    .A2(_02355_),
    .B(_02399_),
    .Y(_01893_));
 BUFx4f_ASAP7_75t_R _17404_ (.A(_08092_),
    .Y(_02400_));
 AND2x6_ASAP7_75t_R _17405_ (.A(_08837_),
    .B(_02353_),
    .Y(_02401_));
 NAND2x2_ASAP7_75t_R _17406_ (.A(_09324_),
    .B(_02401_),
    .Y(_02402_));
 BUFx10_ASAP7_75t_R _17407_ (.A(_02402_),
    .Y(_02403_));
 INVx1_ASAP7_75t_R _17408_ (.A(_00029_),
    .Y(_02404_));
 NAND2x2_ASAP7_75t_R _17409_ (.A(_08114_),
    .B(_02401_),
    .Y(_02405_));
 OA22x2_ASAP7_75t_R _17410_ (.A1(_02404_),
    .A2(_02401_),
    .B1(_02405_),
    .B2(_09330_),
    .Y(_02406_));
 OA21x2_ASAP7_75t_R _17411_ (.A1(_02400_),
    .A2(_02403_),
    .B(_02406_),
    .Y(_01894_));
 NAND2x2_ASAP7_75t_R _17412_ (.A(_08838_),
    .B(_02353_),
    .Y(_02407_));
 BUFx12f_ASAP7_75t_R _17413_ (.A(_02407_),
    .Y(_02408_));
 AND3x2_ASAP7_75t_R _17414_ (.A(_09425_),
    .B(_08847_),
    .C(_02362_),
    .Y(_02409_));
 BUFx12f_ASAP7_75t_R _17415_ (.A(_02409_),
    .Y(_02410_));
 BUFx6f_ASAP7_75t_R _17416_ (.A(_08155_),
    .Y(_02411_));
 AOI22x1_ASAP7_75t_R _17417_ (.A1(_00761_),
    .A2(_02408_),
    .B1(_02410_),
    .B2(_02411_),
    .Y(_02412_));
 OA21x2_ASAP7_75t_R _17418_ (.A1(_09251_),
    .A2(_02403_),
    .B(_02412_),
    .Y(_01895_));
 BUFx6f_ASAP7_75t_R _17419_ (.A(_08184_),
    .Y(_02413_));
 AOI22x1_ASAP7_75t_R _17420_ (.A1(_00728_),
    .A2(_02408_),
    .B1(_02410_),
    .B2(_02413_),
    .Y(_02414_));
 OA21x2_ASAP7_75t_R _17421_ (.A1(_09257_),
    .A2(_02403_),
    .B(_02414_),
    .Y(_01896_));
 BUFx3_ASAP7_75t_R _17422_ (.A(_08190_),
    .Y(_02415_));
 OA222x2_ASAP7_75t_R _17423_ (.A1(_05769_),
    .A2(_02401_),
    .B1(_02402_),
    .B2(_09260_),
    .C1(_02405_),
    .C2(_02415_),
    .Y(_01897_));
 BUFx4f_ASAP7_75t_R _17424_ (.A(_08210_),
    .Y(_02416_));
 OA222x2_ASAP7_75t_R _17425_ (.A1(_05613_),
    .A2(_02401_),
    .B1(_02402_),
    .B2(_09261_),
    .C1(_02405_),
    .C2(_02416_),
    .Y(_01898_));
 BUFx6f_ASAP7_75t_R _17426_ (.A(_08242_),
    .Y(_02417_));
 AOI22x1_ASAP7_75t_R _17427_ (.A1(_00629_),
    .A2(_02408_),
    .B1(_02410_),
    .B2(_02417_),
    .Y(_02418_));
 OA21x2_ASAP7_75t_R _17428_ (.A1(_09262_),
    .A2(_02403_),
    .B(_02418_),
    .Y(_01899_));
 BUFx10_ASAP7_75t_R _17429_ (.A(_08258_),
    .Y(_02419_));
 AOI22x1_ASAP7_75t_R _17430_ (.A1(_00595_),
    .A2(_02408_),
    .B1(_02410_),
    .B2(_02419_),
    .Y(_02420_));
 OA21x2_ASAP7_75t_R _17431_ (.A1(_09264_),
    .A2(_02403_),
    .B(_02420_),
    .Y(_01900_));
 BUFx6f_ASAP7_75t_R _17432_ (.A(_08286_),
    .Y(_02421_));
 AOI22x1_ASAP7_75t_R _17433_ (.A1(_00562_),
    .A2(_02408_),
    .B1(_02410_),
    .B2(_02421_),
    .Y(_02422_));
 OA21x2_ASAP7_75t_R _17434_ (.A1(_09266_),
    .A2(_02403_),
    .B(_02422_),
    .Y(_01901_));
 BUFx16f_ASAP7_75t_R _17435_ (.A(_02407_),
    .Y(_02423_));
 BUFx6f_ASAP7_75t_R _17436_ (.A(_08307_),
    .Y(_02424_));
 AOI22x1_ASAP7_75t_R _17437_ (.A1(_00529_),
    .A2(_02423_),
    .B1(_02410_),
    .B2(_02424_),
    .Y(_02425_));
 OA21x2_ASAP7_75t_R _17438_ (.A1(_09268_),
    .A2(_02403_),
    .B(_02425_),
    .Y(_01902_));
 BUFx6f_ASAP7_75t_R _17439_ (.A(_08326_),
    .Y(_02426_));
 AOI22x1_ASAP7_75t_R _17440_ (.A1(_00496_),
    .A2(_02423_),
    .B1(_02410_),
    .B2(_02426_),
    .Y(_02427_));
 OA21x2_ASAP7_75t_R _17441_ (.A1(_09271_),
    .A2(_02403_),
    .B(_02427_),
    .Y(_01903_));
 BUFx6f_ASAP7_75t_R _17442_ (.A(_08347_),
    .Y(_02428_));
 AOI22x1_ASAP7_75t_R _17443_ (.A1(_00463_),
    .A2(_02423_),
    .B1(_02410_),
    .B2(_02428_),
    .Y(_02429_));
 OA21x2_ASAP7_75t_R _17444_ (.A1(_09273_),
    .A2(_02403_),
    .B(_02429_),
    .Y(_01904_));
 NAND2x1_ASAP7_75t_R _17445_ (.A(_01061_),
    .B(_02408_),
    .Y(_02430_));
 OA21x2_ASAP7_75t_R _17446_ (.A1(_09275_),
    .A2(_02408_),
    .B(_02430_),
    .Y(_01905_));
 BUFx6f_ASAP7_75t_R _17447_ (.A(_08381_),
    .Y(_02431_));
 AOI22x1_ASAP7_75t_R _17448_ (.A1(_00430_),
    .A2(_02423_),
    .B1(_02410_),
    .B2(_02431_),
    .Y(_02432_));
 OA21x2_ASAP7_75t_R _17449_ (.A1(_09277_),
    .A2(_02403_),
    .B(_02432_),
    .Y(_01906_));
 BUFx6f_ASAP7_75t_R _17450_ (.A(_08400_),
    .Y(_02433_));
 BUFx6f_ASAP7_75t_R _17451_ (.A(_02407_),
    .Y(_02434_));
 NAND2x1_ASAP7_75t_R _17452_ (.A(_00397_),
    .B(_02434_),
    .Y(_02435_));
 OA221x2_ASAP7_75t_R _17453_ (.A1(_02433_),
    .A2(_02408_),
    .B1(_02402_),
    .B2(_09279_),
    .C(_02435_),
    .Y(_01907_));
 BUFx4f_ASAP7_75t_R _17454_ (.A(_02402_),
    .Y(_02436_));
 BUFx6f_ASAP7_75t_R _17455_ (.A(_02409_),
    .Y(_02437_));
 BUFx6f_ASAP7_75t_R _17456_ (.A(_08419_),
    .Y(_02438_));
 AOI22x1_ASAP7_75t_R _17457_ (.A1(_00364_),
    .A2(_02423_),
    .B1(_02437_),
    .B2(_02438_),
    .Y(_02439_));
 OA21x2_ASAP7_75t_R _17458_ (.A1(_09282_),
    .A2(_02436_),
    .B(_02439_),
    .Y(_01908_));
 BUFx6f_ASAP7_75t_R _17459_ (.A(_08437_),
    .Y(_02440_));
 AOI22x1_ASAP7_75t_R _17460_ (.A1(_00330_),
    .A2(_02423_),
    .B1(_02437_),
    .B2(_02440_),
    .Y(_02441_));
 OA21x2_ASAP7_75t_R _17461_ (.A1(_09286_),
    .A2(_02436_),
    .B(_02441_),
    .Y(_01909_));
 BUFx6f_ASAP7_75t_R _17462_ (.A(_08458_),
    .Y(_02442_));
 AOI22x1_ASAP7_75t_R _17463_ (.A1(_00297_),
    .A2(_02423_),
    .B1(_02437_),
    .B2(_02442_),
    .Y(_02443_));
 OA21x2_ASAP7_75t_R _17464_ (.A1(_09288_),
    .A2(_02436_),
    .B(_02443_),
    .Y(_01910_));
 BUFx6f_ASAP7_75t_R _17465_ (.A(_08476_),
    .Y(_02444_));
 AOI22x1_ASAP7_75t_R _17466_ (.A1(_00264_),
    .A2(_02423_),
    .B1(_02437_),
    .B2(_02444_),
    .Y(_02445_));
 OA21x2_ASAP7_75t_R _17467_ (.A1(_09290_),
    .A2(_02436_),
    .B(_02445_),
    .Y(_01911_));
 BUFx6f_ASAP7_75t_R _17468_ (.A(_08494_),
    .Y(_02446_));
 AOI22x1_ASAP7_75t_R _17469_ (.A1(_00230_),
    .A2(_02423_),
    .B1(_02437_),
    .B2(_02446_),
    .Y(_02447_));
 OA21x2_ASAP7_75t_R _17470_ (.A1(_09292_),
    .A2(_02436_),
    .B(_02447_),
    .Y(_01912_));
 BUFx6f_ASAP7_75t_R _17471_ (.A(_08511_),
    .Y(_02448_));
 AOI22x1_ASAP7_75t_R _17472_ (.A1(_00197_),
    .A2(_02423_),
    .B1(_02437_),
    .B2(_02448_),
    .Y(_02449_));
 OA21x2_ASAP7_75t_R _17473_ (.A1(_09294_),
    .A2(_02436_),
    .B(_02449_),
    .Y(_01913_));
 BUFx4f_ASAP7_75t_R _17474_ (.A(_08517_),
    .Y(_02450_));
 OA222x2_ASAP7_75t_R _17475_ (.A1(_03993_),
    .A2(_02401_),
    .B1(_02402_),
    .B2(_09296_),
    .C1(_02405_),
    .C2(_02450_),
    .Y(_01914_));
 BUFx6f_ASAP7_75t_R _17476_ (.A(_08545_),
    .Y(_02451_));
 AOI22x1_ASAP7_75t_R _17477_ (.A1(_00130_),
    .A2(_02434_),
    .B1(_02437_),
    .B2(_02451_),
    .Y(_02452_));
 OA21x2_ASAP7_75t_R _17478_ (.A1(_09297_),
    .A2(_02436_),
    .B(_02452_),
    .Y(_01915_));
 NOR2x1_ASAP7_75t_R _17479_ (.A(_01028_),
    .B(_02401_),
    .Y(_02453_));
 AO21x1_ASAP7_75t_R _17480_ (.A1(_09299_),
    .A2(_02401_),
    .B(_02453_),
    .Y(_01916_));
 BUFx3_ASAP7_75t_R _17481_ (.A(_08564_),
    .Y(_02454_));
 AND3x1_ASAP7_75t_R _17482_ (.A(_09503_),
    .B(_08873_),
    .C(_02362_),
    .Y(_02455_));
 NOR2x1_ASAP7_75t_R _17483_ (.A(_00096_),
    .B(_02401_),
    .Y(_02456_));
 AO221x1_ASAP7_75t_R _17484_ (.A1(_02454_),
    .A2(_02401_),
    .B1(_02455_),
    .B2(_09302_),
    .C(_02456_),
    .Y(_01917_));
 BUFx6f_ASAP7_75t_R _17485_ (.A(_08590_),
    .Y(_02457_));
 AND2x2_ASAP7_75t_R _17486_ (.A(_00064_),
    .B(_02434_),
    .Y(_02458_));
 AOI221x1_ASAP7_75t_R _17487_ (.A1(_02457_),
    .A2(_02455_),
    .B1(_02410_),
    .B2(_09304_),
    .C(_02458_),
    .Y(_01918_));
 BUFx10_ASAP7_75t_R _17488_ (.A(_08603_),
    .Y(_02459_));
 AOI22x1_ASAP7_75t_R _17489_ (.A1(_00995_),
    .A2(_02434_),
    .B1(_02437_),
    .B2(_02459_),
    .Y(_02460_));
 OA21x2_ASAP7_75t_R _17490_ (.A1(_09306_),
    .A2(_02436_),
    .B(_02460_),
    .Y(_01919_));
 BUFx6f_ASAP7_75t_R _17491_ (.A(_08618_),
    .Y(_02461_));
 NAND2x1_ASAP7_75t_R _17492_ (.A(_00962_),
    .B(_02434_),
    .Y(_02462_));
 OA221x2_ASAP7_75t_R _17493_ (.A1(_09308_),
    .A2(_02408_),
    .B1(_02402_),
    .B2(_02461_),
    .C(_02462_),
    .Y(_01920_));
 BUFx6f_ASAP7_75t_R _17494_ (.A(_08630_),
    .Y(_02463_));
 NAND2x1_ASAP7_75t_R _17495_ (.A(_00928_),
    .B(_02434_),
    .Y(_02464_));
 OA221x2_ASAP7_75t_R _17496_ (.A1(_02463_),
    .A2(_02408_),
    .B1(_02402_),
    .B2(_09310_),
    .C(_02464_),
    .Y(_01921_));
 BUFx10_ASAP7_75t_R _17497_ (.A(_08643_),
    .Y(_02465_));
 AOI22x1_ASAP7_75t_R _17498_ (.A1(_00895_),
    .A2(_02434_),
    .B1(_02437_),
    .B2(_02465_),
    .Y(_02466_));
 OA21x2_ASAP7_75t_R _17499_ (.A1(_09312_),
    .A2(_02436_),
    .B(_02466_),
    .Y(_01922_));
 NAND2x1_ASAP7_75t_R _17500_ (.A(_00861_),
    .B(_02407_),
    .Y(_02467_));
 OA21x2_ASAP7_75t_R _17501_ (.A1(_09315_),
    .A2(_02434_),
    .B(_02467_),
    .Y(_02468_));
 OA21x2_ASAP7_75t_R _17502_ (.A1(_09314_),
    .A2(_02436_),
    .B(_02468_),
    .Y(_01923_));
 BUFx10_ASAP7_75t_R _17503_ (.A(_08669_),
    .Y(_02469_));
 AOI22x1_ASAP7_75t_R _17504_ (.A1(_00828_),
    .A2(_02434_),
    .B1(_02437_),
    .B2(_02469_),
    .Y(_02470_));
 OA21x2_ASAP7_75t_R _17505_ (.A1(_09318_),
    .A2(_02402_),
    .B(_02470_),
    .Y(_01924_));
 NAND2x1_ASAP7_75t_R _17506_ (.A(_00794_),
    .B(_02407_),
    .Y(_02471_));
 OA21x2_ASAP7_75t_R _17507_ (.A1(_09321_),
    .A2(_02434_),
    .B(_02471_),
    .Y(_02472_));
 OA21x2_ASAP7_75t_R _17508_ (.A1(_09320_),
    .A2(_02402_),
    .B(_02472_),
    .Y(_01925_));
 AND2x6_ASAP7_75t_R _17509_ (.A(_08097_),
    .B(_08777_),
    .Y(_02473_));
 NAND2x2_ASAP7_75t_R _17510_ (.A(_09324_),
    .B(_02473_),
    .Y(_02474_));
 BUFx10_ASAP7_75t_R _17511_ (.A(_02474_),
    .Y(_02475_));
 NAND2x2_ASAP7_75t_R _17512_ (.A(_08115_),
    .B(_02473_),
    .Y(_02476_));
 NAND2x2_ASAP7_75t_R _17513_ (.A(_08098_),
    .B(_08777_),
    .Y(_02477_));
 NAND2x1_ASAP7_75t_R _17514_ (.A(_00002_),
    .B(_02477_),
    .Y(_02478_));
 OA21x2_ASAP7_75t_R _17515_ (.A1(_08111_),
    .A2(_02476_),
    .B(_02478_),
    .Y(_02479_));
 OA21x2_ASAP7_75t_R _17516_ (.A1(_02400_),
    .A2(_02475_),
    .B(_02479_),
    .Y(_01926_));
 BUFx4f_ASAP7_75t_R _17517_ (.A(_08143_),
    .Y(_02480_));
 BUFx12f_ASAP7_75t_R _17518_ (.A(_02477_),
    .Y(_02481_));
 AND3x2_ASAP7_75t_R _17519_ (.A(_08117_),
    .B(_08701_),
    .C(_09175_),
    .Y(_02482_));
 BUFx12f_ASAP7_75t_R _17520_ (.A(_02482_),
    .Y(_02483_));
 AOI22x1_ASAP7_75t_R _17521_ (.A1(_00734_),
    .A2(_02481_),
    .B1(_02483_),
    .B2(_02411_),
    .Y(_02484_));
 OA21x2_ASAP7_75t_R _17522_ (.A1(_02480_),
    .A2(_02475_),
    .B(_02484_),
    .Y(_01927_));
 BUFx4f_ASAP7_75t_R _17523_ (.A(_08178_),
    .Y(_02485_));
 AOI22x1_ASAP7_75t_R _17524_ (.A1(_00701_),
    .A2(_02481_),
    .B1(_02483_),
    .B2(_02413_),
    .Y(_02486_));
 OA21x2_ASAP7_75t_R _17525_ (.A1(_02485_),
    .A2(_02475_),
    .B(_02486_),
    .Y(_01928_));
 INVx1_ASAP7_75t_R _17526_ (.A(_00668_),
    .Y(_02487_));
 BUFx3_ASAP7_75t_R _17527_ (.A(_08206_),
    .Y(_02488_));
 OA222x2_ASAP7_75t_R _17528_ (.A1(_02487_),
    .A2(_02473_),
    .B1(_02474_),
    .B2(_02488_),
    .C1(_02476_),
    .C2(_02415_),
    .Y(_01929_));
 INVx1_ASAP7_75t_R _17529_ (.A(_00635_),
    .Y(_02489_));
 BUFx4f_ASAP7_75t_R _17530_ (.A(_08224_),
    .Y(_02490_));
 OA222x2_ASAP7_75t_R _17531_ (.A1(_02489_),
    .A2(_02473_),
    .B1(_02474_),
    .B2(_02490_),
    .C1(_02476_),
    .C2(_02416_),
    .Y(_01930_));
 BUFx4f_ASAP7_75t_R _17532_ (.A(_08240_),
    .Y(_02491_));
 AOI22x1_ASAP7_75t_R _17533_ (.A1(_00602_),
    .A2(_02481_),
    .B1(_02483_),
    .B2(_02417_),
    .Y(_02492_));
 OA21x2_ASAP7_75t_R _17534_ (.A1(_02491_),
    .A2(_02475_),
    .B(_02492_),
    .Y(_01931_));
 BUFx4f_ASAP7_75t_R _17535_ (.A(_08256_),
    .Y(_02493_));
 AOI22x1_ASAP7_75t_R _17536_ (.A1(_00568_),
    .A2(_02481_),
    .B1(_02483_),
    .B2(_02419_),
    .Y(_02494_));
 OA21x2_ASAP7_75t_R _17537_ (.A1(_02493_),
    .A2(_02475_),
    .B(_02494_),
    .Y(_01932_));
 BUFx4f_ASAP7_75t_R _17538_ (.A(_08279_),
    .Y(_02495_));
 AOI22x1_ASAP7_75t_R _17539_ (.A1(_00535_),
    .A2(_02481_),
    .B1(_02483_),
    .B2(_02421_),
    .Y(_02496_));
 OA21x2_ASAP7_75t_R _17540_ (.A1(_02495_),
    .A2(_02475_),
    .B(_02496_),
    .Y(_01933_));
 BUFx4f_ASAP7_75t_R _17541_ (.A(_08301_),
    .Y(_02497_));
 BUFx16f_ASAP7_75t_R _17542_ (.A(_02477_),
    .Y(_02498_));
 AOI22x1_ASAP7_75t_R _17543_ (.A1(_00502_),
    .A2(_02498_),
    .B1(_02483_),
    .B2(_02424_),
    .Y(_02499_));
 OA21x2_ASAP7_75t_R _17544_ (.A1(_02497_),
    .A2(_02475_),
    .B(_02499_),
    .Y(_01934_));
 BUFx3_ASAP7_75t_R _17545_ (.A(_08323_),
    .Y(_02500_));
 AOI22x1_ASAP7_75t_R _17546_ (.A1(_00469_),
    .A2(_02498_),
    .B1(_02483_),
    .B2(_02426_),
    .Y(_02501_));
 OA21x2_ASAP7_75t_R _17547_ (.A1(_02500_),
    .A2(_02475_),
    .B(_02501_),
    .Y(_01935_));
 BUFx4f_ASAP7_75t_R _17548_ (.A(_08344_),
    .Y(_02502_));
 AOI22x1_ASAP7_75t_R _17549_ (.A1(_00436_),
    .A2(_02498_),
    .B1(_02483_),
    .B2(_02428_),
    .Y(_02503_));
 OA21x2_ASAP7_75t_R _17550_ (.A1(_02502_),
    .A2(_02475_),
    .B(_02503_),
    .Y(_01936_));
 BUFx4f_ASAP7_75t_R _17551_ (.A(_08364_),
    .Y(_02504_));
 NAND2x1_ASAP7_75t_R _17552_ (.A(_01034_),
    .B(_02481_),
    .Y(_02505_));
 OA21x2_ASAP7_75t_R _17553_ (.A1(_02504_),
    .A2(_02481_),
    .B(_02505_),
    .Y(_01937_));
 BUFx4f_ASAP7_75t_R _17554_ (.A(_08378_),
    .Y(_02506_));
 AOI22x1_ASAP7_75t_R _17555_ (.A1(_00403_),
    .A2(_02498_),
    .B1(_02483_),
    .B2(_02431_),
    .Y(_02507_));
 OA21x2_ASAP7_75t_R _17556_ (.A1(_02506_),
    .A2(_02475_),
    .B(_02507_),
    .Y(_01938_));
 BUFx6f_ASAP7_75t_R _17557_ (.A(_08396_),
    .Y(_02508_));
 BUFx6f_ASAP7_75t_R _17558_ (.A(_02477_),
    .Y(_02509_));
 NAND2x1_ASAP7_75t_R _17559_ (.A(_00370_),
    .B(_02509_),
    .Y(_02510_));
 OA221x2_ASAP7_75t_R _17560_ (.A1(_02433_),
    .A2(_02481_),
    .B1(_02474_),
    .B2(_02508_),
    .C(_02510_),
    .Y(_01939_));
 BUFx3_ASAP7_75t_R _17561_ (.A(_08415_),
    .Y(_02511_));
 BUFx4f_ASAP7_75t_R _17562_ (.A(_02474_),
    .Y(_02512_));
 BUFx6f_ASAP7_75t_R _17563_ (.A(_02482_),
    .Y(_02513_));
 AOI22x1_ASAP7_75t_R _17564_ (.A1(_00337_),
    .A2(_02498_),
    .B1(_02513_),
    .B2(_02438_),
    .Y(_02514_));
 OA21x2_ASAP7_75t_R _17565_ (.A1(_02511_),
    .A2(_02512_),
    .B(_02514_),
    .Y(_01940_));
 BUFx3_ASAP7_75t_R _17566_ (.A(_08434_),
    .Y(_02515_));
 AOI22x1_ASAP7_75t_R _17567_ (.A1(_00303_),
    .A2(_02498_),
    .B1(_02513_),
    .B2(_02440_),
    .Y(_02516_));
 OA21x2_ASAP7_75t_R _17568_ (.A1(_02515_),
    .A2(_02512_),
    .B(_02516_),
    .Y(_01941_));
 BUFx4f_ASAP7_75t_R _17569_ (.A(_08455_),
    .Y(_02517_));
 AOI22x1_ASAP7_75t_R _17570_ (.A1(_00270_),
    .A2(_02498_),
    .B1(_02513_),
    .B2(_02442_),
    .Y(_02518_));
 OA21x2_ASAP7_75t_R _17571_ (.A1(_02517_),
    .A2(_02512_),
    .B(_02518_),
    .Y(_01942_));
 BUFx4f_ASAP7_75t_R _17572_ (.A(_08472_),
    .Y(_02519_));
 AOI22x1_ASAP7_75t_R _17573_ (.A1(_00237_),
    .A2(_02498_),
    .B1(_02513_),
    .B2(_02444_),
    .Y(_02520_));
 OA21x2_ASAP7_75t_R _17574_ (.A1(_02519_),
    .A2(_02512_),
    .B(_02520_),
    .Y(_01943_));
 BUFx4f_ASAP7_75t_R _17575_ (.A(_08491_),
    .Y(_02521_));
 AOI22x1_ASAP7_75t_R _17576_ (.A1(_00203_),
    .A2(_02498_),
    .B1(_02513_),
    .B2(_02446_),
    .Y(_02522_));
 OA21x2_ASAP7_75t_R _17577_ (.A1(_02521_),
    .A2(_02512_),
    .B(_02522_),
    .Y(_01944_));
 BUFx4f_ASAP7_75t_R _17578_ (.A(_08508_),
    .Y(_02523_));
 AOI22x1_ASAP7_75t_R _17579_ (.A1(_00170_),
    .A2(_02498_),
    .B1(_02513_),
    .B2(_02448_),
    .Y(_02524_));
 OA21x2_ASAP7_75t_R _17580_ (.A1(_02523_),
    .A2(_02512_),
    .B(_02524_),
    .Y(_01945_));
 BUFx4f_ASAP7_75t_R _17581_ (.A(_08531_),
    .Y(_02525_));
 OA222x2_ASAP7_75t_R _17582_ (.A1(_04014_),
    .A2(_02473_),
    .B1(_02474_),
    .B2(_02525_),
    .C1(_02476_),
    .C2(_02450_),
    .Y(_01946_));
 BUFx4f_ASAP7_75t_R _17583_ (.A(_08542_),
    .Y(_02526_));
 AOI22x1_ASAP7_75t_R _17584_ (.A1(_00103_),
    .A2(_02509_),
    .B1(_02513_),
    .B2(_02451_),
    .Y(_02527_));
 OA21x2_ASAP7_75t_R _17585_ (.A1(_02526_),
    .A2(_02512_),
    .B(_02527_),
    .Y(_01947_));
 BUFx6f_ASAP7_75t_R _17586_ (.A(_08560_),
    .Y(_02528_));
 NOR2x1_ASAP7_75t_R _17587_ (.A(_01001_),
    .B(_02473_),
    .Y(_02529_));
 AO21x1_ASAP7_75t_R _17588_ (.A1(_02528_),
    .A2(_02473_),
    .B(_02529_),
    .Y(_01948_));
 AND3x1_ASAP7_75t_R _17589_ (.A(_08145_),
    .B(_08577_),
    .C(_09175_),
    .Y(_02530_));
 BUFx4f_ASAP7_75t_R _17590_ (.A(_08576_),
    .Y(_02531_));
 NOR2x1_ASAP7_75t_R _17591_ (.A(_00069_),
    .B(_02473_),
    .Y(_02532_));
 AO221x1_ASAP7_75t_R _17592_ (.A1(_02454_),
    .A2(_02473_),
    .B1(_02530_),
    .B2(_02531_),
    .C(_02532_),
    .Y(_01949_));
 BUFx6f_ASAP7_75t_R _17593_ (.A(_08594_),
    .Y(_02533_));
 AND2x2_ASAP7_75t_R _17594_ (.A(_00037_),
    .B(_02509_),
    .Y(_02534_));
 AOI221x1_ASAP7_75t_R _17595_ (.A1(_02457_),
    .A2(_02530_),
    .B1(_02483_),
    .B2(_02533_),
    .C(_02534_),
    .Y(_01950_));
 BUFx4f_ASAP7_75t_R _17596_ (.A(_08601_),
    .Y(_02535_));
 AOI22x1_ASAP7_75t_R _17597_ (.A1(_00968_),
    .A2(_02509_),
    .B1(_02513_),
    .B2(_02459_),
    .Y(_02536_));
 OA21x2_ASAP7_75t_R _17598_ (.A1(_02535_),
    .A2(_02512_),
    .B(_02536_),
    .Y(_01951_));
 BUFx6f_ASAP7_75t_R _17599_ (.A(_08609_),
    .Y(_02537_));
 NAND2x1_ASAP7_75t_R _17600_ (.A(_00935_),
    .B(_02509_),
    .Y(_02538_));
 OA221x2_ASAP7_75t_R _17601_ (.A1(_02537_),
    .A2(_02481_),
    .B1(_02474_),
    .B2(_02461_),
    .C(_02538_),
    .Y(_01952_));
 BUFx6f_ASAP7_75t_R _17602_ (.A(_08628_),
    .Y(_02539_));
 NAND2x1_ASAP7_75t_R _17603_ (.A(_00901_),
    .B(_02509_),
    .Y(_02540_));
 OA221x2_ASAP7_75t_R _17604_ (.A1(_02463_),
    .A2(_02481_),
    .B1(_02474_),
    .B2(_02539_),
    .C(_02540_),
    .Y(_01953_));
 BUFx4f_ASAP7_75t_R _17605_ (.A(_08641_),
    .Y(_02541_));
 AOI22x1_ASAP7_75t_R _17606_ (.A1(_00868_),
    .A2(_02509_),
    .B1(_02513_),
    .B2(_02465_),
    .Y(_02542_));
 OA21x2_ASAP7_75t_R _17607_ (.A1(_02541_),
    .A2(_02512_),
    .B(_02542_),
    .Y(_01954_));
 BUFx4f_ASAP7_75t_R _17608_ (.A(_08654_),
    .Y(_02543_));
 BUFx4f_ASAP7_75t_R _17609_ (.A(_08656_),
    .Y(_02544_));
 NAND2x1_ASAP7_75t_R _17610_ (.A(_00834_),
    .B(_02477_),
    .Y(_02545_));
 OA21x2_ASAP7_75t_R _17611_ (.A1(_02544_),
    .A2(_02509_),
    .B(_02545_),
    .Y(_02546_));
 OA21x2_ASAP7_75t_R _17612_ (.A1(_02543_),
    .A2(_02512_),
    .B(_02546_),
    .Y(_01955_));
 BUFx4f_ASAP7_75t_R _17613_ (.A(_08667_),
    .Y(_02547_));
 AOI22x1_ASAP7_75t_R _17614_ (.A1(_00801_),
    .A2(_02509_),
    .B1(_02513_),
    .B2(_02469_),
    .Y(_02548_));
 OA21x2_ASAP7_75t_R _17615_ (.A1(_02547_),
    .A2(_02474_),
    .B(_02548_),
    .Y(_01956_));
 BUFx4f_ASAP7_75t_R _17616_ (.A(_08680_),
    .Y(_02549_));
 BUFx4f_ASAP7_75t_R _17617_ (.A(_08684_),
    .Y(_02550_));
 NAND2x1_ASAP7_75t_R _17618_ (.A(_00767_),
    .B(_02477_),
    .Y(_02551_));
 OA21x2_ASAP7_75t_R _17619_ (.A1(_02550_),
    .A2(_02509_),
    .B(_02551_),
    .Y(_02552_));
 OA21x2_ASAP7_75t_R _17620_ (.A1(_02549_),
    .A2(_02474_),
    .B(_02552_),
    .Y(_01957_));
 AND2x6_ASAP7_75t_R _17621_ (.A(_08097_),
    .B(_02353_),
    .Y(_02553_));
 NAND2x2_ASAP7_75t_R _17622_ (.A(_08606_),
    .B(_02553_),
    .Y(_02554_));
 BUFx10_ASAP7_75t_R _17623_ (.A(_02554_),
    .Y(_02555_));
 NAND2x2_ASAP7_75t_R _17624_ (.A(_08115_),
    .B(_02553_),
    .Y(_02556_));
 NAND2x2_ASAP7_75t_R _17625_ (.A(_08098_),
    .B(_02353_),
    .Y(_02557_));
 NAND2x1_ASAP7_75t_R _17626_ (.A(_00030_),
    .B(_02557_),
    .Y(_02558_));
 OA21x2_ASAP7_75t_R _17627_ (.A1(_08793_),
    .A2(_02556_),
    .B(_02558_),
    .Y(_02559_));
 OA21x2_ASAP7_75t_R _17628_ (.A1(_02400_),
    .A2(_02555_),
    .B(_02559_),
    .Y(_01958_));
 BUFx16f_ASAP7_75t_R _17629_ (.A(_02557_),
    .Y(_02560_));
 AND3x2_ASAP7_75t_R _17630_ (.A(_08117_),
    .B(_08701_),
    .C(_02362_),
    .Y(_02561_));
 BUFx12f_ASAP7_75t_R _17631_ (.A(_02561_),
    .Y(_02562_));
 AOI22x1_ASAP7_75t_R _17632_ (.A1(_00762_),
    .A2(_02560_),
    .B1(_02562_),
    .B2(_02411_),
    .Y(_02563_));
 OA21x2_ASAP7_75t_R _17633_ (.A1(_02480_),
    .A2(_02555_),
    .B(_02563_),
    .Y(_01959_));
 AOI22x1_ASAP7_75t_R _17634_ (.A1(_00729_),
    .A2(_02560_),
    .B1(_02562_),
    .B2(_02413_),
    .Y(_02564_));
 OA21x2_ASAP7_75t_R _17635_ (.A1(_02485_),
    .A2(_02555_),
    .B(_02564_),
    .Y(_01960_));
 OA222x2_ASAP7_75t_R _17636_ (.A1(_05764_),
    .A2(_02553_),
    .B1(_02554_),
    .B2(_02488_),
    .C1(_02556_),
    .C2(_02415_),
    .Y(_01961_));
 INVx1_ASAP7_75t_R _17637_ (.A(_00663_),
    .Y(_02565_));
 OA222x2_ASAP7_75t_R _17638_ (.A1(_02565_),
    .A2(_02553_),
    .B1(_02554_),
    .B2(_02490_),
    .C1(_02556_),
    .C2(_02416_),
    .Y(_01962_));
 AOI22x1_ASAP7_75t_R _17639_ (.A1(_00630_),
    .A2(_02560_),
    .B1(_02562_),
    .B2(_02417_),
    .Y(_02566_));
 OA21x2_ASAP7_75t_R _17640_ (.A1(_02491_),
    .A2(_02555_),
    .B(_02566_),
    .Y(_01963_));
 AOI22x1_ASAP7_75t_R _17641_ (.A1(_00596_),
    .A2(_02560_),
    .B1(_02562_),
    .B2(_02419_),
    .Y(_02567_));
 OA21x2_ASAP7_75t_R _17642_ (.A1(_02493_),
    .A2(_02555_),
    .B(_02567_),
    .Y(_01964_));
 AOI22x1_ASAP7_75t_R _17643_ (.A1(_00563_),
    .A2(_02560_),
    .B1(_02562_),
    .B2(_02421_),
    .Y(_02568_));
 OA21x2_ASAP7_75t_R _17644_ (.A1(_02495_),
    .A2(_02555_),
    .B(_02568_),
    .Y(_01965_));
 BUFx16f_ASAP7_75t_R _17645_ (.A(_02557_),
    .Y(_02569_));
 AOI22x1_ASAP7_75t_R _17646_ (.A1(_00530_),
    .A2(_02569_),
    .B1(_02562_),
    .B2(_02424_),
    .Y(_02570_));
 OA21x2_ASAP7_75t_R _17647_ (.A1(_02497_),
    .A2(_02555_),
    .B(_02570_),
    .Y(_01966_));
 AOI22x1_ASAP7_75t_R _17648_ (.A1(_00497_),
    .A2(_02569_),
    .B1(_02562_),
    .B2(_02426_),
    .Y(_02571_));
 OA21x2_ASAP7_75t_R _17649_ (.A1(_02500_),
    .A2(_02555_),
    .B(_02571_),
    .Y(_01967_));
 AOI22x1_ASAP7_75t_R _17650_ (.A1(_00464_),
    .A2(_02569_),
    .B1(_02562_),
    .B2(_02428_),
    .Y(_02572_));
 OA21x2_ASAP7_75t_R _17651_ (.A1(_02502_),
    .A2(_02555_),
    .B(_02572_),
    .Y(_01968_));
 NAND2x1_ASAP7_75t_R _17652_ (.A(_01062_),
    .B(_02560_),
    .Y(_02573_));
 OA21x2_ASAP7_75t_R _17653_ (.A1(_02504_),
    .A2(_02560_),
    .B(_02573_),
    .Y(_01969_));
 AOI22x1_ASAP7_75t_R _17654_ (.A1(_00431_),
    .A2(_02569_),
    .B1(_02562_),
    .B2(_02431_),
    .Y(_02574_));
 OA21x2_ASAP7_75t_R _17655_ (.A1(_02506_),
    .A2(_02555_),
    .B(_02574_),
    .Y(_01970_));
 BUFx6f_ASAP7_75t_R _17656_ (.A(_02557_),
    .Y(_02575_));
 NAND2x1_ASAP7_75t_R _17657_ (.A(_00398_),
    .B(_02575_),
    .Y(_02576_));
 OA221x2_ASAP7_75t_R _17658_ (.A1(_02433_),
    .A2(_02560_),
    .B1(_02554_),
    .B2(_02508_),
    .C(_02576_),
    .Y(_01971_));
 BUFx4f_ASAP7_75t_R _17659_ (.A(_02554_),
    .Y(_02577_));
 BUFx6f_ASAP7_75t_R _17660_ (.A(_02561_),
    .Y(_02578_));
 AOI22x1_ASAP7_75t_R _17661_ (.A1(_00365_),
    .A2(_02569_),
    .B1(_02578_),
    .B2(_02438_),
    .Y(_02579_));
 OA21x2_ASAP7_75t_R _17662_ (.A1(_02511_),
    .A2(_02577_),
    .B(_02579_),
    .Y(_01972_));
 AOI22x1_ASAP7_75t_R _17663_ (.A1(_00331_),
    .A2(_02569_),
    .B1(_02578_),
    .B2(_02440_),
    .Y(_02580_));
 OA21x2_ASAP7_75t_R _17664_ (.A1(_02515_),
    .A2(_02577_),
    .B(_02580_),
    .Y(_01973_));
 AOI22x1_ASAP7_75t_R _17665_ (.A1(_00298_),
    .A2(_02569_),
    .B1(_02578_),
    .B2(_02442_),
    .Y(_02581_));
 OA21x2_ASAP7_75t_R _17666_ (.A1(_02517_),
    .A2(_02577_),
    .B(_02581_),
    .Y(_01974_));
 AOI22x1_ASAP7_75t_R _17667_ (.A1(_00265_),
    .A2(_02569_),
    .B1(_02578_),
    .B2(_02444_),
    .Y(_02582_));
 OA21x2_ASAP7_75t_R _17668_ (.A1(_02519_),
    .A2(_02577_),
    .B(_02582_),
    .Y(_01975_));
 AOI22x1_ASAP7_75t_R _17669_ (.A1(_00231_),
    .A2(_02569_),
    .B1(_02578_),
    .B2(_02446_),
    .Y(_02583_));
 OA21x2_ASAP7_75t_R _17670_ (.A1(_02521_),
    .A2(_02577_),
    .B(_02583_),
    .Y(_01976_));
 AOI22x1_ASAP7_75t_R _17671_ (.A1(_00198_),
    .A2(_02569_),
    .B1(_02578_),
    .B2(_02448_),
    .Y(_02584_));
 OA21x2_ASAP7_75t_R _17672_ (.A1(_02523_),
    .A2(_02577_),
    .B(_02584_),
    .Y(_01977_));
 INVx1_ASAP7_75t_R _17673_ (.A(_00164_),
    .Y(_02585_));
 OA222x2_ASAP7_75t_R _17674_ (.A1(_02585_),
    .A2(_02553_),
    .B1(_02554_),
    .B2(_02525_),
    .C1(_02556_),
    .C2(_02450_),
    .Y(_01978_));
 AOI22x1_ASAP7_75t_R _17675_ (.A1(_00131_),
    .A2(_02575_),
    .B1(_02578_),
    .B2(_02451_),
    .Y(_02586_));
 OA21x2_ASAP7_75t_R _17676_ (.A1(_02526_),
    .A2(_02577_),
    .B(_02586_),
    .Y(_01979_));
 NOR2x1_ASAP7_75t_R _17677_ (.A(_01029_),
    .B(_02553_),
    .Y(_02587_));
 AO21x1_ASAP7_75t_R _17678_ (.A1(_02528_),
    .A2(_02553_),
    .B(_02587_),
    .Y(_01980_));
 AND3x1_ASAP7_75t_R _17679_ (.A(_08145_),
    .B(_08577_),
    .C(_02362_),
    .Y(_02588_));
 NOR2x1_ASAP7_75t_R _17680_ (.A(_00097_),
    .B(_02553_),
    .Y(_02589_));
 AO221x1_ASAP7_75t_R _17681_ (.A1(_02454_),
    .A2(_02553_),
    .B1(_02588_),
    .B2(_02531_),
    .C(_02589_),
    .Y(_01981_));
 AND2x2_ASAP7_75t_R _17682_ (.A(_00065_),
    .B(_02575_),
    .Y(_02590_));
 AOI221x1_ASAP7_75t_R _17683_ (.A1(_02457_),
    .A2(_02588_),
    .B1(_02562_),
    .B2(_02533_),
    .C(_02590_),
    .Y(_01982_));
 AOI22x1_ASAP7_75t_R _17684_ (.A1(_00996_),
    .A2(_02575_),
    .B1(_02578_),
    .B2(_02459_),
    .Y(_02591_));
 OA21x2_ASAP7_75t_R _17685_ (.A1(_02535_),
    .A2(_02577_),
    .B(_02591_),
    .Y(_01983_));
 NAND2x1_ASAP7_75t_R _17686_ (.A(_00963_),
    .B(_02575_),
    .Y(_02592_));
 OA221x2_ASAP7_75t_R _17687_ (.A1(_02537_),
    .A2(_02560_),
    .B1(_02554_),
    .B2(_02461_),
    .C(_02592_),
    .Y(_01984_));
 NAND2x1_ASAP7_75t_R _17688_ (.A(_00929_),
    .B(_02575_),
    .Y(_02593_));
 OA221x2_ASAP7_75t_R _17689_ (.A1(_02463_),
    .A2(_02560_),
    .B1(_02554_),
    .B2(_02539_),
    .C(_02593_),
    .Y(_01985_));
 AOI22x1_ASAP7_75t_R _17690_ (.A1(_00896_),
    .A2(_02575_),
    .B1(_02578_),
    .B2(_02465_),
    .Y(_02594_));
 OA21x2_ASAP7_75t_R _17691_ (.A1(_02541_),
    .A2(_02577_),
    .B(_02594_),
    .Y(_01986_));
 NAND2x1_ASAP7_75t_R _17692_ (.A(_00862_),
    .B(_02557_),
    .Y(_02595_));
 OA21x2_ASAP7_75t_R _17693_ (.A1(_02544_),
    .A2(_02575_),
    .B(_02595_),
    .Y(_02596_));
 OA21x2_ASAP7_75t_R _17694_ (.A1(_02543_),
    .A2(_02577_),
    .B(_02596_),
    .Y(_01987_));
 AOI22x1_ASAP7_75t_R _17695_ (.A1(_00829_),
    .A2(_02575_),
    .B1(_02578_),
    .B2(_02469_),
    .Y(_02597_));
 OA21x2_ASAP7_75t_R _17696_ (.A1(_02547_),
    .A2(_02554_),
    .B(_02597_),
    .Y(_01988_));
 NAND2x1_ASAP7_75t_R _17697_ (.A(_00795_),
    .B(_02557_),
    .Y(_02598_));
 OA21x2_ASAP7_75t_R _17698_ (.A1(_02550_),
    .A2(_02575_),
    .B(_02598_),
    .Y(_02599_));
 OA21x2_ASAP7_75t_R _17699_ (.A1(_02549_),
    .A2(_02554_),
    .B(_02599_),
    .Y(_01989_));
 AND2x6_ASAP7_75t_R _17700_ (.A(_08689_),
    .B(_02353_),
    .Y(_02600_));
 NAND2x2_ASAP7_75t_R _17701_ (.A(_08606_),
    .B(_02600_),
    .Y(_02601_));
 BUFx10_ASAP7_75t_R _17702_ (.A(_02601_),
    .Y(_02602_));
 NAND2x2_ASAP7_75t_R _17703_ (.A(_08114_),
    .B(_02600_),
    .Y(_02603_));
 OA22x2_ASAP7_75t_R _17704_ (.A1(_03148_),
    .A2(_02600_),
    .B1(_02603_),
    .B2(_09330_),
    .Y(_02604_));
 OA21x2_ASAP7_75t_R _17705_ (.A1(_02400_),
    .A2(_02602_),
    .B(_02604_),
    .Y(_01990_));
 NAND2x2_ASAP7_75t_R _17706_ (.A(_08694_),
    .B(_02362_),
    .Y(_02605_));
 BUFx12f_ASAP7_75t_R _17707_ (.A(_02605_),
    .Y(_02606_));
 AND3x2_ASAP7_75t_R _17708_ (.A(_09425_),
    .B(_08694_),
    .C(_02362_),
    .Y(_02607_));
 BUFx12f_ASAP7_75t_R _17709_ (.A(_02607_),
    .Y(_02608_));
 AOI22x1_ASAP7_75t_R _17710_ (.A1(_00763_),
    .A2(_02606_),
    .B1(_02608_),
    .B2(_02411_),
    .Y(_02609_));
 OA21x2_ASAP7_75t_R _17711_ (.A1(_02480_),
    .A2(_02602_),
    .B(_02609_),
    .Y(_01991_));
 AOI22x1_ASAP7_75t_R _17712_ (.A1(_00730_),
    .A2(_02606_),
    .B1(_02608_),
    .B2(_02413_),
    .Y(_02610_));
 OA21x2_ASAP7_75t_R _17713_ (.A1(_02485_),
    .A2(_02602_),
    .B(_02610_),
    .Y(_01992_));
 OA222x2_ASAP7_75t_R _17714_ (.A1(_05765_),
    .A2(_02600_),
    .B1(_02601_),
    .B2(_02488_),
    .C1(_02603_),
    .C2(_02415_),
    .Y(_01993_));
 INVx1_ASAP7_75t_R _17715_ (.A(_00664_),
    .Y(_02611_));
 OA222x2_ASAP7_75t_R _17716_ (.A1(_02611_),
    .A2(_02600_),
    .B1(_02601_),
    .B2(_02490_),
    .C1(_02603_),
    .C2(_02416_),
    .Y(_01994_));
 AOI22x1_ASAP7_75t_R _17717_ (.A1(_00631_),
    .A2(_02606_),
    .B1(_02608_),
    .B2(_02417_),
    .Y(_02612_));
 OA21x2_ASAP7_75t_R _17718_ (.A1(_02491_),
    .A2(_02602_),
    .B(_02612_),
    .Y(_01995_));
 AOI22x1_ASAP7_75t_R _17719_ (.A1(_00597_),
    .A2(_02606_),
    .B1(_02608_),
    .B2(_02419_),
    .Y(_02613_));
 OA21x2_ASAP7_75t_R _17720_ (.A1(_02493_),
    .A2(_02602_),
    .B(_02613_),
    .Y(_01996_));
 AOI22x1_ASAP7_75t_R _17721_ (.A1(_00564_),
    .A2(_02606_),
    .B1(_02608_),
    .B2(_02421_),
    .Y(_02614_));
 OA21x2_ASAP7_75t_R _17722_ (.A1(_02495_),
    .A2(_02602_),
    .B(_02614_),
    .Y(_01997_));
 BUFx16f_ASAP7_75t_R _17723_ (.A(_02605_),
    .Y(_02615_));
 AOI22x1_ASAP7_75t_R _17724_ (.A1(_00531_),
    .A2(_02615_),
    .B1(_02608_),
    .B2(_02424_),
    .Y(_02616_));
 OA21x2_ASAP7_75t_R _17725_ (.A1(_02497_),
    .A2(_02602_),
    .B(_02616_),
    .Y(_01998_));
 AOI22x1_ASAP7_75t_R _17726_ (.A1(_00498_),
    .A2(_02615_),
    .B1(_02608_),
    .B2(_02426_),
    .Y(_02617_));
 OA21x2_ASAP7_75t_R _17727_ (.A1(_02500_),
    .A2(_02602_),
    .B(_02617_),
    .Y(_01999_));
 AOI22x1_ASAP7_75t_R _17728_ (.A1(_00465_),
    .A2(_02615_),
    .B1(_02608_),
    .B2(_02428_),
    .Y(_02618_));
 OA21x2_ASAP7_75t_R _17729_ (.A1(_02502_),
    .A2(_02602_),
    .B(_02618_),
    .Y(_02000_));
 NAND2x1_ASAP7_75t_R _17730_ (.A(_01063_),
    .B(_02606_),
    .Y(_02619_));
 OA21x2_ASAP7_75t_R _17731_ (.A1(_02504_),
    .A2(_02606_),
    .B(_02619_),
    .Y(_02001_));
 AOI22x1_ASAP7_75t_R _17732_ (.A1(_00432_),
    .A2(_02615_),
    .B1(_02608_),
    .B2(_02431_),
    .Y(_02620_));
 OA21x2_ASAP7_75t_R _17733_ (.A1(_02506_),
    .A2(_02602_),
    .B(_02620_),
    .Y(_02002_));
 BUFx6f_ASAP7_75t_R _17734_ (.A(_02605_),
    .Y(_02621_));
 NAND2x1_ASAP7_75t_R _17735_ (.A(_00399_),
    .B(_02621_),
    .Y(_02622_));
 OA221x2_ASAP7_75t_R _17736_ (.A1(_02433_),
    .A2(_02606_),
    .B1(_02601_),
    .B2(_02508_),
    .C(_02622_),
    .Y(_02003_));
 BUFx4f_ASAP7_75t_R _17737_ (.A(_02601_),
    .Y(_02623_));
 BUFx6f_ASAP7_75t_R _17738_ (.A(_02607_),
    .Y(_02624_));
 AOI22x1_ASAP7_75t_R _17739_ (.A1(_00366_),
    .A2(_02615_),
    .B1(_02624_),
    .B2(_02438_),
    .Y(_02625_));
 OA21x2_ASAP7_75t_R _17740_ (.A1(_02511_),
    .A2(_02623_),
    .B(_02625_),
    .Y(_02004_));
 AOI22x1_ASAP7_75t_R _17741_ (.A1(_00332_),
    .A2(_02615_),
    .B1(_02624_),
    .B2(_02440_),
    .Y(_02626_));
 OA21x2_ASAP7_75t_R _17742_ (.A1(_02515_),
    .A2(_02623_),
    .B(_02626_),
    .Y(_02005_));
 AOI22x1_ASAP7_75t_R _17743_ (.A1(_00299_),
    .A2(_02615_),
    .B1(_02624_),
    .B2(_02442_),
    .Y(_02627_));
 OA21x2_ASAP7_75t_R _17744_ (.A1(_02517_),
    .A2(_02623_),
    .B(_02627_),
    .Y(_02006_));
 AOI22x1_ASAP7_75t_R _17745_ (.A1(_00266_),
    .A2(_02615_),
    .B1(_02624_),
    .B2(_02444_),
    .Y(_02628_));
 OA21x2_ASAP7_75t_R _17746_ (.A1(_02519_),
    .A2(_02623_),
    .B(_02628_),
    .Y(_02007_));
 AOI22x1_ASAP7_75t_R _17747_ (.A1(_00232_),
    .A2(_02615_),
    .B1(_02624_),
    .B2(_02446_),
    .Y(_02629_));
 OA21x2_ASAP7_75t_R _17748_ (.A1(_02521_),
    .A2(_02623_),
    .B(_02629_),
    .Y(_02008_));
 AOI22x1_ASAP7_75t_R _17749_ (.A1(_00199_),
    .A2(_02615_),
    .B1(_02624_),
    .B2(_02448_),
    .Y(_02630_));
 OA21x2_ASAP7_75t_R _17750_ (.A1(_02523_),
    .A2(_02623_),
    .B(_02630_),
    .Y(_02009_));
 INVx1_ASAP7_75t_R _17751_ (.A(_00165_),
    .Y(_02631_));
 OA222x2_ASAP7_75t_R _17752_ (.A1(_02631_),
    .A2(_02600_),
    .B1(_02601_),
    .B2(_02525_),
    .C1(_02603_),
    .C2(_02450_),
    .Y(_02010_));
 AOI22x1_ASAP7_75t_R _17753_ (.A1(_00132_),
    .A2(_02621_),
    .B1(_02624_),
    .B2(_02451_),
    .Y(_02632_));
 OA21x2_ASAP7_75t_R _17754_ (.A1(_02526_),
    .A2(_02623_),
    .B(_02632_),
    .Y(_02011_));
 NOR2x1_ASAP7_75t_R _17755_ (.A(_01030_),
    .B(_02600_),
    .Y(_02633_));
 AO21x1_ASAP7_75t_R _17756_ (.A1(_02528_),
    .A2(_02600_),
    .B(_02633_),
    .Y(_02012_));
 AND3x1_ASAP7_75t_R _17757_ (.A(_09503_),
    .B(_08750_),
    .C(_02362_),
    .Y(_02634_));
 NOR2x1_ASAP7_75t_R _17758_ (.A(_00098_),
    .B(_02600_),
    .Y(_02635_));
 AO221x1_ASAP7_75t_R _17759_ (.A1(_02454_),
    .A2(_02600_),
    .B1(_02634_),
    .B2(_02531_),
    .C(_02635_),
    .Y(_02013_));
 AND2x2_ASAP7_75t_R _17760_ (.A(_00066_),
    .B(_02621_),
    .Y(_02636_));
 AOI221x1_ASAP7_75t_R _17761_ (.A1(_02457_),
    .A2(_02634_),
    .B1(_02608_),
    .B2(_02533_),
    .C(_02636_),
    .Y(_02014_));
 AOI22x1_ASAP7_75t_R _17762_ (.A1(_00997_),
    .A2(_02621_),
    .B1(_02624_),
    .B2(_02459_),
    .Y(_02637_));
 OA21x2_ASAP7_75t_R _17763_ (.A1(_02535_),
    .A2(_02623_),
    .B(_02637_),
    .Y(_02015_));
 NAND2x1_ASAP7_75t_R _17764_ (.A(_00964_),
    .B(_02621_),
    .Y(_02638_));
 OA221x2_ASAP7_75t_R _17765_ (.A1(_02537_),
    .A2(_02606_),
    .B1(_02601_),
    .B2(_02461_),
    .C(_02638_),
    .Y(_02016_));
 NAND2x1_ASAP7_75t_R _17766_ (.A(_00930_),
    .B(_02621_),
    .Y(_02639_));
 OA221x2_ASAP7_75t_R _17767_ (.A1(_02463_),
    .A2(_02606_),
    .B1(_02601_),
    .B2(_02539_),
    .C(_02639_),
    .Y(_02017_));
 AOI22x1_ASAP7_75t_R _17768_ (.A1(_00897_),
    .A2(_02621_),
    .B1(_02624_),
    .B2(_02465_),
    .Y(_02640_));
 OA21x2_ASAP7_75t_R _17769_ (.A1(_02541_),
    .A2(_02623_),
    .B(_02640_),
    .Y(_02018_));
 AO21x1_ASAP7_75t_R _17770_ (.A1(_08749_),
    .A2(_02362_),
    .B(_06230_),
    .Y(_02641_));
 OA21x2_ASAP7_75t_R _17771_ (.A1(_02544_),
    .A2(_02621_),
    .B(_02641_),
    .Y(_02642_));
 OA21x2_ASAP7_75t_R _17772_ (.A1(_02543_),
    .A2(_02623_),
    .B(_02642_),
    .Y(_02019_));
 AOI22x1_ASAP7_75t_R _17773_ (.A1(_00830_),
    .A2(_02621_),
    .B1(_02624_),
    .B2(_02469_),
    .Y(_02643_));
 OA21x2_ASAP7_75t_R _17774_ (.A1(_02547_),
    .A2(_02601_),
    .B(_02643_),
    .Y(_02020_));
 NAND2x1_ASAP7_75t_R _17775_ (.A(_00796_),
    .B(_02605_),
    .Y(_02644_));
 OA21x2_ASAP7_75t_R _17776_ (.A1(_02550_),
    .A2(_02621_),
    .B(_02644_),
    .Y(_02645_));
 OA21x2_ASAP7_75t_R _17777_ (.A1(_02549_),
    .A2(_02601_),
    .B(_02645_),
    .Y(_02021_));
 AND2x6_ASAP7_75t_R _17778_ (.A(_08689_),
    .B(_08777_),
    .Y(_02646_));
 NAND2x2_ASAP7_75t_R _17779_ (.A(_08606_),
    .B(_02646_),
    .Y(_02647_));
 BUFx6f_ASAP7_75t_R _17780_ (.A(_02647_),
    .Y(_02648_));
 NAND2x2_ASAP7_75t_R _17781_ (.A(_08114_),
    .B(_02646_),
    .Y(_02649_));
 OA22x2_ASAP7_75t_R _17782_ (.A1(_03314_),
    .A2(_02646_),
    .B1(_02649_),
    .B2(_09330_),
    .Y(_02650_));
 OA21x2_ASAP7_75t_R _17783_ (.A1(_02400_),
    .A2(_02648_),
    .B(_02650_),
    .Y(_02022_));
 NAND2x2_ASAP7_75t_R _17784_ (.A(_08694_),
    .B(_08777_),
    .Y(_02651_));
 BUFx6f_ASAP7_75t_R _17785_ (.A(_02651_),
    .Y(_02652_));
 BUFx12f_ASAP7_75t_R _17786_ (.A(_02652_),
    .Y(_02653_));
 AND3x2_ASAP7_75t_R _17787_ (.A(_09425_),
    .B(_08694_),
    .C(_08777_),
    .Y(_02654_));
 BUFx12f_ASAP7_75t_R _17788_ (.A(_02654_),
    .Y(_02655_));
 AOI22x1_ASAP7_75t_R _17789_ (.A1(_00735_),
    .A2(_02653_),
    .B1(_02655_),
    .B2(_02411_),
    .Y(_02656_));
 OA21x2_ASAP7_75t_R _17790_ (.A1(_02480_),
    .A2(_02648_),
    .B(_02656_),
    .Y(_02023_));
 AOI22x1_ASAP7_75t_R _17791_ (.A1(_00702_),
    .A2(_02653_),
    .B1(_02655_),
    .B2(_02413_),
    .Y(_02657_));
 OA21x2_ASAP7_75t_R _17792_ (.A1(_02485_),
    .A2(_02648_),
    .B(_02657_),
    .Y(_02024_));
 INVx1_ASAP7_75t_R _17793_ (.A(_00669_),
    .Y(_02658_));
 OA222x2_ASAP7_75t_R _17794_ (.A1(_02658_),
    .A2(_02646_),
    .B1(_02647_),
    .B2(_02488_),
    .C1(_02649_),
    .C2(_02415_),
    .Y(_02025_));
 INVx1_ASAP7_75t_R _17795_ (.A(_00636_),
    .Y(_02659_));
 OA222x2_ASAP7_75t_R _17796_ (.A1(_02659_),
    .A2(_02646_),
    .B1(_02647_),
    .B2(_02490_),
    .C1(_02649_),
    .C2(_02416_),
    .Y(_02026_));
 AOI22x1_ASAP7_75t_R _17797_ (.A1(_00603_),
    .A2(_02653_),
    .B1(_02655_),
    .B2(_02417_),
    .Y(_02660_));
 OA21x2_ASAP7_75t_R _17798_ (.A1(_02491_),
    .A2(_02648_),
    .B(_02660_),
    .Y(_02027_));
 AOI22x1_ASAP7_75t_R _17799_ (.A1(_00569_),
    .A2(_02653_),
    .B1(_02655_),
    .B2(_02419_),
    .Y(_02661_));
 OA21x2_ASAP7_75t_R _17800_ (.A1(_02493_),
    .A2(_02648_),
    .B(_02661_),
    .Y(_02028_));
 AOI22x1_ASAP7_75t_R _17801_ (.A1(_00536_),
    .A2(_02653_),
    .B1(_02655_),
    .B2(_02421_),
    .Y(_02662_));
 OA21x2_ASAP7_75t_R _17802_ (.A1(_02495_),
    .A2(_02648_),
    .B(_02662_),
    .Y(_02029_));
 BUFx12f_ASAP7_75t_R _17803_ (.A(_02651_),
    .Y(_02663_));
 AOI22x1_ASAP7_75t_R _17804_ (.A1(_00503_),
    .A2(_02663_),
    .B1(_02655_),
    .B2(_02424_),
    .Y(_02664_));
 OA21x2_ASAP7_75t_R _17805_ (.A1(_02497_),
    .A2(_02648_),
    .B(_02664_),
    .Y(_02030_));
 AOI22x1_ASAP7_75t_R _17806_ (.A1(_00470_),
    .A2(_02663_),
    .B1(_02655_),
    .B2(_02426_),
    .Y(_02665_));
 OA21x2_ASAP7_75t_R _17807_ (.A1(_02500_),
    .A2(_02648_),
    .B(_02665_),
    .Y(_02031_));
 AOI22x1_ASAP7_75t_R _17808_ (.A1(_00437_),
    .A2(_02663_),
    .B1(_02655_),
    .B2(_02428_),
    .Y(_02666_));
 OA21x2_ASAP7_75t_R _17809_ (.A1(_02502_),
    .A2(_02648_),
    .B(_02666_),
    .Y(_02032_));
 AO21x1_ASAP7_75t_R _17810_ (.A1(_09141_),
    .A2(_09175_),
    .B(_06804_),
    .Y(_02667_));
 OA21x2_ASAP7_75t_R _17811_ (.A1(_02504_),
    .A2(_02653_),
    .B(_02667_),
    .Y(_02033_));
 AOI22x1_ASAP7_75t_R _17812_ (.A1(_00404_),
    .A2(_02663_),
    .B1(_02655_),
    .B2(_02431_),
    .Y(_02668_));
 OA21x2_ASAP7_75t_R _17813_ (.A1(_02506_),
    .A2(_02648_),
    .B(_02668_),
    .Y(_02034_));
 AO21x1_ASAP7_75t_R _17814_ (.A1(_09141_),
    .A2(_09175_),
    .B(_04773_),
    .Y(_02669_));
 OA221x2_ASAP7_75t_R _17815_ (.A1(_02433_),
    .A2(_02653_),
    .B1(_02647_),
    .B2(_02508_),
    .C(_02669_),
    .Y(_02035_));
 BUFx4f_ASAP7_75t_R _17816_ (.A(_02647_),
    .Y(_02670_));
 BUFx6f_ASAP7_75t_R _17817_ (.A(_02654_),
    .Y(_02671_));
 AOI22x1_ASAP7_75t_R _17818_ (.A1(_00338_),
    .A2(_02663_),
    .B1(_02671_),
    .B2(_02438_),
    .Y(_02672_));
 OA21x2_ASAP7_75t_R _17819_ (.A1(_02511_),
    .A2(_02670_),
    .B(_02672_),
    .Y(_02036_));
 AOI22x1_ASAP7_75t_R _17820_ (.A1(_00304_),
    .A2(_02663_),
    .B1(_02671_),
    .B2(_02440_),
    .Y(_02673_));
 OA21x2_ASAP7_75t_R _17821_ (.A1(_02515_),
    .A2(_02670_),
    .B(_02673_),
    .Y(_02037_));
 AOI22x1_ASAP7_75t_R _17822_ (.A1(_00271_),
    .A2(_02663_),
    .B1(_02671_),
    .B2(_02442_),
    .Y(_02674_));
 OA21x2_ASAP7_75t_R _17823_ (.A1(_02517_),
    .A2(_02670_),
    .B(_02674_),
    .Y(_02038_));
 AOI22x1_ASAP7_75t_R _17824_ (.A1(_00238_),
    .A2(_02663_),
    .B1(_02671_),
    .B2(_02444_),
    .Y(_02675_));
 OA21x2_ASAP7_75t_R _17825_ (.A1(_02519_),
    .A2(_02670_),
    .B(_02675_),
    .Y(_02039_));
 AOI22x1_ASAP7_75t_R _17826_ (.A1(_00204_),
    .A2(_02663_),
    .B1(_02671_),
    .B2(_02446_),
    .Y(_02676_));
 OA21x2_ASAP7_75t_R _17827_ (.A1(_02521_),
    .A2(_02670_),
    .B(_02676_),
    .Y(_02040_));
 AOI22x1_ASAP7_75t_R _17828_ (.A1(_00171_),
    .A2(_02663_),
    .B1(_02671_),
    .B2(_02448_),
    .Y(_02677_));
 OA21x2_ASAP7_75t_R _17829_ (.A1(_02523_),
    .A2(_02670_),
    .B(_02677_),
    .Y(_02041_));
 OA222x2_ASAP7_75t_R _17830_ (.A1(_04016_),
    .A2(_02646_),
    .B1(_02647_),
    .B2(_02525_),
    .C1(_02649_),
    .C2(_02450_),
    .Y(_02042_));
 AOI22x1_ASAP7_75t_R _17831_ (.A1(_00104_),
    .A2(_02652_),
    .B1(_02671_),
    .B2(_02451_),
    .Y(_02678_));
 OA21x2_ASAP7_75t_R _17832_ (.A1(_02526_),
    .A2(_02670_),
    .B(_02678_),
    .Y(_02043_));
 NOR2x1_ASAP7_75t_R _17833_ (.A(_01002_),
    .B(_02646_),
    .Y(_02679_));
 AO21x1_ASAP7_75t_R _17834_ (.A1(_02528_),
    .A2(_02646_),
    .B(_02679_),
    .Y(_02044_));
 INVx1_ASAP7_75t_R _17835_ (.A(_00070_),
    .Y(_02680_));
 AND3x1_ASAP7_75t_R _17836_ (.A(_09503_),
    .B(_08750_),
    .C(_09175_),
    .Y(_02681_));
 AND2x2_ASAP7_75t_R _17837_ (.A(_02454_),
    .B(_02646_),
    .Y(_02682_));
 AO221x1_ASAP7_75t_R _17838_ (.A1(_02680_),
    .A2(_02653_),
    .B1(_02681_),
    .B2(_02531_),
    .C(_02682_),
    .Y(_02045_));
 AND2x2_ASAP7_75t_R _17839_ (.A(_00038_),
    .B(_02652_),
    .Y(_02683_));
 AOI221x1_ASAP7_75t_R _17840_ (.A1(_02457_),
    .A2(_02681_),
    .B1(_02655_),
    .B2(_02533_),
    .C(_02683_),
    .Y(_02046_));
 AOI22x1_ASAP7_75t_R _17841_ (.A1(_00969_),
    .A2(_02652_),
    .B1(_02671_),
    .B2(_02459_),
    .Y(_02684_));
 OA21x2_ASAP7_75t_R _17842_ (.A1(_02535_),
    .A2(_02670_),
    .B(_02684_),
    .Y(_02047_));
 NAND2x1_ASAP7_75t_R _17843_ (.A(_00936_),
    .B(_02652_),
    .Y(_02685_));
 OA221x2_ASAP7_75t_R _17844_ (.A1(_02537_),
    .A2(_02653_),
    .B1(_02647_),
    .B2(_02461_),
    .C(_02685_),
    .Y(_02048_));
 AO21x1_ASAP7_75t_R _17845_ (.A1(_09141_),
    .A2(_09175_),
    .B(_06376_),
    .Y(_02686_));
 OA221x2_ASAP7_75t_R _17846_ (.A1(_02463_),
    .A2(_02653_),
    .B1(_02647_),
    .B2(_02539_),
    .C(_02686_),
    .Y(_02049_));
 AOI22x1_ASAP7_75t_R _17847_ (.A1(_00869_),
    .A2(_02652_),
    .B1(_02671_),
    .B2(_02465_),
    .Y(_02687_));
 OA21x2_ASAP7_75t_R _17848_ (.A1(_02541_),
    .A2(_02670_),
    .B(_02687_),
    .Y(_02050_));
 NAND2x1_ASAP7_75t_R _17849_ (.A(_00835_),
    .B(_02652_),
    .Y(_02688_));
 OA21x2_ASAP7_75t_R _17850_ (.A1(_02544_),
    .A2(_02652_),
    .B(_02688_),
    .Y(_02689_));
 OA21x2_ASAP7_75t_R _17851_ (.A1(_02543_),
    .A2(_02670_),
    .B(_02689_),
    .Y(_02051_));
 AOI22x1_ASAP7_75t_R _17852_ (.A1(_00802_),
    .A2(_02652_),
    .B1(_02671_),
    .B2(_02469_),
    .Y(_02690_));
 OA21x2_ASAP7_75t_R _17853_ (.A1(_02547_),
    .A2(_02647_),
    .B(_02690_),
    .Y(_02052_));
 AO21x1_ASAP7_75t_R _17854_ (.A1(_08749_),
    .A2(_09175_),
    .B(_06014_),
    .Y(_02691_));
 OA21x2_ASAP7_75t_R _17855_ (.A1(_02550_),
    .A2(_02652_),
    .B(_02691_),
    .Y(_02692_));
 OA21x2_ASAP7_75t_R _17856_ (.A1(_02549_),
    .A2(_02647_),
    .B(_02692_),
    .Y(_02053_));
 NOR2x2_ASAP7_75t_R _17857_ (.A(_08100_),
    .B(_08776_),
    .Y(_02693_));
 AND2x6_ASAP7_75t_R _17858_ (.A(_08787_),
    .B(_02693_),
    .Y(_02694_));
 NAND2x2_ASAP7_75t_R _17859_ (.A(_08606_),
    .B(_02694_),
    .Y(_02695_));
 BUFx6f_ASAP7_75t_R _17860_ (.A(_02695_),
    .Y(_02696_));
 INVx1_ASAP7_75t_R _17861_ (.A(_00004_),
    .Y(_02697_));
 NAND2x2_ASAP7_75t_R _17862_ (.A(_08114_),
    .B(_02694_),
    .Y(_02698_));
 OA22x2_ASAP7_75t_R _17863_ (.A1(_02697_),
    .A2(_02694_),
    .B1(_02698_),
    .B2(_09330_),
    .Y(_02699_));
 OA21x2_ASAP7_75t_R _17864_ (.A1(_02400_),
    .A2(_02696_),
    .B(_02699_),
    .Y(_02054_));
 BUFx4f_ASAP7_75t_R _17865_ (.A(_02693_),
    .Y(_02700_));
 NAND2x2_ASAP7_75t_R _17866_ (.A(_08795_),
    .B(_02700_),
    .Y(_02701_));
 BUFx12f_ASAP7_75t_R _17867_ (.A(_02701_),
    .Y(_02702_));
 AND3x2_ASAP7_75t_R _17868_ (.A(_09425_),
    .B(_08795_),
    .C(_02700_),
    .Y(_02703_));
 BUFx12f_ASAP7_75t_R _17869_ (.A(_02703_),
    .Y(_02704_));
 AOI22x1_ASAP7_75t_R _17870_ (.A1(_00736_),
    .A2(_02702_),
    .B1(_02704_),
    .B2(_02411_),
    .Y(_02705_));
 OA21x2_ASAP7_75t_R _17871_ (.A1(_02480_),
    .A2(_02696_),
    .B(_02705_),
    .Y(_02055_));
 AOI22x1_ASAP7_75t_R _17872_ (.A1(_00703_),
    .A2(_02702_),
    .B1(_02704_),
    .B2(_02413_),
    .Y(_02706_));
 OA21x2_ASAP7_75t_R _17873_ (.A1(_02485_),
    .A2(_02696_),
    .B(_02706_),
    .Y(_02056_));
 OA222x2_ASAP7_75t_R _17874_ (.A1(_05722_),
    .A2(_02694_),
    .B1(_02695_),
    .B2(_02488_),
    .C1(_02698_),
    .C2(_02415_),
    .Y(_02057_));
 OA222x2_ASAP7_75t_R _17875_ (.A1(_05642_),
    .A2(_02694_),
    .B1(_02695_),
    .B2(_02490_),
    .C1(_02698_),
    .C2(_02416_),
    .Y(_02058_));
 AOI22x1_ASAP7_75t_R _17876_ (.A1(_00604_),
    .A2(_02702_),
    .B1(_02704_),
    .B2(_02417_),
    .Y(_02707_));
 OA21x2_ASAP7_75t_R _17877_ (.A1(_02491_),
    .A2(_02696_),
    .B(_02707_),
    .Y(_02059_));
 AOI22x1_ASAP7_75t_R _17878_ (.A1(_00570_),
    .A2(_02702_),
    .B1(_02704_),
    .B2(_02419_),
    .Y(_02708_));
 OA21x2_ASAP7_75t_R _17879_ (.A1(_02493_),
    .A2(_02696_),
    .B(_02708_),
    .Y(_02060_));
 BUFx12f_ASAP7_75t_R _17880_ (.A(_02701_),
    .Y(_02709_));
 AOI22x1_ASAP7_75t_R _17881_ (.A1(_00537_),
    .A2(_02709_),
    .B1(_02704_),
    .B2(_02421_),
    .Y(_02710_));
 OA21x2_ASAP7_75t_R _17882_ (.A1(_02495_),
    .A2(_02696_),
    .B(_02710_),
    .Y(_02061_));
 AOI22x1_ASAP7_75t_R _17883_ (.A1(_00504_),
    .A2(_02709_),
    .B1(_02704_),
    .B2(_02424_),
    .Y(_02711_));
 OA21x2_ASAP7_75t_R _17884_ (.A1(_02497_),
    .A2(_02696_),
    .B(_02711_),
    .Y(_02062_));
 AOI22x1_ASAP7_75t_R _17885_ (.A1(_00471_),
    .A2(_02709_),
    .B1(_02704_),
    .B2(_02426_),
    .Y(_02712_));
 OA21x2_ASAP7_75t_R _17886_ (.A1(_02500_),
    .A2(_02696_),
    .B(_02712_),
    .Y(_02063_));
 AOI22x1_ASAP7_75t_R _17887_ (.A1(_00438_),
    .A2(_02709_),
    .B1(_02704_),
    .B2(_02428_),
    .Y(_02713_));
 OA21x2_ASAP7_75t_R _17888_ (.A1(_02502_),
    .A2(_02696_),
    .B(_02713_),
    .Y(_02064_));
 NAND2x1_ASAP7_75t_R _17889_ (.A(_01036_),
    .B(_02702_),
    .Y(_02714_));
 OA21x2_ASAP7_75t_R _17890_ (.A1(_02504_),
    .A2(_02702_),
    .B(_02714_),
    .Y(_02065_));
 AOI22x1_ASAP7_75t_R _17891_ (.A1(_00405_),
    .A2(_02709_),
    .B1(_02704_),
    .B2(_02431_),
    .Y(_02715_));
 OA21x2_ASAP7_75t_R _17892_ (.A1(_02506_),
    .A2(_02696_),
    .B(_02715_),
    .Y(_02066_));
 BUFx6f_ASAP7_75t_R _17893_ (.A(_02701_),
    .Y(_02716_));
 NAND2x1_ASAP7_75t_R _17894_ (.A(_00372_),
    .B(_02716_),
    .Y(_02717_));
 OA221x2_ASAP7_75t_R _17895_ (.A1(_02433_),
    .A2(_02702_),
    .B1(_02695_),
    .B2(_02508_),
    .C(_02717_),
    .Y(_02067_));
 BUFx4f_ASAP7_75t_R _17896_ (.A(_02695_),
    .Y(_02718_));
 BUFx6f_ASAP7_75t_R _17897_ (.A(_02703_),
    .Y(_02719_));
 AOI22x1_ASAP7_75t_R _17898_ (.A1(_00339_),
    .A2(_02709_),
    .B1(_02719_),
    .B2(_02438_),
    .Y(_02720_));
 OA21x2_ASAP7_75t_R _17899_ (.A1(_02511_),
    .A2(_02718_),
    .B(_02720_),
    .Y(_02068_));
 AOI22x1_ASAP7_75t_R _17900_ (.A1(_00305_),
    .A2(_02709_),
    .B1(_02719_),
    .B2(_02440_),
    .Y(_02721_));
 OA21x2_ASAP7_75t_R _17901_ (.A1(_02515_),
    .A2(_02718_),
    .B(_02721_),
    .Y(_02069_));
 AOI22x1_ASAP7_75t_R _17902_ (.A1(_00272_),
    .A2(_02709_),
    .B1(_02719_),
    .B2(_02442_),
    .Y(_02722_));
 OA21x2_ASAP7_75t_R _17903_ (.A1(_02517_),
    .A2(_02718_),
    .B(_02722_),
    .Y(_02070_));
 AOI22x1_ASAP7_75t_R _17904_ (.A1(_00239_),
    .A2(_02709_),
    .B1(_02719_),
    .B2(_02444_),
    .Y(_02723_));
 OA21x2_ASAP7_75t_R _17905_ (.A1(_02519_),
    .A2(_02718_),
    .B(_02723_),
    .Y(_02071_));
 AOI22x1_ASAP7_75t_R _17906_ (.A1(_00205_),
    .A2(_02709_),
    .B1(_02719_),
    .B2(_02446_),
    .Y(_02724_));
 OA21x2_ASAP7_75t_R _17907_ (.A1(_02521_),
    .A2(_02718_),
    .B(_02724_),
    .Y(_02072_));
 AOI22x1_ASAP7_75t_R _17908_ (.A1(_00172_),
    .A2(_02716_),
    .B1(_02719_),
    .B2(_02448_),
    .Y(_02725_));
 OA21x2_ASAP7_75t_R _17909_ (.A1(_02523_),
    .A2(_02718_),
    .B(_02725_),
    .Y(_02073_));
 OA222x2_ASAP7_75t_R _17910_ (.A1(_04008_),
    .A2(_02694_),
    .B1(_02695_),
    .B2(_02525_),
    .C1(_02698_),
    .C2(_02450_),
    .Y(_02074_));
 AOI22x1_ASAP7_75t_R _17911_ (.A1(_00105_),
    .A2(_02716_),
    .B1(_02719_),
    .B2(_02451_),
    .Y(_02726_));
 OA21x2_ASAP7_75t_R _17912_ (.A1(_02526_),
    .A2(_02718_),
    .B(_02726_),
    .Y(_02075_));
 NOR2x1_ASAP7_75t_R _17913_ (.A(_01003_),
    .B(_02694_),
    .Y(_02727_));
 AO21x1_ASAP7_75t_R _17914_ (.A1(_02528_),
    .A2(_02694_),
    .B(_02727_),
    .Y(_02076_));
 AND3x2_ASAP7_75t_R _17915_ (.A(_09503_),
    .B(_08788_),
    .C(_02700_),
    .Y(_02728_));
 AND2x2_ASAP7_75t_R _17916_ (.A(_08564_),
    .B(_02694_),
    .Y(_02729_));
 AO221x1_ASAP7_75t_R _17917_ (.A1(_03758_),
    .A2(_02702_),
    .B1(_02728_),
    .B2(_02531_),
    .C(_02729_),
    .Y(_02077_));
 AND2x2_ASAP7_75t_R _17918_ (.A(_00039_),
    .B(_02701_),
    .Y(_02730_));
 AOI221x1_ASAP7_75t_R _17919_ (.A1(_02457_),
    .A2(_02728_),
    .B1(_02704_),
    .B2(_02533_),
    .C(_02730_),
    .Y(_02078_));
 AOI22x1_ASAP7_75t_R _17920_ (.A1(_00970_),
    .A2(_02716_),
    .B1(_02719_),
    .B2(_02459_),
    .Y(_02731_));
 OA21x2_ASAP7_75t_R _17921_ (.A1(_02535_),
    .A2(_02718_),
    .B(_02731_),
    .Y(_02079_));
 NAND2x1_ASAP7_75t_R _17922_ (.A(_00937_),
    .B(_02716_),
    .Y(_02732_));
 OA221x2_ASAP7_75t_R _17923_ (.A1(_02537_),
    .A2(_02702_),
    .B1(_02695_),
    .B2(_02461_),
    .C(_02732_),
    .Y(_02080_));
 NAND2x1_ASAP7_75t_R _17924_ (.A(_00903_),
    .B(_02716_),
    .Y(_02733_));
 OA221x2_ASAP7_75t_R _17925_ (.A1(_02463_),
    .A2(_02702_),
    .B1(_02695_),
    .B2(_02539_),
    .C(_02733_),
    .Y(_02081_));
 AOI22x1_ASAP7_75t_R _17926_ (.A1(_00870_),
    .A2(_02716_),
    .B1(_02719_),
    .B2(_02465_),
    .Y(_02734_));
 OA21x2_ASAP7_75t_R _17927_ (.A1(_02541_),
    .A2(_02718_),
    .B(_02734_),
    .Y(_02082_));
 NAND2x1_ASAP7_75t_R _17928_ (.A(_00836_),
    .B(_02701_),
    .Y(_02735_));
 OA21x2_ASAP7_75t_R _17929_ (.A1(_02544_),
    .A2(_02716_),
    .B(_02735_),
    .Y(_02736_));
 OA21x2_ASAP7_75t_R _17930_ (.A1(_02543_),
    .A2(_02718_),
    .B(_02736_),
    .Y(_02083_));
 AOI22x1_ASAP7_75t_R _17931_ (.A1(_00803_),
    .A2(_02716_),
    .B1(_02719_),
    .B2(_02469_),
    .Y(_02737_));
 OA21x2_ASAP7_75t_R _17932_ (.A1(_02547_),
    .A2(_02695_),
    .B(_02737_),
    .Y(_02084_));
 NAND2x1_ASAP7_75t_R _17933_ (.A(_00769_),
    .B(_02701_),
    .Y(_02738_));
 OA21x2_ASAP7_75t_R _17934_ (.A1(_02550_),
    .A2(_02716_),
    .B(_02738_),
    .Y(_02739_));
 OA21x2_ASAP7_75t_R _17935_ (.A1(_02549_),
    .A2(_02695_),
    .B(_02739_),
    .Y(_02085_));
 AND2x6_ASAP7_75t_R _17936_ (.A(_08838_),
    .B(_02693_),
    .Y(_02740_));
 NAND2x2_ASAP7_75t_R _17937_ (.A(_08606_),
    .B(_02740_),
    .Y(_02741_));
 BUFx6f_ASAP7_75t_R _17938_ (.A(_02741_),
    .Y(_02742_));
 NAND2x2_ASAP7_75t_R _17939_ (.A(_08937_),
    .B(_02740_),
    .Y(_02743_));
 NAND2x2_ASAP7_75t_R _17940_ (.A(_08838_),
    .B(_02693_),
    .Y(_02744_));
 BUFx6f_ASAP7_75t_R _17941_ (.A(_02744_),
    .Y(_02745_));
 NAND2x1_ASAP7_75t_R _17942_ (.A(_00005_),
    .B(_02745_),
    .Y(_02746_));
 OA21x2_ASAP7_75t_R _17943_ (.A1(_08793_),
    .A2(_02743_),
    .B(_02746_),
    .Y(_02747_));
 OA21x2_ASAP7_75t_R _17944_ (.A1(_02400_),
    .A2(_02742_),
    .B(_02747_),
    .Y(_02086_));
 BUFx12f_ASAP7_75t_R _17945_ (.A(_02744_),
    .Y(_02748_));
 AND3x2_ASAP7_75t_R _17946_ (.A(_09425_),
    .B(_08847_),
    .C(_02700_),
    .Y(_02749_));
 BUFx12_ASAP7_75t_R _17947_ (.A(_02749_),
    .Y(_02750_));
 AOI22x1_ASAP7_75t_R _17948_ (.A1(_00737_),
    .A2(_02748_),
    .B1(_02750_),
    .B2(_02411_),
    .Y(_02751_));
 OA21x2_ASAP7_75t_R _17949_ (.A1(_02480_),
    .A2(_02742_),
    .B(_02751_),
    .Y(_02087_));
 AOI22x1_ASAP7_75t_R _17950_ (.A1(_00704_),
    .A2(_02748_),
    .B1(_02750_),
    .B2(_02413_),
    .Y(_02752_));
 OA21x2_ASAP7_75t_R _17951_ (.A1(_02485_),
    .A2(_02742_),
    .B(_02752_),
    .Y(_02088_));
 OA222x2_ASAP7_75t_R _17952_ (.A1(_05723_),
    .A2(_02740_),
    .B1(_02741_),
    .B2(_02488_),
    .C1(_02743_),
    .C2(_02415_),
    .Y(_02089_));
 OA222x2_ASAP7_75t_R _17953_ (.A1(_05643_),
    .A2(_02740_),
    .B1(_02741_),
    .B2(_02490_),
    .C1(_02743_),
    .C2(_02416_),
    .Y(_02090_));
 AOI22x1_ASAP7_75t_R _17954_ (.A1(_00605_),
    .A2(_02748_),
    .B1(_02750_),
    .B2(_02417_),
    .Y(_02753_));
 OA21x2_ASAP7_75t_R _17955_ (.A1(_02491_),
    .A2(_02742_),
    .B(_02753_),
    .Y(_02091_));
 AOI22x1_ASAP7_75t_R _17956_ (.A1(_00571_),
    .A2(_02748_),
    .B1(_02750_),
    .B2(_02419_),
    .Y(_02754_));
 OA21x2_ASAP7_75t_R _17957_ (.A1(_02493_),
    .A2(_02742_),
    .B(_02754_),
    .Y(_02092_));
 AOI22x1_ASAP7_75t_R _17958_ (.A1(_00538_),
    .A2(_02748_),
    .B1(_02750_),
    .B2(_02421_),
    .Y(_02755_));
 OA21x2_ASAP7_75t_R _17959_ (.A1(_02495_),
    .A2(_02742_),
    .B(_02755_),
    .Y(_02093_));
 BUFx12f_ASAP7_75t_R _17960_ (.A(_02744_),
    .Y(_02756_));
 AOI22x1_ASAP7_75t_R _17961_ (.A1(_00505_),
    .A2(_02756_),
    .B1(_02750_),
    .B2(_02424_),
    .Y(_02757_));
 OA21x2_ASAP7_75t_R _17962_ (.A1(_02497_),
    .A2(_02742_),
    .B(_02757_),
    .Y(_02094_));
 AOI22x1_ASAP7_75t_R _17963_ (.A1(_00472_),
    .A2(_02756_),
    .B1(_02750_),
    .B2(_02426_),
    .Y(_02758_));
 OA21x2_ASAP7_75t_R _17964_ (.A1(_02500_),
    .A2(_02742_),
    .B(_02758_),
    .Y(_02095_));
 AOI22x1_ASAP7_75t_R _17965_ (.A1(_00439_),
    .A2(_02756_),
    .B1(_02750_),
    .B2(_02428_),
    .Y(_02759_));
 OA21x2_ASAP7_75t_R _17966_ (.A1(_02502_),
    .A2(_02742_),
    .B(_02759_),
    .Y(_02096_));
 NAND2x1_ASAP7_75t_R _17967_ (.A(_01037_),
    .B(_02748_),
    .Y(_02760_));
 OA21x2_ASAP7_75t_R _17968_ (.A1(_02504_),
    .A2(_02748_),
    .B(_02760_),
    .Y(_02097_));
 AOI22x1_ASAP7_75t_R _17969_ (.A1(_00406_),
    .A2(_02756_),
    .B1(_02750_),
    .B2(_02431_),
    .Y(_02761_));
 OA21x2_ASAP7_75t_R _17970_ (.A1(_02506_),
    .A2(_02742_),
    .B(_02761_),
    .Y(_02098_));
 AO21x1_ASAP7_75t_R _17971_ (.A1(_09051_),
    .A2(_02700_),
    .B(_04780_),
    .Y(_02762_));
 OA221x2_ASAP7_75t_R _17972_ (.A1(_02433_),
    .A2(_02748_),
    .B1(_02741_),
    .B2(_02508_),
    .C(_02762_),
    .Y(_02099_));
 BUFx4f_ASAP7_75t_R _17973_ (.A(_02741_),
    .Y(_02763_));
 BUFx6f_ASAP7_75t_R _17974_ (.A(_02749_),
    .Y(_02764_));
 AOI22x1_ASAP7_75t_R _17975_ (.A1(_00340_),
    .A2(_02756_),
    .B1(_02764_),
    .B2(_02438_),
    .Y(_02765_));
 OA21x2_ASAP7_75t_R _17976_ (.A1(_02511_),
    .A2(_02763_),
    .B(_02765_),
    .Y(_02100_));
 AOI22x1_ASAP7_75t_R _17977_ (.A1(_00306_),
    .A2(_02756_),
    .B1(_02764_),
    .B2(_02440_),
    .Y(_02766_));
 OA21x2_ASAP7_75t_R _17978_ (.A1(_02515_),
    .A2(_02763_),
    .B(_02766_),
    .Y(_02101_));
 AOI22x1_ASAP7_75t_R _17979_ (.A1(_00273_),
    .A2(_02756_),
    .B1(_02764_),
    .B2(_02442_),
    .Y(_02767_));
 OA21x2_ASAP7_75t_R _17980_ (.A1(_02517_),
    .A2(_02763_),
    .B(_02767_),
    .Y(_02102_));
 AOI22x1_ASAP7_75t_R _17981_ (.A1(_00240_),
    .A2(_02756_),
    .B1(_02764_),
    .B2(_02444_),
    .Y(_02768_));
 OA21x2_ASAP7_75t_R _17982_ (.A1(_02519_),
    .A2(_02763_),
    .B(_02768_),
    .Y(_02103_));
 AOI22x1_ASAP7_75t_R _17983_ (.A1(_00206_),
    .A2(_02756_),
    .B1(_02764_),
    .B2(_02446_),
    .Y(_02769_));
 OA21x2_ASAP7_75t_R _17984_ (.A1(_02521_),
    .A2(_02763_),
    .B(_02769_),
    .Y(_02104_));
 AOI22x1_ASAP7_75t_R _17985_ (.A1(_00173_),
    .A2(_02756_),
    .B1(_02764_),
    .B2(_02448_),
    .Y(_02770_));
 OA21x2_ASAP7_75t_R _17986_ (.A1(_02523_),
    .A2(_02763_),
    .B(_02770_),
    .Y(_02105_));
 OA222x2_ASAP7_75t_R _17987_ (.A1(_04010_),
    .A2(_02740_),
    .B1(_02741_),
    .B2(_02525_),
    .C1(_02743_),
    .C2(_02450_),
    .Y(_02106_));
 AOI22x1_ASAP7_75t_R _17988_ (.A1(_00106_),
    .A2(_02745_),
    .B1(_02764_),
    .B2(_02451_),
    .Y(_02771_));
 OA21x2_ASAP7_75t_R _17989_ (.A1(_02526_),
    .A2(_02763_),
    .B(_02771_),
    .Y(_02107_));
 NOR2x1_ASAP7_75t_R _17990_ (.A(_01004_),
    .B(_02740_),
    .Y(_02772_));
 AO21x1_ASAP7_75t_R _17991_ (.A1(_02528_),
    .A2(_02740_),
    .B(_02772_),
    .Y(_02108_));
 AND3x1_ASAP7_75t_R _17992_ (.A(_09503_),
    .B(_08873_),
    .C(_02700_),
    .Y(_02773_));
 NOR2x1_ASAP7_75t_R _17993_ (.A(_00072_),
    .B(_02740_),
    .Y(_02774_));
 AO221x1_ASAP7_75t_R _17994_ (.A1(_02454_),
    .A2(_02740_),
    .B1(_02773_),
    .B2(_02531_),
    .C(_02774_),
    .Y(_02109_));
 AND2x2_ASAP7_75t_R _17995_ (.A(_00040_),
    .B(_02745_),
    .Y(_02775_));
 AOI221x1_ASAP7_75t_R _17996_ (.A1(_02457_),
    .A2(_02773_),
    .B1(_02750_),
    .B2(_02533_),
    .C(_02775_),
    .Y(_02110_));
 AOI22x1_ASAP7_75t_R _17997_ (.A1(_00971_),
    .A2(_02745_),
    .B1(_02764_),
    .B2(_02459_),
    .Y(_02776_));
 OA21x2_ASAP7_75t_R _17998_ (.A1(_02535_),
    .A2(_02763_),
    .B(_02776_),
    .Y(_02111_));
 NAND2x1_ASAP7_75t_R _17999_ (.A(_00938_),
    .B(_02745_),
    .Y(_02777_));
 OA221x2_ASAP7_75t_R _18000_ (.A1(_02537_),
    .A2(_02748_),
    .B1(_02741_),
    .B2(_02461_),
    .C(_02777_),
    .Y(_02112_));
 NAND2x1_ASAP7_75t_R _18001_ (.A(_00904_),
    .B(_02745_),
    .Y(_02778_));
 OA221x2_ASAP7_75t_R _18002_ (.A1(_02463_),
    .A2(_02748_),
    .B1(_02741_),
    .B2(_02539_),
    .C(_02778_),
    .Y(_02113_));
 AOI22x1_ASAP7_75t_R _18003_ (.A1(_00871_),
    .A2(_02745_),
    .B1(_02764_),
    .B2(_02465_),
    .Y(_02779_));
 OA21x2_ASAP7_75t_R _18004_ (.A1(_02541_),
    .A2(_02763_),
    .B(_02779_),
    .Y(_02114_));
 NAND2x1_ASAP7_75t_R _18005_ (.A(_00837_),
    .B(_02744_),
    .Y(_02780_));
 OA21x2_ASAP7_75t_R _18006_ (.A1(_02544_),
    .A2(_02745_),
    .B(_02780_),
    .Y(_02781_));
 OA21x2_ASAP7_75t_R _18007_ (.A1(_02543_),
    .A2(_02763_),
    .B(_02781_),
    .Y(_02115_));
 AOI22x1_ASAP7_75t_R _18008_ (.A1(_00804_),
    .A2(_02745_),
    .B1(_02764_),
    .B2(_02469_),
    .Y(_02782_));
 OA21x2_ASAP7_75t_R _18009_ (.A1(_02547_),
    .A2(_02741_),
    .B(_02782_),
    .Y(_02116_));
 NAND2x1_ASAP7_75t_R _18010_ (.A(_00770_),
    .B(_02744_),
    .Y(_02783_));
 OA21x2_ASAP7_75t_R _18011_ (.A1(_02550_),
    .A2(_02745_),
    .B(_02783_),
    .Y(_02784_));
 OA21x2_ASAP7_75t_R _18012_ (.A1(_02549_),
    .A2(_02741_),
    .B(_02784_),
    .Y(_02117_));
 AND2x6_ASAP7_75t_R _18013_ (.A(_08097_),
    .B(_02693_),
    .Y(_02785_));
 NAND2x2_ASAP7_75t_R _18014_ (.A(_08606_),
    .B(_02785_),
    .Y(_02786_));
 BUFx10_ASAP7_75t_R _18015_ (.A(_02786_),
    .Y(_02787_));
 NAND2x2_ASAP7_75t_R _18016_ (.A(_08937_),
    .B(_02785_),
    .Y(_02788_));
 NAND2x2_ASAP7_75t_R _18017_ (.A(_08098_),
    .B(_02693_),
    .Y(_02789_));
 NAND2x1_ASAP7_75t_R _18018_ (.A(_00006_),
    .B(_02789_),
    .Y(_02790_));
 OA21x2_ASAP7_75t_R _18019_ (.A1(_08793_),
    .A2(_02788_),
    .B(_02790_),
    .Y(_02791_));
 OA21x2_ASAP7_75t_R _18020_ (.A1(_02400_),
    .A2(_02787_),
    .B(_02791_),
    .Y(_02118_));
 BUFx12f_ASAP7_75t_R _18021_ (.A(_02789_),
    .Y(_02792_));
 AND3x2_ASAP7_75t_R _18022_ (.A(_08117_),
    .B(_08701_),
    .C(_02700_),
    .Y(_02793_));
 BUFx12f_ASAP7_75t_R _18023_ (.A(_02793_),
    .Y(_02794_));
 AOI22x1_ASAP7_75t_R _18024_ (.A1(_00738_),
    .A2(_02792_),
    .B1(_02794_),
    .B2(_02411_),
    .Y(_02795_));
 OA21x2_ASAP7_75t_R _18025_ (.A1(_02480_),
    .A2(_02787_),
    .B(_02795_),
    .Y(_02119_));
 AOI22x1_ASAP7_75t_R _18026_ (.A1(_00705_),
    .A2(_02792_),
    .B1(_02794_),
    .B2(_02413_),
    .Y(_02796_));
 OA21x2_ASAP7_75t_R _18027_ (.A1(_02485_),
    .A2(_02787_),
    .B(_02796_),
    .Y(_02120_));
 INVx1_ASAP7_75t_R _18028_ (.A(_00672_),
    .Y(_02797_));
 OA222x2_ASAP7_75t_R _18029_ (.A1(_02797_),
    .A2(_02785_),
    .B1(_02786_),
    .B2(_02488_),
    .C1(_02788_),
    .C2(_02415_),
    .Y(_02121_));
 INVx1_ASAP7_75t_R _18030_ (.A(_00639_),
    .Y(_02798_));
 OA222x2_ASAP7_75t_R _18031_ (.A1(_02798_),
    .A2(_02785_),
    .B1(_02786_),
    .B2(_02490_),
    .C1(_02788_),
    .C2(_02416_),
    .Y(_02122_));
 AOI22x1_ASAP7_75t_R _18032_ (.A1(_00606_),
    .A2(_02792_),
    .B1(_02794_),
    .B2(_02417_),
    .Y(_02799_));
 OA21x2_ASAP7_75t_R _18033_ (.A1(_02491_),
    .A2(_02787_),
    .B(_02799_),
    .Y(_02123_));
 AOI22x1_ASAP7_75t_R _18034_ (.A1(_00572_),
    .A2(_02792_),
    .B1(_02794_),
    .B2(_02419_),
    .Y(_02800_));
 OA21x2_ASAP7_75t_R _18035_ (.A1(_02493_),
    .A2(_02787_),
    .B(_02800_),
    .Y(_02124_));
 AOI22x1_ASAP7_75t_R _18036_ (.A1(_00539_),
    .A2(_02792_),
    .B1(_02794_),
    .B2(_02421_),
    .Y(_02801_));
 OA21x2_ASAP7_75t_R _18037_ (.A1(_02495_),
    .A2(_02787_),
    .B(_02801_),
    .Y(_02125_));
 BUFx16f_ASAP7_75t_R _18038_ (.A(_02789_),
    .Y(_02802_));
 AOI22x1_ASAP7_75t_R _18039_ (.A1(_00506_),
    .A2(_02802_),
    .B1(_02794_),
    .B2(_02424_),
    .Y(_02803_));
 OA21x2_ASAP7_75t_R _18040_ (.A1(_02497_),
    .A2(_02787_),
    .B(_02803_),
    .Y(_02126_));
 AOI22x1_ASAP7_75t_R _18041_ (.A1(_00473_),
    .A2(_02802_),
    .B1(_02794_),
    .B2(_02426_),
    .Y(_02804_));
 OA21x2_ASAP7_75t_R _18042_ (.A1(_02500_),
    .A2(_02787_),
    .B(_02804_),
    .Y(_02127_));
 AOI22x1_ASAP7_75t_R _18043_ (.A1(_00440_),
    .A2(_02802_),
    .B1(_02794_),
    .B2(_02428_),
    .Y(_02805_));
 OA21x2_ASAP7_75t_R _18044_ (.A1(_02502_),
    .A2(_02787_),
    .B(_02805_),
    .Y(_02128_));
 NAND2x1_ASAP7_75t_R _18045_ (.A(_01038_),
    .B(_02792_),
    .Y(_02806_));
 OA21x2_ASAP7_75t_R _18046_ (.A1(_02504_),
    .A2(_02792_),
    .B(_02806_),
    .Y(_02129_));
 AOI22x1_ASAP7_75t_R _18047_ (.A1(_00407_),
    .A2(_02802_),
    .B1(_02794_),
    .B2(_02431_),
    .Y(_02807_));
 OA21x2_ASAP7_75t_R _18048_ (.A1(_02506_),
    .A2(_02787_),
    .B(_02807_),
    .Y(_02130_));
 BUFx6f_ASAP7_75t_R _18049_ (.A(_02789_),
    .Y(_02808_));
 NAND2x1_ASAP7_75t_R _18050_ (.A(_00374_),
    .B(_02808_),
    .Y(_02809_));
 OA221x2_ASAP7_75t_R _18051_ (.A1(_02433_),
    .A2(_02792_),
    .B1(_02786_),
    .B2(_02508_),
    .C(_02809_),
    .Y(_02131_));
 BUFx4f_ASAP7_75t_R _18052_ (.A(_02786_),
    .Y(_02810_));
 BUFx6f_ASAP7_75t_R _18053_ (.A(_02793_),
    .Y(_02811_));
 AOI22x1_ASAP7_75t_R _18054_ (.A1(_00341_),
    .A2(_02802_),
    .B1(_02811_),
    .B2(_02438_),
    .Y(_02812_));
 OA21x2_ASAP7_75t_R _18055_ (.A1(_02511_),
    .A2(_02810_),
    .B(_02812_),
    .Y(_02132_));
 AOI22x1_ASAP7_75t_R _18056_ (.A1(_00307_),
    .A2(_02802_),
    .B1(_02811_),
    .B2(_02440_),
    .Y(_02813_));
 OA21x2_ASAP7_75t_R _18057_ (.A1(_02515_),
    .A2(_02810_),
    .B(_02813_),
    .Y(_02133_));
 AOI22x1_ASAP7_75t_R _18058_ (.A1(_00274_),
    .A2(_02802_),
    .B1(_02811_),
    .B2(_02442_),
    .Y(_02814_));
 OA21x2_ASAP7_75t_R _18059_ (.A1(_02517_),
    .A2(_02810_),
    .B(_02814_),
    .Y(_02134_));
 AOI22x1_ASAP7_75t_R _18060_ (.A1(_00241_),
    .A2(_02802_),
    .B1(_02811_),
    .B2(_02444_),
    .Y(_02815_));
 OA21x2_ASAP7_75t_R _18061_ (.A1(_02519_),
    .A2(_02810_),
    .B(_02815_),
    .Y(_02135_));
 AOI22x1_ASAP7_75t_R _18062_ (.A1(_00207_),
    .A2(_02802_),
    .B1(_02811_),
    .B2(_02446_),
    .Y(_02816_));
 OA21x2_ASAP7_75t_R _18063_ (.A1(_02521_),
    .A2(_02810_),
    .B(_02816_),
    .Y(_02136_));
 AOI22x1_ASAP7_75t_R _18064_ (.A1(_00174_),
    .A2(_02802_),
    .B1(_02811_),
    .B2(_02448_),
    .Y(_02817_));
 OA21x2_ASAP7_75t_R _18065_ (.A1(_02523_),
    .A2(_02810_),
    .B(_02817_),
    .Y(_02137_));
 INVx1_ASAP7_75t_R _18066_ (.A(_00140_),
    .Y(_02818_));
 OA222x2_ASAP7_75t_R _18067_ (.A1(_02818_),
    .A2(_02785_),
    .B1(_02786_),
    .B2(_02525_),
    .C1(_02788_),
    .C2(_02450_),
    .Y(_02138_));
 AOI22x1_ASAP7_75t_R _18068_ (.A1(_00107_),
    .A2(_02808_),
    .B1(_02811_),
    .B2(_02451_),
    .Y(_02819_));
 OA21x2_ASAP7_75t_R _18069_ (.A1(_02526_),
    .A2(_02810_),
    .B(_02819_),
    .Y(_02139_));
 NOR2x1_ASAP7_75t_R _18070_ (.A(_01005_),
    .B(_02785_),
    .Y(_02820_));
 AO21x1_ASAP7_75t_R _18071_ (.A1(_02528_),
    .A2(_02785_),
    .B(_02820_),
    .Y(_02140_));
 AND3x1_ASAP7_75t_R _18072_ (.A(_08145_),
    .B(_08577_),
    .C(_02700_),
    .Y(_02821_));
 NOR2x1_ASAP7_75t_R _18073_ (.A(_00073_),
    .B(_02785_),
    .Y(_02822_));
 AO221x1_ASAP7_75t_R _18074_ (.A1(_02454_),
    .A2(_02785_),
    .B1(_02821_),
    .B2(_02531_),
    .C(_02822_),
    .Y(_02141_));
 AND2x2_ASAP7_75t_R _18075_ (.A(_00041_),
    .B(_02808_),
    .Y(_02823_));
 AOI221x1_ASAP7_75t_R _18076_ (.A1(_02457_),
    .A2(_02821_),
    .B1(_02794_),
    .B2(_02533_),
    .C(_02823_),
    .Y(_02142_));
 AOI22x1_ASAP7_75t_R _18077_ (.A1(_00972_),
    .A2(_02808_),
    .B1(_02811_),
    .B2(_02459_),
    .Y(_02824_));
 OA21x2_ASAP7_75t_R _18078_ (.A1(_02535_),
    .A2(_02810_),
    .B(_02824_),
    .Y(_02143_));
 NAND2x1_ASAP7_75t_R _18079_ (.A(_00939_),
    .B(_02808_),
    .Y(_02825_));
 OA221x2_ASAP7_75t_R _18080_ (.A1(_02537_),
    .A2(_02792_),
    .B1(_02786_),
    .B2(_02461_),
    .C(_02825_),
    .Y(_02144_));
 NAND2x1_ASAP7_75t_R _18081_ (.A(_00905_),
    .B(_02808_),
    .Y(_02826_));
 OA221x2_ASAP7_75t_R _18082_ (.A1(_02463_),
    .A2(_02792_),
    .B1(_02786_),
    .B2(_02539_),
    .C(_02826_),
    .Y(_02145_));
 AOI22x1_ASAP7_75t_R _18083_ (.A1(_00872_),
    .A2(_02808_),
    .B1(_02811_),
    .B2(_02465_),
    .Y(_02827_));
 OA21x2_ASAP7_75t_R _18084_ (.A1(_02541_),
    .A2(_02810_),
    .B(_02827_),
    .Y(_02146_));
 NAND2x1_ASAP7_75t_R _18085_ (.A(_00838_),
    .B(_02789_),
    .Y(_02828_));
 OA21x2_ASAP7_75t_R _18086_ (.A1(_02544_),
    .A2(_02808_),
    .B(_02828_),
    .Y(_02829_));
 OA21x2_ASAP7_75t_R _18087_ (.A1(_02543_),
    .A2(_02810_),
    .B(_02829_),
    .Y(_02147_));
 AOI22x1_ASAP7_75t_R _18088_ (.A1(_00805_),
    .A2(_02808_),
    .B1(_02811_),
    .B2(_02469_),
    .Y(_02830_));
 OA21x2_ASAP7_75t_R _18089_ (.A1(_02547_),
    .A2(_02786_),
    .B(_02830_),
    .Y(_02148_));
 NAND2x1_ASAP7_75t_R _18090_ (.A(_00771_),
    .B(_02789_),
    .Y(_02831_));
 OA21x2_ASAP7_75t_R _18091_ (.A1(_02550_),
    .A2(_02808_),
    .B(_02831_),
    .Y(_02832_));
 OA21x2_ASAP7_75t_R _18092_ (.A1(_02549_),
    .A2(_02786_),
    .B(_02832_),
    .Y(_02149_));
 AND2x6_ASAP7_75t_R _18093_ (.A(_08689_),
    .B(_02693_),
    .Y(_02833_));
 NAND2x2_ASAP7_75t_R _18094_ (.A(_08606_),
    .B(_02833_),
    .Y(_02834_));
 BUFx10_ASAP7_75t_R _18095_ (.A(_02834_),
    .Y(_02835_));
 NAND2x2_ASAP7_75t_R _18096_ (.A(_08114_),
    .B(_02833_),
    .Y(_02836_));
 OA22x2_ASAP7_75t_R _18097_ (.A1(_03035_),
    .A2(_02833_),
    .B1(_02836_),
    .B2(_09330_),
    .Y(_02837_));
 OA21x2_ASAP7_75t_R _18098_ (.A1(_02400_),
    .A2(_02835_),
    .B(_02837_),
    .Y(_02150_));
 NAND2x2_ASAP7_75t_R _18099_ (.A(_08694_),
    .B(_02693_),
    .Y(_02838_));
 BUFx12f_ASAP7_75t_R _18100_ (.A(_02838_),
    .Y(_02839_));
 AND3x2_ASAP7_75t_R _18101_ (.A(_08701_),
    .B(_08694_),
    .C(_02700_),
    .Y(_02840_));
 BUFx12f_ASAP7_75t_R _18102_ (.A(_02840_),
    .Y(_02841_));
 AOI22x1_ASAP7_75t_R _18103_ (.A1(_00739_),
    .A2(_02839_),
    .B1(_02841_),
    .B2(_02411_),
    .Y(_02842_));
 OA21x2_ASAP7_75t_R _18104_ (.A1(_02480_),
    .A2(_02835_),
    .B(_02842_),
    .Y(_02151_));
 AOI22x1_ASAP7_75t_R _18105_ (.A1(_00706_),
    .A2(_02839_),
    .B1(_02841_),
    .B2(_02413_),
    .Y(_02843_));
 OA21x2_ASAP7_75t_R _18106_ (.A1(_02485_),
    .A2(_02835_),
    .B(_02843_),
    .Y(_02152_));
 INVx1_ASAP7_75t_R _18107_ (.A(_00673_),
    .Y(_02844_));
 OA222x2_ASAP7_75t_R _18108_ (.A1(_02844_),
    .A2(_02833_),
    .B1(_02834_),
    .B2(_02488_),
    .C1(_02836_),
    .C2(_02415_),
    .Y(_02153_));
 INVx1_ASAP7_75t_R _18109_ (.A(_00640_),
    .Y(_02845_));
 OA222x2_ASAP7_75t_R _18110_ (.A1(_02845_),
    .A2(_02833_),
    .B1(_02834_),
    .B2(_02490_),
    .C1(_02836_),
    .C2(_02416_),
    .Y(_02154_));
 AOI22x1_ASAP7_75t_R _18111_ (.A1(_00607_),
    .A2(_02839_),
    .B1(_02841_),
    .B2(_02417_),
    .Y(_02846_));
 OA21x2_ASAP7_75t_R _18112_ (.A1(_02491_),
    .A2(_02835_),
    .B(_02846_),
    .Y(_02155_));
 AOI22x1_ASAP7_75t_R _18113_ (.A1(_00573_),
    .A2(_02839_),
    .B1(_02841_),
    .B2(_02419_),
    .Y(_02847_));
 OA21x2_ASAP7_75t_R _18114_ (.A1(_02493_),
    .A2(_02835_),
    .B(_02847_),
    .Y(_02156_));
 AOI22x1_ASAP7_75t_R _18115_ (.A1(_00540_),
    .A2(_02839_),
    .B1(_02841_),
    .B2(_02421_),
    .Y(_02848_));
 OA21x2_ASAP7_75t_R _18116_ (.A1(_02495_),
    .A2(_02835_),
    .B(_02848_),
    .Y(_02157_));
 BUFx16f_ASAP7_75t_R _18117_ (.A(_02838_),
    .Y(_02849_));
 AOI22x1_ASAP7_75t_R _18118_ (.A1(_00507_),
    .A2(_02849_),
    .B1(_02841_),
    .B2(_02424_),
    .Y(_02850_));
 OA21x2_ASAP7_75t_R _18119_ (.A1(_02497_),
    .A2(_02835_),
    .B(_02850_),
    .Y(_02158_));
 AOI22x1_ASAP7_75t_R _18120_ (.A1(_00474_),
    .A2(_02849_),
    .B1(_02841_),
    .B2(_02426_),
    .Y(_02851_));
 OA21x2_ASAP7_75t_R _18121_ (.A1(_02500_),
    .A2(_02835_),
    .B(_02851_),
    .Y(_02159_));
 AOI22x1_ASAP7_75t_R _18122_ (.A1(_00441_),
    .A2(_02849_),
    .B1(_02841_),
    .B2(_02428_),
    .Y(_02852_));
 OA21x2_ASAP7_75t_R _18123_ (.A1(_02502_),
    .A2(_02835_),
    .B(_02852_),
    .Y(_02160_));
 NAND2x1_ASAP7_75t_R _18124_ (.A(_01039_),
    .B(_02839_),
    .Y(_02853_));
 OA21x2_ASAP7_75t_R _18125_ (.A1(_02504_),
    .A2(_02839_),
    .B(_02853_),
    .Y(_02161_));
 AOI22x1_ASAP7_75t_R _18126_ (.A1(_00408_),
    .A2(_02849_),
    .B1(_02841_),
    .B2(_02431_),
    .Y(_02854_));
 OA21x2_ASAP7_75t_R _18127_ (.A1(_02506_),
    .A2(_02835_),
    .B(_02854_),
    .Y(_02162_));
 BUFx6f_ASAP7_75t_R _18128_ (.A(_02838_),
    .Y(_02855_));
 NAND2x1_ASAP7_75t_R _18129_ (.A(_00375_),
    .B(_02855_),
    .Y(_02856_));
 OA221x2_ASAP7_75t_R _18130_ (.A1(_02433_),
    .A2(_02839_),
    .B1(_02834_),
    .B2(_02508_),
    .C(_02856_),
    .Y(_02163_));
 BUFx4f_ASAP7_75t_R _18131_ (.A(_02834_),
    .Y(_02857_));
 BUFx6f_ASAP7_75t_R _18132_ (.A(_02840_),
    .Y(_02858_));
 AOI22x1_ASAP7_75t_R _18133_ (.A1(_00342_),
    .A2(_02849_),
    .B1(_02858_),
    .B2(_02438_),
    .Y(_02859_));
 OA21x2_ASAP7_75t_R _18134_ (.A1(_02511_),
    .A2(_02857_),
    .B(_02859_),
    .Y(_02164_));
 AOI22x1_ASAP7_75t_R _18135_ (.A1(_00308_),
    .A2(_02849_),
    .B1(_02858_),
    .B2(_02440_),
    .Y(_02860_));
 OA21x2_ASAP7_75t_R _18136_ (.A1(_02515_),
    .A2(_02857_),
    .B(_02860_),
    .Y(_02165_));
 AOI22x1_ASAP7_75t_R _18137_ (.A1(_00275_),
    .A2(_02849_),
    .B1(_02858_),
    .B2(_02442_),
    .Y(_02861_));
 OA21x2_ASAP7_75t_R _18138_ (.A1(_02517_),
    .A2(_02857_),
    .B(_02861_),
    .Y(_02166_));
 AOI22x1_ASAP7_75t_R _18139_ (.A1(_00242_),
    .A2(_02849_),
    .B1(_02858_),
    .B2(_02444_),
    .Y(_02862_));
 OA21x2_ASAP7_75t_R _18140_ (.A1(_02519_),
    .A2(_02857_),
    .B(_02862_),
    .Y(_02167_));
 AOI22x1_ASAP7_75t_R _18141_ (.A1(_00208_),
    .A2(_02849_),
    .B1(_02858_),
    .B2(_02446_),
    .Y(_02863_));
 OA21x2_ASAP7_75t_R _18142_ (.A1(_02521_),
    .A2(_02857_),
    .B(_02863_),
    .Y(_02168_));
 AOI22x1_ASAP7_75t_R _18143_ (.A1(_00175_),
    .A2(_02849_),
    .B1(_02858_),
    .B2(_02448_),
    .Y(_02864_));
 OA21x2_ASAP7_75t_R _18144_ (.A1(_02523_),
    .A2(_02857_),
    .B(_02864_),
    .Y(_02169_));
 INVx1_ASAP7_75t_R _18145_ (.A(_00141_),
    .Y(_02865_));
 OA222x2_ASAP7_75t_R _18146_ (.A1(_02865_),
    .A2(_02833_),
    .B1(_02834_),
    .B2(_02525_),
    .C1(_02836_),
    .C2(_02450_),
    .Y(_02170_));
 AOI22x1_ASAP7_75t_R _18147_ (.A1(_00108_),
    .A2(_02855_),
    .B1(_02858_),
    .B2(_02451_),
    .Y(_02866_));
 OA21x2_ASAP7_75t_R _18148_ (.A1(_02526_),
    .A2(_02857_),
    .B(_02866_),
    .Y(_02171_));
 NOR2x1_ASAP7_75t_R _18149_ (.A(_01006_),
    .B(_02833_),
    .Y(_02867_));
 AO21x1_ASAP7_75t_R _18150_ (.A1(_02528_),
    .A2(_02833_),
    .B(_02867_),
    .Y(_02172_));
 AND3x1_ASAP7_75t_R _18151_ (.A(_09503_),
    .B(_08750_),
    .C(_02700_),
    .Y(_02868_));
 NOR2x1_ASAP7_75t_R _18152_ (.A(_00074_),
    .B(_02833_),
    .Y(_02869_));
 AO221x1_ASAP7_75t_R _18153_ (.A1(_02454_),
    .A2(_02833_),
    .B1(_02868_),
    .B2(_02531_),
    .C(_02869_),
    .Y(_02173_));
 AND2x2_ASAP7_75t_R _18154_ (.A(_00042_),
    .B(_02855_),
    .Y(_02870_));
 AOI221x1_ASAP7_75t_R _18155_ (.A1(_02457_),
    .A2(_02868_),
    .B1(_02841_),
    .B2(_02533_),
    .C(_02870_),
    .Y(_02174_));
 AOI22x1_ASAP7_75t_R _18156_ (.A1(_00973_),
    .A2(_02855_),
    .B1(_02858_),
    .B2(_02459_),
    .Y(_02871_));
 OA21x2_ASAP7_75t_R _18157_ (.A1(_02535_),
    .A2(_02857_),
    .B(_02871_),
    .Y(_02175_));
 NAND2x1_ASAP7_75t_R _18158_ (.A(_00940_),
    .B(_02855_),
    .Y(_02872_));
 OA221x2_ASAP7_75t_R _18159_ (.A1(_02537_),
    .A2(_02839_),
    .B1(_02834_),
    .B2(_02461_),
    .C(_02872_),
    .Y(_02176_));
 NAND2x1_ASAP7_75t_R _18160_ (.A(_00906_),
    .B(_02855_),
    .Y(_02873_));
 OA221x2_ASAP7_75t_R _18161_ (.A1(_02463_),
    .A2(_02839_),
    .B1(_02834_),
    .B2(_02539_),
    .C(_02873_),
    .Y(_02177_));
 AOI22x1_ASAP7_75t_R _18162_ (.A1(_00873_),
    .A2(_02855_),
    .B1(_02858_),
    .B2(_02465_),
    .Y(_02874_));
 OA21x2_ASAP7_75t_R _18163_ (.A1(_02541_),
    .A2(_02857_),
    .B(_02874_),
    .Y(_02178_));
 NAND2x1_ASAP7_75t_R _18164_ (.A(_00839_),
    .B(_02838_),
    .Y(_02875_));
 OA21x2_ASAP7_75t_R _18165_ (.A1(_02544_),
    .A2(_02855_),
    .B(_02875_),
    .Y(_02876_));
 OA21x2_ASAP7_75t_R _18166_ (.A1(_02543_),
    .A2(_02857_),
    .B(_02876_),
    .Y(_02179_));
 AOI22x1_ASAP7_75t_R _18167_ (.A1(_00806_),
    .A2(_02855_),
    .B1(_02858_),
    .B2(_02469_),
    .Y(_02877_));
 OA21x2_ASAP7_75t_R _18168_ (.A1(_02547_),
    .A2(_02834_),
    .B(_02877_),
    .Y(_02180_));
 NAND2x1_ASAP7_75t_R _18169_ (.A(_00772_),
    .B(_02838_),
    .Y(_02878_));
 OA21x2_ASAP7_75t_R _18170_ (.A1(_02550_),
    .A2(_02855_),
    .B(_02878_),
    .Y(_02879_));
 OA21x2_ASAP7_75t_R _18171_ (.A1(_02549_),
    .A2(_02834_),
    .B(_02879_),
    .Y(_02181_));
 AND2x6_ASAP7_75t_R _18172_ (.A(_08102_),
    .B(_08787_),
    .Y(_02880_));
 NAND2x2_ASAP7_75t_R _18173_ (.A(_08606_),
    .B(_02880_),
    .Y(_02881_));
 BUFx10_ASAP7_75t_R _18174_ (.A(_02881_),
    .Y(_02882_));
 NAND2x2_ASAP7_75t_R _18175_ (.A(_08114_),
    .B(_02880_),
    .Y(_02883_));
 OA22x2_ASAP7_75t_R _18176_ (.A1(_03129_),
    .A2(_02880_),
    .B1(_02883_),
    .B2(_08110_),
    .Y(_02884_));
 OA21x2_ASAP7_75t_R _18177_ (.A1(_02400_),
    .A2(_02882_),
    .B(_02884_),
    .Y(_02182_));
 NAND2x2_ASAP7_75t_R _18178_ (.A(_08102_),
    .B(_08795_),
    .Y(_02885_));
 BUFx12f_ASAP7_75t_R _18179_ (.A(_02885_),
    .Y(_02886_));
 AND3x2_ASAP7_75t_R _18180_ (.A(_08146_),
    .B(_08701_),
    .C(_08795_),
    .Y(_02887_));
 BUFx12f_ASAP7_75t_R _18181_ (.A(_02887_),
    .Y(_02888_));
 AOI22x1_ASAP7_75t_R _18182_ (.A1(_00740_),
    .A2(_02886_),
    .B1(_02888_),
    .B2(_02411_),
    .Y(_02889_));
 OA21x2_ASAP7_75t_R _18183_ (.A1(_02480_),
    .A2(_02882_),
    .B(_02889_),
    .Y(_02183_));
 AOI22x1_ASAP7_75t_R _18184_ (.A1(_00707_),
    .A2(_02886_),
    .B1(_02888_),
    .B2(_02413_),
    .Y(_02890_));
 OA21x2_ASAP7_75t_R _18185_ (.A1(_02485_),
    .A2(_02882_),
    .B(_02890_),
    .Y(_02184_));
 INVx1_ASAP7_75t_R _18186_ (.A(_00674_),
    .Y(_02891_));
 OA222x2_ASAP7_75t_R _18187_ (.A1(_02891_),
    .A2(_02880_),
    .B1(_02881_),
    .B2(_02488_),
    .C1(_02883_),
    .C2(_02415_),
    .Y(_02185_));
 INVx1_ASAP7_75t_R _18188_ (.A(_00641_),
    .Y(_02892_));
 OA222x2_ASAP7_75t_R _18189_ (.A1(_02892_),
    .A2(_02880_),
    .B1(_02881_),
    .B2(_02490_),
    .C1(_02883_),
    .C2(_02416_),
    .Y(_02186_));
 AOI22x1_ASAP7_75t_R _18190_ (.A1(_00608_),
    .A2(_02886_),
    .B1(_02888_),
    .B2(_02417_),
    .Y(_02893_));
 OA21x2_ASAP7_75t_R _18191_ (.A1(_02491_),
    .A2(_02882_),
    .B(_02893_),
    .Y(_02187_));
 AOI22x1_ASAP7_75t_R _18192_ (.A1(_00574_),
    .A2(_02886_),
    .B1(_02888_),
    .B2(_02419_),
    .Y(_02894_));
 OA21x2_ASAP7_75t_R _18193_ (.A1(_02493_),
    .A2(_02882_),
    .B(_02894_),
    .Y(_02188_));
 AOI22x1_ASAP7_75t_R _18194_ (.A1(_00541_),
    .A2(_02886_),
    .B1(_02888_),
    .B2(_02421_),
    .Y(_02895_));
 OA21x2_ASAP7_75t_R _18195_ (.A1(_02495_),
    .A2(_02882_),
    .B(_02895_),
    .Y(_02189_));
 BUFx16f_ASAP7_75t_R _18196_ (.A(_02885_),
    .Y(_02896_));
 AOI22x1_ASAP7_75t_R _18197_ (.A1(_00508_),
    .A2(_02896_),
    .B1(_02888_),
    .B2(_02424_),
    .Y(_02897_));
 OA21x2_ASAP7_75t_R _18198_ (.A1(_02497_),
    .A2(_02882_),
    .B(_02897_),
    .Y(_02190_));
 AOI22x1_ASAP7_75t_R _18199_ (.A1(_00475_),
    .A2(_02896_),
    .B1(_02888_),
    .B2(_02426_),
    .Y(_02898_));
 OA21x2_ASAP7_75t_R _18200_ (.A1(_02500_),
    .A2(_02882_),
    .B(_02898_),
    .Y(_02191_));
 AOI22x1_ASAP7_75t_R _18201_ (.A1(_00442_),
    .A2(_02896_),
    .B1(_02888_),
    .B2(_02428_),
    .Y(_02899_));
 OA21x2_ASAP7_75t_R _18202_ (.A1(_02502_),
    .A2(_02882_),
    .B(_02899_),
    .Y(_02192_));
 NAND2x1_ASAP7_75t_R _18203_ (.A(_01040_),
    .B(_02886_),
    .Y(_02900_));
 OA21x2_ASAP7_75t_R _18204_ (.A1(_02504_),
    .A2(_02886_),
    .B(_02900_),
    .Y(_02193_));
 AOI22x1_ASAP7_75t_R _18205_ (.A1(_00409_),
    .A2(_02896_),
    .B1(_02888_),
    .B2(_02431_),
    .Y(_02901_));
 OA21x2_ASAP7_75t_R _18206_ (.A1(_02506_),
    .A2(_02882_),
    .B(_02901_),
    .Y(_02194_));
 BUFx6f_ASAP7_75t_R _18207_ (.A(_02885_),
    .Y(_02902_));
 NAND2x1_ASAP7_75t_R _18208_ (.A(_00376_),
    .B(_02902_),
    .Y(_02903_));
 OA221x2_ASAP7_75t_R _18209_ (.A1(_02433_),
    .A2(_02886_),
    .B1(_02881_),
    .B2(_02508_),
    .C(_02903_),
    .Y(_02195_));
 BUFx4f_ASAP7_75t_R _18210_ (.A(_02881_),
    .Y(_02904_));
 BUFx6f_ASAP7_75t_R _18211_ (.A(_02887_),
    .Y(_02905_));
 AOI22x1_ASAP7_75t_R _18212_ (.A1(_00343_),
    .A2(_02896_),
    .B1(_02905_),
    .B2(_02438_),
    .Y(_02906_));
 OA21x2_ASAP7_75t_R _18213_ (.A1(_02511_),
    .A2(_02904_),
    .B(_02906_),
    .Y(_02196_));
 AOI22x1_ASAP7_75t_R _18214_ (.A1(_00309_),
    .A2(_02896_),
    .B1(_02905_),
    .B2(_02440_),
    .Y(_02907_));
 OA21x2_ASAP7_75t_R _18215_ (.A1(_02515_),
    .A2(_02904_),
    .B(_02907_),
    .Y(_02197_));
 AOI22x1_ASAP7_75t_R _18216_ (.A1(_00276_),
    .A2(_02896_),
    .B1(_02905_),
    .B2(_02442_),
    .Y(_02908_));
 OA21x2_ASAP7_75t_R _18217_ (.A1(_02517_),
    .A2(_02904_),
    .B(_02908_),
    .Y(_02198_));
 AOI22x1_ASAP7_75t_R _18218_ (.A1(_00243_),
    .A2(_02896_),
    .B1(_02905_),
    .B2(_02444_),
    .Y(_02909_));
 OA21x2_ASAP7_75t_R _18219_ (.A1(_02519_),
    .A2(_02904_),
    .B(_02909_),
    .Y(_02199_));
 AOI22x1_ASAP7_75t_R _18220_ (.A1(_00209_),
    .A2(_02896_),
    .B1(_02905_),
    .B2(_02446_),
    .Y(_02910_));
 OA21x2_ASAP7_75t_R _18221_ (.A1(_02521_),
    .A2(_02904_),
    .B(_02910_),
    .Y(_02200_));
 AOI22x1_ASAP7_75t_R _18222_ (.A1(_00176_),
    .A2(_02896_),
    .B1(_02905_),
    .B2(_02448_),
    .Y(_02911_));
 OA21x2_ASAP7_75t_R _18223_ (.A1(_02523_),
    .A2(_02904_),
    .B(_02911_),
    .Y(_02201_));
 INVx1_ASAP7_75t_R _18224_ (.A(_00142_),
    .Y(_02912_));
 OA222x2_ASAP7_75t_R _18225_ (.A1(_02912_),
    .A2(_02880_),
    .B1(_02881_),
    .B2(_02525_),
    .C1(_02883_),
    .C2(_02450_),
    .Y(_02202_));
 AOI22x1_ASAP7_75t_R _18226_ (.A1(_00109_),
    .A2(_02902_),
    .B1(_02905_),
    .B2(_02451_),
    .Y(_02913_));
 OA21x2_ASAP7_75t_R _18227_ (.A1(_02526_),
    .A2(_02904_),
    .B(_02913_),
    .Y(_02203_));
 NOR2x1_ASAP7_75t_R _18228_ (.A(_01007_),
    .B(_02880_),
    .Y(_02914_));
 AO21x1_ASAP7_75t_R _18229_ (.A1(_02528_),
    .A2(_02880_),
    .B(_02914_),
    .Y(_02204_));
 AND3x1_ASAP7_75t_R _18230_ (.A(_08146_),
    .B(_08577_),
    .C(_08788_),
    .Y(_02915_));
 NOR2x1_ASAP7_75t_R _18231_ (.A(_00075_),
    .B(_02880_),
    .Y(_02916_));
 AO221x1_ASAP7_75t_R _18232_ (.A1(_02454_),
    .A2(_02880_),
    .B1(_02915_),
    .B2(_02531_),
    .C(_02916_),
    .Y(_02205_));
 AND2x2_ASAP7_75t_R _18233_ (.A(_00043_),
    .B(_02902_),
    .Y(_02917_));
 AOI221x1_ASAP7_75t_R _18234_ (.A1(_02457_),
    .A2(_02915_),
    .B1(_02888_),
    .B2(_02533_),
    .C(_02917_),
    .Y(_02206_));
 AOI22x1_ASAP7_75t_R _18235_ (.A1(_00974_),
    .A2(_02902_),
    .B1(_02905_),
    .B2(_02459_),
    .Y(_02918_));
 OA21x2_ASAP7_75t_R _18236_ (.A1(_02535_),
    .A2(_02904_),
    .B(_02918_),
    .Y(_02207_));
 NAND2x1_ASAP7_75t_R _18237_ (.A(_00941_),
    .B(_02902_),
    .Y(_02919_));
 OA221x2_ASAP7_75t_R _18238_ (.A1(_02537_),
    .A2(_02886_),
    .B1(_02881_),
    .B2(_02461_),
    .C(_02919_),
    .Y(_02208_));
 NAND2x1_ASAP7_75t_R _18239_ (.A(_00907_),
    .B(_02902_),
    .Y(_02920_));
 OA221x2_ASAP7_75t_R _18240_ (.A1(_02463_),
    .A2(_02886_),
    .B1(_02881_),
    .B2(_02539_),
    .C(_02920_),
    .Y(_02209_));
 AOI22x1_ASAP7_75t_R _18241_ (.A1(_00874_),
    .A2(_02902_),
    .B1(_02905_),
    .B2(_02465_),
    .Y(_02921_));
 OA21x2_ASAP7_75t_R _18242_ (.A1(_02541_),
    .A2(_02904_),
    .B(_02921_),
    .Y(_02210_));
 NAND2x1_ASAP7_75t_R _18243_ (.A(_00840_),
    .B(_02885_),
    .Y(_02922_));
 OA21x2_ASAP7_75t_R _18244_ (.A1(_02544_),
    .A2(_02902_),
    .B(_02922_),
    .Y(_02923_));
 OA21x2_ASAP7_75t_R _18245_ (.A1(_02543_),
    .A2(_02904_),
    .B(_02923_),
    .Y(_02211_));
 AOI22x1_ASAP7_75t_R _18246_ (.A1(_00807_),
    .A2(_02902_),
    .B1(_02905_),
    .B2(_02469_),
    .Y(_02924_));
 OA21x2_ASAP7_75t_R _18247_ (.A1(_02547_),
    .A2(_02881_),
    .B(_02924_),
    .Y(_02212_));
 NAND2x1_ASAP7_75t_R _18248_ (.A(_00773_),
    .B(_02885_),
    .Y(_02925_));
 OA21x2_ASAP7_75t_R _18249_ (.A1(_02550_),
    .A2(_02902_),
    .B(_02925_),
    .Y(_02926_));
 OA21x2_ASAP7_75t_R _18250_ (.A1(_02549_),
    .A2(_02881_),
    .B(_02926_),
    .Y(_02213_));
 AND2x6_ASAP7_75t_R _18251_ (.A(_08102_),
    .B(_08838_),
    .Y(_02927_));
 NAND2x2_ASAP7_75t_R _18252_ (.A(_08606_),
    .B(_02927_),
    .Y(_02928_));
 BUFx6f_ASAP7_75t_R _18253_ (.A(_02928_),
    .Y(_02929_));
 NAND2x2_ASAP7_75t_R _18254_ (.A(_08937_),
    .B(_02927_),
    .Y(_02930_));
 NAND2x2_ASAP7_75t_R _18255_ (.A(_08102_),
    .B(_08847_),
    .Y(_02931_));
 NAND2x1_ASAP7_75t_R _18256_ (.A(_00009_),
    .B(_02931_),
    .Y(_02932_));
 OA21x2_ASAP7_75t_R _18257_ (.A1(_08793_),
    .A2(_02930_),
    .B(_02932_),
    .Y(_02933_));
 OA21x2_ASAP7_75t_R _18258_ (.A1(_08092_),
    .A2(_02929_),
    .B(_02933_),
    .Y(_02214_));
 BUFx12f_ASAP7_75t_R _18259_ (.A(_02931_),
    .Y(_02934_));
 AND3x2_ASAP7_75t_R _18260_ (.A(_08146_),
    .B(_08113_),
    .C(_08847_),
    .Y(_02935_));
 BUFx12f_ASAP7_75t_R _18261_ (.A(_02935_),
    .Y(_02936_));
 AOI22x1_ASAP7_75t_R _18262_ (.A1(_00741_),
    .A2(_02934_),
    .B1(_02936_),
    .B2(_08155_),
    .Y(_02937_));
 OA21x2_ASAP7_75t_R _18263_ (.A1(_02480_),
    .A2(_02929_),
    .B(_02937_),
    .Y(_02215_));
 AOI22x1_ASAP7_75t_R _18264_ (.A1(_00708_),
    .A2(_02934_),
    .B1(_02936_),
    .B2(_08184_),
    .Y(_02938_));
 OA21x2_ASAP7_75t_R _18265_ (.A1(_02485_),
    .A2(_02929_),
    .B(_02938_),
    .Y(_02216_));
 INVx1_ASAP7_75t_R _18266_ (.A(_00675_),
    .Y(_02939_));
 OA222x2_ASAP7_75t_R _18267_ (.A1(_02939_),
    .A2(_02927_),
    .B1(_02928_),
    .B2(_02488_),
    .C1(_02930_),
    .C2(_08190_),
    .Y(_02217_));
 INVx1_ASAP7_75t_R _18268_ (.A(_00642_),
    .Y(_02940_));
 OA222x2_ASAP7_75t_R _18269_ (.A1(_02940_),
    .A2(_02927_),
    .B1(_02928_),
    .B2(_02490_),
    .C1(_02930_),
    .C2(_08210_),
    .Y(_02218_));
 AOI22x1_ASAP7_75t_R _18270_ (.A1(_00609_),
    .A2(_02934_),
    .B1(_02936_),
    .B2(_08242_),
    .Y(_02941_));
 OA21x2_ASAP7_75t_R _18271_ (.A1(_02491_),
    .A2(_02929_),
    .B(_02941_),
    .Y(_02219_));
 AOI22x1_ASAP7_75t_R _18272_ (.A1(_00575_),
    .A2(_02934_),
    .B1(_02936_),
    .B2(_08258_),
    .Y(_02942_));
 OA21x2_ASAP7_75t_R _18273_ (.A1(_02493_),
    .A2(_02929_),
    .B(_02942_),
    .Y(_02220_));
 AOI22x1_ASAP7_75t_R _18274_ (.A1(_00542_),
    .A2(_02934_),
    .B1(_02936_),
    .B2(_08286_),
    .Y(_02943_));
 OA21x2_ASAP7_75t_R _18275_ (.A1(_02495_),
    .A2(_02929_),
    .B(_02943_),
    .Y(_02221_));
 BUFx12f_ASAP7_75t_R _18276_ (.A(_02931_),
    .Y(_02944_));
 AOI22x1_ASAP7_75t_R _18277_ (.A1(_00509_),
    .A2(_02944_),
    .B1(_02936_),
    .B2(_08307_),
    .Y(_02945_));
 OA21x2_ASAP7_75t_R _18278_ (.A1(_02497_),
    .A2(_02929_),
    .B(_02945_),
    .Y(_02222_));
 AOI22x1_ASAP7_75t_R _18279_ (.A1(_00476_),
    .A2(_02944_),
    .B1(_02936_),
    .B2(_08326_),
    .Y(_02946_));
 OA21x2_ASAP7_75t_R _18280_ (.A1(_02500_),
    .A2(_02929_),
    .B(_02946_),
    .Y(_02223_));
 AOI22x1_ASAP7_75t_R _18281_ (.A1(_00443_),
    .A2(_02944_),
    .B1(_02936_),
    .B2(_08347_),
    .Y(_02947_));
 OA21x2_ASAP7_75t_R _18282_ (.A1(_02502_),
    .A2(_02929_),
    .B(_02947_),
    .Y(_02224_));
 NAND2x1_ASAP7_75t_R _18283_ (.A(_01041_),
    .B(_02934_),
    .Y(_02948_));
 OA21x2_ASAP7_75t_R _18284_ (.A1(_02504_),
    .A2(_02934_),
    .B(_02948_),
    .Y(_02225_));
 AOI22x1_ASAP7_75t_R _18285_ (.A1(_00410_),
    .A2(_02944_),
    .B1(_02936_),
    .B2(_08381_),
    .Y(_02949_));
 OA21x2_ASAP7_75t_R _18286_ (.A1(_02506_),
    .A2(_02929_),
    .B(_02949_),
    .Y(_02226_));
 BUFx6f_ASAP7_75t_R _18287_ (.A(_02931_),
    .Y(_02950_));
 NAND2x1_ASAP7_75t_R _18288_ (.A(_00377_),
    .B(_02950_),
    .Y(_02951_));
 OA221x2_ASAP7_75t_R _18289_ (.A1(_08400_),
    .A2(_02934_),
    .B1(_02928_),
    .B2(_02508_),
    .C(_02951_),
    .Y(_02227_));
 BUFx4f_ASAP7_75t_R _18290_ (.A(_02928_),
    .Y(_02952_));
 BUFx6f_ASAP7_75t_R _18291_ (.A(_02935_),
    .Y(_02953_));
 AOI22x1_ASAP7_75t_R _18292_ (.A1(_00344_),
    .A2(_02944_),
    .B1(_02953_),
    .B2(_08419_),
    .Y(_02954_));
 OA21x2_ASAP7_75t_R _18293_ (.A1(_02511_),
    .A2(_02952_),
    .B(_02954_),
    .Y(_02228_));
 AOI22x1_ASAP7_75t_R _18294_ (.A1(_00310_),
    .A2(_02944_),
    .B1(_02953_),
    .B2(_08437_),
    .Y(_02955_));
 OA21x2_ASAP7_75t_R _18295_ (.A1(_02515_),
    .A2(_02952_),
    .B(_02955_),
    .Y(_02229_));
 AOI22x1_ASAP7_75t_R _18296_ (.A1(_00277_),
    .A2(_02944_),
    .B1(_02953_),
    .B2(_08458_),
    .Y(_02956_));
 OA21x2_ASAP7_75t_R _18297_ (.A1(_02517_),
    .A2(_02952_),
    .B(_02956_),
    .Y(_02230_));
 AOI22x1_ASAP7_75t_R _18298_ (.A1(_00244_),
    .A2(_02944_),
    .B1(_02953_),
    .B2(_08476_),
    .Y(_02957_));
 OA21x2_ASAP7_75t_R _18299_ (.A1(_02519_),
    .A2(_02952_),
    .B(_02957_),
    .Y(_02231_));
 AOI22x1_ASAP7_75t_R _18300_ (.A1(_00210_),
    .A2(_02944_),
    .B1(_02953_),
    .B2(_08494_),
    .Y(_02958_));
 OA21x2_ASAP7_75t_R _18301_ (.A1(_02521_),
    .A2(_02952_),
    .B(_02958_),
    .Y(_02232_));
 AOI22x1_ASAP7_75t_R _18302_ (.A1(_00177_),
    .A2(_02944_),
    .B1(_02953_),
    .B2(_08511_),
    .Y(_02959_));
 OA21x2_ASAP7_75t_R _18303_ (.A1(_02523_),
    .A2(_02952_),
    .B(_02959_),
    .Y(_02233_));
 INVx1_ASAP7_75t_R _18304_ (.A(_00143_),
    .Y(_02960_));
 OA222x2_ASAP7_75t_R _18305_ (.A1(_02960_),
    .A2(_02927_),
    .B1(_02928_),
    .B2(_02525_),
    .C1(_02930_),
    .C2(_08517_),
    .Y(_02234_));
 AOI22x1_ASAP7_75t_R _18306_ (.A1(_00110_),
    .A2(_02950_),
    .B1(_02953_),
    .B2(_08545_),
    .Y(_02961_));
 OA21x2_ASAP7_75t_R _18307_ (.A1(_02526_),
    .A2(_02952_),
    .B(_02961_),
    .Y(_02235_));
 NOR2x1_ASAP7_75t_R _18308_ (.A(_01008_),
    .B(_02927_),
    .Y(_02962_));
 AO21x1_ASAP7_75t_R _18309_ (.A1(_02528_),
    .A2(_02927_),
    .B(_02962_),
    .Y(_02236_));
 AND3x1_ASAP7_75t_R _18310_ (.A(_08146_),
    .B(_08106_),
    .C(_08873_),
    .Y(_02963_));
 NOR2x1_ASAP7_75t_R _18311_ (.A(_00076_),
    .B(_02927_),
    .Y(_02964_));
 AO221x1_ASAP7_75t_R _18312_ (.A1(_02454_),
    .A2(_02927_),
    .B1(_02963_),
    .B2(_02531_),
    .C(_02964_),
    .Y(_02237_));
 AND2x2_ASAP7_75t_R _18313_ (.A(_00044_),
    .B(_02950_),
    .Y(_02965_));
 AOI221x1_ASAP7_75t_R _18314_ (.A1(_08590_),
    .A2(_02963_),
    .B1(_02936_),
    .B2(_02533_),
    .C(_02965_),
    .Y(_02238_));
 AOI22x1_ASAP7_75t_R _18315_ (.A1(_00975_),
    .A2(_02950_),
    .B1(_02953_),
    .B2(_08603_),
    .Y(_02966_));
 OA21x2_ASAP7_75t_R _18316_ (.A1(_02535_),
    .A2(_02952_),
    .B(_02966_),
    .Y(_02239_));
 NAND2x1_ASAP7_75t_R _18317_ (.A(_00942_),
    .B(_02950_),
    .Y(_02967_));
 OA221x2_ASAP7_75t_R _18318_ (.A1(_02537_),
    .A2(_02934_),
    .B1(_02928_),
    .B2(_08618_),
    .C(_02967_),
    .Y(_02240_));
 NAND2x1_ASAP7_75t_R _18319_ (.A(_00908_),
    .B(_02950_),
    .Y(_02968_));
 OA221x2_ASAP7_75t_R _18320_ (.A1(_08630_),
    .A2(_02934_),
    .B1(_02928_),
    .B2(_02539_),
    .C(_02968_),
    .Y(_02241_));
 AOI22x1_ASAP7_75t_R _18321_ (.A1(_00875_),
    .A2(_02950_),
    .B1(_02953_),
    .B2(_08643_),
    .Y(_02969_));
 OA21x2_ASAP7_75t_R _18322_ (.A1(_02541_),
    .A2(_02952_),
    .B(_02969_),
    .Y(_02242_));
 AO21x1_ASAP7_75t_R _18323_ (.A1(_08146_),
    .A2(_08873_),
    .B(_06194_),
    .Y(_02970_));
 OA21x2_ASAP7_75t_R _18324_ (.A1(_02544_),
    .A2(_02950_),
    .B(_02970_),
    .Y(_02971_));
 OA21x2_ASAP7_75t_R _18325_ (.A1(_02543_),
    .A2(_02952_),
    .B(_02971_),
    .Y(_02243_));
 AOI22x1_ASAP7_75t_R _18326_ (.A1(_00808_),
    .A2(_02950_),
    .B1(_02953_),
    .B2(_08669_),
    .Y(_02972_));
 OA21x2_ASAP7_75t_R _18327_ (.A1(_02547_),
    .A2(_02928_),
    .B(_02972_),
    .Y(_02244_));
 NAND2x1_ASAP7_75t_R _18328_ (.A(_00774_),
    .B(_02931_),
    .Y(_02973_));
 OA21x2_ASAP7_75t_R _18329_ (.A1(_02550_),
    .A2(_02950_),
    .B(_02973_),
    .Y(_02974_));
 OA21x2_ASAP7_75t_R _18330_ (.A1(_02549_),
    .A2(_02928_),
    .B(_02974_),
    .Y(_02245_));
 BUFx4f_ASAP7_75t_R _18331_ (.A(_08069_),
    .Y(_02975_));
 AO21x1_ASAP7_75t_R _18332_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08138_),
    .Y(_02976_));
 OA21x2_ASAP7_75t_R _18333_ (.A1(_02975_),
    .A2(_08126_),
    .B(_02976_),
    .Y(\riscv.dp.ISRmux.d0[10] ));
 AO21x1_ASAP7_75t_R _18334_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08174_),
    .Y(_02977_));
 OA21x2_ASAP7_75t_R _18335_ (.A1(_02975_),
    .A2(_08161_),
    .B(_02977_),
    .Y(\riscv.dp.ISRmux.d0[11] ));
 AO21x1_ASAP7_75t_R _18336_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08200_),
    .Y(_02978_));
 OA21x2_ASAP7_75t_R _18337_ (.A1(_02975_),
    .A2(_08193_),
    .B(_02978_),
    .Y(\riscv.dp.ISRmux.d0[12] ));
 AO21x1_ASAP7_75t_R _18338_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08220_),
    .Y(_02979_));
 OA21x2_ASAP7_75t_R _18339_ (.A1(_02975_),
    .A2(_08215_),
    .B(_02979_),
    .Y(\riscv.dp.ISRmux.d0[13] ));
 AO21x1_ASAP7_75t_R _18340_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08236_),
    .Y(_02980_));
 OA21x2_ASAP7_75t_R _18341_ (.A1(_02975_),
    .A2(_08227_),
    .B(_02980_),
    .Y(\riscv.dp.ISRmux.d0[14] ));
 AO21x1_ASAP7_75t_R _18342_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08252_),
    .Y(_02981_));
 OA21x2_ASAP7_75t_R _18343_ (.A1(_02975_),
    .A2(_08246_),
    .B(_02981_),
    .Y(\riscv.dp.ISRmux.d0[15] ));
 AO21x1_ASAP7_75t_R _18344_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08274_),
    .Y(_02982_));
 OA21x2_ASAP7_75t_R _18345_ (.A1(_02975_),
    .A2(_08263_),
    .B(_02982_),
    .Y(\riscv.dp.ISRmux.d0[16] ));
 AO21x1_ASAP7_75t_R _18346_ (.A1(_08071_),
    .A2(_08072_),
    .B(_08297_),
    .Y(_02983_));
 OA21x2_ASAP7_75t_R _18347_ (.A1(_02975_),
    .A2(_08291_),
    .B(_02983_),
    .Y(\riscv.dp.ISRmux.d0[17] ));
 BUFx3_ASAP7_75t_R _18348_ (.A(_08064_),
    .Y(_02984_));
 BUFx3_ASAP7_75t_R _18349_ (.A(_08068_),
    .Y(_02985_));
 AO21x1_ASAP7_75t_R _18350_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08318_),
    .Y(_02986_));
 OA21x2_ASAP7_75t_R _18351_ (.A1(_02975_),
    .A2(_08311_),
    .B(_02986_),
    .Y(\riscv.dp.ISRmux.d0[18] ));
 BUFx3_ASAP7_75t_R _18352_ (.A(_08069_),
    .Y(_02987_));
 AO21x1_ASAP7_75t_R _18353_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08339_),
    .Y(_02988_));
 OA21x2_ASAP7_75t_R _18354_ (.A1(_02987_),
    .A2(_08332_),
    .B(_02988_),
    .Y(\riscv.dp.ISRmux.d0[19] ));
 AO21x1_ASAP7_75t_R _18355_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08373_),
    .Y(_02989_));
 OA21x2_ASAP7_75t_R _18356_ (.A1(_02987_),
    .A2(_08367_),
    .B(_02989_),
    .Y(\riscv.dp.ISRmux.d0[20] ));
 AO21x1_ASAP7_75t_R _18357_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08392_),
    .Y(_02990_));
 OA21x2_ASAP7_75t_R _18358_ (.A1(_02987_),
    .A2(_08385_),
    .B(_02990_),
    .Y(\riscv.dp.ISRmux.d0[21] ));
 AO21x1_ASAP7_75t_R _18359_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08411_),
    .Y(_02991_));
 OA21x2_ASAP7_75t_R _18360_ (.A1(_02987_),
    .A2(_08405_),
    .B(_02991_),
    .Y(\riscv.dp.ISRmux.d0[22] ));
 AO21x1_ASAP7_75t_R _18361_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08430_),
    .Y(_02992_));
 OA21x2_ASAP7_75t_R _18362_ (.A1(_02987_),
    .A2(_08425_),
    .B(_02992_),
    .Y(\riscv.dp.ISRmux.d0[23] ));
 AO21x1_ASAP7_75t_R _18363_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08451_),
    .Y(_02993_));
 OA21x2_ASAP7_75t_R _18364_ (.A1(_02987_),
    .A2(_08442_),
    .B(_02993_),
    .Y(\riscv.dp.ISRmux.d0[24] ));
 AO21x1_ASAP7_75t_R _18365_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08468_),
    .Y(_02994_));
 OA21x2_ASAP7_75t_R _18366_ (.A1(_02987_),
    .A2(_08462_),
    .B(_02994_),
    .Y(\riscv.dp.ISRmux.d0[25] ));
 AO21x1_ASAP7_75t_R _18367_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08487_),
    .Y(_02995_));
 OA21x2_ASAP7_75t_R _18368_ (.A1(_02987_),
    .A2(_08480_),
    .B(_02995_),
    .Y(\riscv.dp.ISRmux.d0[26] ));
 AO21x1_ASAP7_75t_R _18369_ (.A1(_02984_),
    .A2(_02985_),
    .B(_08504_),
    .Y(_02996_));
 OA21x2_ASAP7_75t_R _18370_ (.A1(_02987_),
    .A2(_08499_),
    .B(_02996_),
    .Y(\riscv.dp.ISRmux.d0[27] ));
 BUFx3_ASAP7_75t_R _18371_ (.A(_08064_),
    .Y(_02997_));
 BUFx3_ASAP7_75t_R _18372_ (.A(_08068_),
    .Y(_02998_));
 AO21x1_ASAP7_75t_R _18373_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08526_),
    .Y(_02999_));
 OA21x2_ASAP7_75t_R _18374_ (.A1(_02987_),
    .A2(_08528_),
    .B(_02999_),
    .Y(\riscv.dp.ISRmux.d0[28] ));
 AO21x1_ASAP7_75t_R _18375_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08538_),
    .Y(_03000_));
 OA21x2_ASAP7_75t_R _18376_ (.A1(_08070_),
    .A2(_08533_),
    .B(_03000_),
    .Y(\riscv.dp.ISRmux.d0[29] ));
 AO21x1_ASAP7_75t_R _18377_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08548_),
    .Y(_03001_));
 OA21x2_ASAP7_75t_R _18378_ (.A1(_09717_),
    .A2(_08069_),
    .B(_03001_),
    .Y(\riscv.dp.ISRmux.d0[2] ));
 AO21x1_ASAP7_75t_R _18379_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08572_),
    .Y(_03002_));
 OA21x2_ASAP7_75t_R _18380_ (.A1(_08070_),
    .A2(_08567_),
    .B(_03002_),
    .Y(\riscv.dp.ISRmux.d0[30] ));
 AO21x1_ASAP7_75t_R _18381_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08587_),
    .Y(_03003_));
 OA21x2_ASAP7_75t_R _18382_ (.A1(_08070_),
    .A2(_08581_),
    .B(_03003_),
    .Y(\riscv.dp.ISRmux.d0[31] ));
 AND3x1_ASAP7_75t_R _18383_ (.A(_01217_),
    .B(_08064_),
    .C(_08068_),
    .Y(_03004_));
 AOI21x1_ASAP7_75t_R _18384_ (.A1(_02975_),
    .A2(_08597_),
    .B(_03004_),
    .Y(\riscv.dp.ISRmux.d0[3] ));
 AO21x1_ASAP7_75t_R _18385_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08612_),
    .Y(_03005_));
 OA21x2_ASAP7_75t_R _18386_ (.A1(_08070_),
    .A2(_08610_),
    .B(_03005_),
    .Y(\riscv.dp.ISRmux.d0[4] ));
 AO21x1_ASAP7_75t_R _18387_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08624_),
    .Y(_03006_));
 OA21x2_ASAP7_75t_R _18388_ (.A1(_08070_),
    .A2(_08621_),
    .B(_03006_),
    .Y(\riscv.dp.ISRmux.d0[5] ));
 AO21x1_ASAP7_75t_R _18389_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08637_),
    .Y(_03007_));
 OA21x2_ASAP7_75t_R _18390_ (.A1(_08070_),
    .A2(_08633_),
    .B(_03007_),
    .Y(\riscv.dp.ISRmux.d0[6] ));
 AND3x1_ASAP7_75t_R _18391_ (.A(_08064_),
    .B(_08068_),
    .C(_08647_),
    .Y(_03008_));
 AO21x1_ASAP7_75t_R _18392_ (.A1(_08069_),
    .A2(_08650_),
    .B(_03008_),
    .Y(\riscv.dp.ISRmux.d0[7] ));
 AO21x1_ASAP7_75t_R _18393_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08663_),
    .Y(_03009_));
 OA21x2_ASAP7_75t_R _18394_ (.A1(_08070_),
    .A2(_08660_),
    .B(_03009_),
    .Y(\riscv.dp.ISRmux.d0[8] ));
 AO21x1_ASAP7_75t_R _18395_ (.A1(_02997_),
    .A2(_02998_),
    .B(_08676_),
    .Y(_03010_));
 OA21x2_ASAP7_75t_R _18396_ (.A1(_08070_),
    .A2(_08673_),
    .B(_03010_),
    .Y(\riscv.dp.ISRmux.d0[9] ));
 NAND2x1_ASAP7_75t_R _18397_ (.A(_03202_),
    .B(_03210_),
    .Y(_03011_));
 AND2x2_ASAP7_75t_R _18398_ (.A(_03199_),
    .B(_03011_),
    .Y(net98));
 AND3x4_ASAP7_75t_R _18399_ (.A(_03218_),
    .B(net64),
    .C(_06942_),
    .Y(_03012_));
 NOR2x2_ASAP7_75t_R _18400_ (.A(_05917_),
    .B(_03012_),
    .Y(net100));
 NOR2x2_ASAP7_75t_R _18401_ (.A(_05829_),
    .B(_03012_),
    .Y(net101));
 OR3x4_ASAP7_75t_R _18402_ (.A(_08049_),
    .B(_03229_),
    .C(_05468_),
    .Y(_03013_));
 AND2x6_ASAP7_75t_R _18403_ (.A(_05715_),
    .B(_03013_),
    .Y(net102));
 AND2x6_ASAP7_75t_R _18404_ (.A(_05610_),
    .B(_03013_),
    .Y(net103));
 AND2x6_ASAP7_75t_R _18405_ (.A(_05518_),
    .B(_03013_),
    .Y(net104));
 AND2x6_ASAP7_75t_R _18406_ (.A(_05417_),
    .B(_03013_),
    .Y(net105));
 AND2x6_ASAP7_75t_R _18407_ (.A(net64),
    .B(_06942_),
    .Y(_03014_));
 BUFx16f_ASAP7_75t_R _18408_ (.A(_03014_),
    .Y(_03015_));
 NOR2x2_ASAP7_75t_R _18409_ (.A(_07962_),
    .B(_03015_),
    .Y(net106));
 NOR2x2_ASAP7_75t_R _18410_ (.A(_05194_),
    .B(_03015_),
    .Y(net107));
 NOR2x2_ASAP7_75t_R _18411_ (.A(_05091_),
    .B(_03015_),
    .Y(net108));
 NOR2x2_ASAP7_75t_R _18412_ (.A(_04976_),
    .B(_03015_),
    .Y(net109));
 NOR2x2_ASAP7_75t_R _18413_ (.A(_04877_),
    .B(_03015_),
    .Y(net111));
 NOR2x2_ASAP7_75t_R _18414_ (.A(_04763_),
    .B(_03015_),
    .Y(net112));
 NOR2x2_ASAP7_75t_R _18415_ (.A(_04656_),
    .B(_03015_),
    .Y(net113));
 NOR2x2_ASAP7_75t_R _18416_ (.A(_04544_),
    .B(_03015_),
    .Y(net114));
 NOR2x2_ASAP7_75t_R _18417_ (.A(_04421_),
    .B(_03015_),
    .Y(net115));
 NOR2x2_ASAP7_75t_R _18418_ (.A(_04313_),
    .B(_03015_),
    .Y(net116));
 NOR2x2_ASAP7_75t_R _18419_ (.A(_07941_),
    .B(_03014_),
    .Y(net117));
 NOR2x2_ASAP7_75t_R _18420_ (.A(_04102_),
    .B(_03014_),
    .Y(net118));
 NOR2x2_ASAP7_75t_R _18421_ (.A(_03960_),
    .B(_03014_),
    .Y(net119));
 NOR2x2_ASAP7_75t_R _18422_ (.A(_03830_),
    .B(_03014_),
    .Y(net120));
 NOR2x2_ASAP7_75t_R _18423_ (.A(_03706_),
    .B(_03014_),
    .Y(net122));
 NOR2x2_ASAP7_75t_R _18424_ (.A(_03640_),
    .B(_03014_),
    .Y(net123));
 NOR2x2_ASAP7_75t_R _18425_ (.A(_06094_),
    .B(_03012_),
    .Y(net129));
 NOR2x2_ASAP7_75t_R _18426_ (.A(_06005_),
    .B(_03012_),
    .Y(net130));
 FAx1_ASAP7_75t_R _18427_ (.SN(_01065_),
    .A(_09548_),
    .B(_09549_),
    .CI(_09550_),
    .CON(_01158_));
 FAx1_ASAP7_75t_R _18428_ (.SN(_01070_),
    .A(_09551_),
    .B(_09552_),
    .CI(_09553_),
    .CON(_01159_));
 HAxp5_ASAP7_75t_R _18429_ (.A(_09555_),
    .B(_09556_),
    .CON(_01160_),
    .SN(_00034_));
 HAxp5_ASAP7_75t_R _18430_ (.A(_09557_),
    .B(_09558_),
    .CON(_01064_),
    .SN(_09559_));
 HAxp5_ASAP7_75t_R _18431_ (.A(_09560_),
    .B(_09561_),
    .CON(_01161_),
    .SN(_01162_));
 HAxp5_ASAP7_75t_R _18432_ (.A(_09562_),
    .B(_09563_),
    .CON(_01163_),
    .SN(_09564_));
 HAxp5_ASAP7_75t_R _18433_ (.A(_09565_),
    .B(_09566_),
    .CON(_00099_),
    .SN(_00100_));
 HAxp5_ASAP7_75t_R _18434_ (.A(_09567_),
    .B(_09568_),
    .CON(_01164_),
    .SN(_09569_));
 HAxp5_ASAP7_75t_R _18435_ (.A(_09570_),
    .B(_09571_),
    .CON(_00133_),
    .SN(_01165_));
 HAxp5_ASAP7_75t_R _18436_ (.A(_09572_),
    .B(_09573_),
    .CON(_01166_),
    .SN(_09574_));
 HAxp5_ASAP7_75t_R _18437_ (.A(_09575_),
    .B(_09576_),
    .CON(_00166_),
    .SN(_00167_));
 HAxp5_ASAP7_75t_R _18438_ (.A(_09577_),
    .B(_09578_),
    .CON(_01167_),
    .SN(_09579_));
 HAxp5_ASAP7_75t_R _18439_ (.A(_09580_),
    .B(_09581_),
    .CON(_00200_),
    .SN(_01168_));
 HAxp5_ASAP7_75t_R _18440_ (.A(_09582_),
    .B(_09583_),
    .CON(_01169_),
    .SN(_09584_));
 HAxp5_ASAP7_75t_R _18441_ (.A(_09585_),
    .B(_09586_),
    .CON(_00233_),
    .SN(_00234_));
 HAxp5_ASAP7_75t_R _18442_ (.A(_09587_),
    .B(_09588_),
    .CON(_01170_),
    .SN(_09589_));
 HAxp5_ASAP7_75t_R _18443_ (.A(_09590_),
    .B(_09591_),
    .CON(_01171_),
    .SN(_00267_));
 HAxp5_ASAP7_75t_R _18444_ (.A(_09592_),
    .B(_09593_),
    .CON(_01172_),
    .SN(_09594_));
 HAxp5_ASAP7_75t_R _18445_ (.A(_09595_),
    .B(_09596_),
    .CON(_01173_),
    .SN(_00300_));
 HAxp5_ASAP7_75t_R _18446_ (.A(_09597_),
    .B(_09598_),
    .CON(_01174_),
    .SN(_09599_));
 HAxp5_ASAP7_75t_R _18447_ (.A(_09600_),
    .B(_09601_),
    .CON(_00333_),
    .SN(_00334_));
 HAxp5_ASAP7_75t_R _18448_ (.A(_09602_),
    .B(_09603_),
    .CON(_01175_),
    .SN(_09604_));
 HAxp5_ASAP7_75t_R _18449_ (.A(_09605_),
    .B(_09606_),
    .CON(_01176_),
    .SN(_00367_));
 HAxp5_ASAP7_75t_R _18450_ (.A(_09607_),
    .B(_09608_),
    .CON(_01177_),
    .SN(_09609_));
 HAxp5_ASAP7_75t_R _18451_ (.A(_09610_),
    .B(_09611_),
    .CON(_01178_),
    .SN(_00400_));
 HAxp5_ASAP7_75t_R _18452_ (.A(_09612_),
    .B(_09613_),
    .CON(_01179_),
    .SN(_09614_));
 HAxp5_ASAP7_75t_R _18453_ (.A(_09615_),
    .B(_09616_),
    .CON(_01180_),
    .SN(_00433_));
 HAxp5_ASAP7_75t_R _18454_ (.A(_09617_),
    .B(_09618_),
    .CON(_01181_),
    .SN(_09619_));
 HAxp5_ASAP7_75t_R _18455_ (.A(_09620_),
    .B(_09621_),
    .CON(_01182_),
    .SN(_00466_));
 HAxp5_ASAP7_75t_R _18456_ (.A(_09622_),
    .B(_09623_),
    .CON(_01183_),
    .SN(_09624_));
 HAxp5_ASAP7_75t_R _18457_ (.A(_09625_),
    .B(_09626_),
    .CON(_01184_),
    .SN(_00499_));
 HAxp5_ASAP7_75t_R _18458_ (.A(_09627_),
    .B(_09628_),
    .CON(_01185_),
    .SN(_09629_));
 HAxp5_ASAP7_75t_R _18459_ (.A(_09630_),
    .B(_09631_),
    .CON(_01186_),
    .SN(_00532_));
 HAxp5_ASAP7_75t_R _18460_ (.A(_09632_),
    .B(_09633_),
    .CON(_01187_),
    .SN(_09634_));
 HAxp5_ASAP7_75t_R _18461_ (.A(_09635_),
    .B(_09636_),
    .CON(_01188_),
    .SN(_00565_));
 HAxp5_ASAP7_75t_R _18462_ (.A(_09637_),
    .B(_09638_),
    .CON(_01189_),
    .SN(_09639_));
 HAxp5_ASAP7_75t_R _18463_ (.A(_09640_),
    .B(_09641_),
    .CON(_00598_),
    .SN(_00599_));
 HAxp5_ASAP7_75t_R _18464_ (.A(_09642_),
    .B(_09643_),
    .CON(_01190_),
    .SN(_09644_));
 HAxp5_ASAP7_75t_R _18465_ (.A(_09645_),
    .B(_09646_),
    .CON(_01191_),
    .SN(_00632_));
 HAxp5_ASAP7_75t_R _18466_ (.A(_09647_),
    .B(_09648_),
    .CON(_01192_),
    .SN(_09649_));
 HAxp5_ASAP7_75t_R _18467_ (.A(_09650_),
    .B(_09651_),
    .CON(_01193_),
    .SN(_00665_));
 HAxp5_ASAP7_75t_R _18468_ (.A(_09652_),
    .B(_09653_),
    .CON(_01194_),
    .SN(_09654_));
 HAxp5_ASAP7_75t_R _18469_ (.A(_09655_),
    .B(_09656_),
    .CON(_01195_),
    .SN(_00698_));
 HAxp5_ASAP7_75t_R _18470_ (.A(_09657_),
    .B(_09658_),
    .CON(_01196_),
    .SN(_09659_));
 HAxp5_ASAP7_75t_R _18471_ (.A(_09660_),
    .B(_09661_),
    .CON(_01197_),
    .SN(_00731_));
 HAxp5_ASAP7_75t_R _18472_ (.A(_09662_),
    .B(_09663_),
    .CON(_01198_),
    .SN(_09664_));
 HAxp5_ASAP7_75t_R _18473_ (.A(_09665_),
    .B(_09666_),
    .CON(_01199_),
    .SN(_00764_));
 HAxp5_ASAP7_75t_R _18474_ (.A(_09667_),
    .B(_09668_),
    .CON(_01200_),
    .SN(_09669_));
 HAxp5_ASAP7_75t_R _18475_ (.A(_09670_),
    .B(_09671_),
    .CON(_00797_),
    .SN(_00798_));
 HAxp5_ASAP7_75t_R _18476_ (.A(_09672_),
    .B(_09673_),
    .CON(_01201_),
    .SN(_09674_));
 HAxp5_ASAP7_75t_R _18477_ (.A(_09675_),
    .B(_09676_),
    .CON(_01202_),
    .SN(_00831_));
 HAxp5_ASAP7_75t_R _18478_ (.A(_09677_),
    .B(_09678_),
    .CON(_01203_),
    .SN(_09679_));
 HAxp5_ASAP7_75t_R _18479_ (.A(_09680_),
    .B(_09681_),
    .CON(_00864_),
    .SN(_00865_));
 HAxp5_ASAP7_75t_R _18480_ (.A(_09682_),
    .B(_09683_),
    .CON(_01204_),
    .SN(_09684_));
 HAxp5_ASAP7_75t_R _18481_ (.A(_09685_),
    .B(_09686_),
    .CON(_01205_),
    .SN(_00898_));
 HAxp5_ASAP7_75t_R _18482_ (.A(_09687_),
    .B(_09688_),
    .CON(_01206_),
    .SN(_09689_));
 HAxp5_ASAP7_75t_R _18483_ (.A(_09690_),
    .B(_09691_),
    .CON(_00931_),
    .SN(_00932_));
 HAxp5_ASAP7_75t_R _18484_ (.A(_09692_),
    .B(_09693_),
    .CON(_01207_),
    .SN(_09694_));
 HAxp5_ASAP7_75t_R _18485_ (.A(_09695_),
    .B(_09696_),
    .CON(_01208_),
    .SN(_00965_));
 HAxp5_ASAP7_75t_R _18486_ (.A(_09697_),
    .B(_09698_),
    .CON(_01209_),
    .SN(_09699_));
 HAxp5_ASAP7_75t_R _18487_ (.A(_09700_),
    .B(_09701_),
    .CON(_01210_),
    .SN(_00998_));
 HAxp5_ASAP7_75t_R _18488_ (.A(_09702_),
    .B(_09703_),
    .CON(_01211_),
    .SN(_09704_));
 HAxp5_ASAP7_75t_R _18489_ (.A(_09706_),
    .B(_09705_),
    .CON(_01212_),
    .SN(_01031_));
 HAxp5_ASAP7_75t_R _18490_ (.A(_09707_),
    .B(_09708_),
    .CON(_01213_),
    .SN(_09709_));
 HAxp5_ASAP7_75t_R _18491_ (.A(_09549_),
    .B(_09550_),
    .CON(_01214_),
    .SN(_01215_));
 HAxp5_ASAP7_75t_R _18492_ (.A(_09710_),
    .B(_09711_),
    .CON(_01216_),
    .SN(_09712_));
 HAxp5_ASAP7_75t_R _18493_ (.A(_09713_),
    .B(_09714_),
    .CON(_09554_),
    .SN(_01067_));
 HAxp5_ASAP7_75t_R _18494_ (.A(_09552_),
    .B(_09553_),
    .CON(_01072_),
    .SN(_01069_));
 HAxp5_ASAP7_75t_R _18495_ (.A(_09715_),
    .B(_09716_),
    .CON(_01074_),
    .SN(_01071_));
 HAxp5_ASAP7_75t_R _18496_ (.A(_09717_),
    .B(_09718_),
    .CON(_00032_),
    .SN(_01217_));
 HAxp5_ASAP7_75t_R _18497_ (.A(net87),
    .B(_09718_),
    .CON(_00033_),
    .SN(_09719_));
 HAxp5_ASAP7_75t_R _18498_ (.A(net87),
    .B(net90),
    .CON(_01218_),
    .SN(_09720_));
 HAxp5_ASAP7_75t_R _18499_ (.A(_09721_),
    .B(_09722_),
    .CON(_01077_),
    .SN(_01073_));
 HAxp5_ASAP7_75t_R _18500_ (.A(_09723_),
    .B(_09724_),
    .CON(_01080_),
    .SN(_01076_));
 HAxp5_ASAP7_75t_R _18501_ (.A(_09725_),
    .B(_09726_),
    .CON(_01083_),
    .SN(_01079_));
 HAxp5_ASAP7_75t_R _18502_ (.A(_09727_),
    .B(_09728_),
    .CON(_01086_),
    .SN(_01082_));
 HAxp5_ASAP7_75t_R _18503_ (.A(_09729_),
    .B(_09730_),
    .CON(_01089_),
    .SN(_01085_));
 HAxp5_ASAP7_75t_R _18504_ (.A(_09731_),
    .B(_09732_),
    .CON(_01092_),
    .SN(_01088_));
 HAxp5_ASAP7_75t_R _18505_ (.A(_09733_),
    .B(_09734_),
    .CON(_01095_),
    .SN(_01091_));
 HAxp5_ASAP7_75t_R _18506_ (.A(_09735_),
    .B(_09736_),
    .CON(_01098_),
    .SN(_01094_));
 HAxp5_ASAP7_75t_R _18507_ (.A(_09737_),
    .B(_09738_),
    .CON(_01101_),
    .SN(_01097_));
 HAxp5_ASAP7_75t_R _18508_ (.A(_09739_),
    .B(_09740_),
    .CON(_01104_),
    .SN(_01100_));
 HAxp5_ASAP7_75t_R _18509_ (.A(_09741_),
    .B(_09742_),
    .CON(_01107_),
    .SN(_01103_));
 HAxp5_ASAP7_75t_R _18510_ (.A(_09743_),
    .B(_09744_),
    .CON(_01110_),
    .SN(_01106_));
 HAxp5_ASAP7_75t_R _18511_ (.A(_09745_),
    .B(_09746_),
    .CON(_01113_),
    .SN(_01109_));
 HAxp5_ASAP7_75t_R _18512_ (.A(_09747_),
    .B(_09748_),
    .CON(_01116_),
    .SN(_01112_));
 HAxp5_ASAP7_75t_R _18513_ (.A(_09749_),
    .B(_09750_),
    .CON(_01119_),
    .SN(_01115_));
 HAxp5_ASAP7_75t_R _18514_ (.A(_09751_),
    .B(_09752_),
    .CON(_01122_),
    .SN(_01118_));
 HAxp5_ASAP7_75t_R _18515_ (.A(_09753_),
    .B(_09754_),
    .CON(_01125_),
    .SN(_01121_));
 HAxp5_ASAP7_75t_R _18516_ (.A(_09755_),
    .B(_09756_),
    .CON(_01128_),
    .SN(_01124_));
 HAxp5_ASAP7_75t_R _18517_ (.A(_09757_),
    .B(_09758_),
    .CON(_01131_),
    .SN(_01127_));
 HAxp5_ASAP7_75t_R _18518_ (.A(_09759_),
    .B(_09760_),
    .CON(_01134_),
    .SN(_01130_));
 HAxp5_ASAP7_75t_R _18519_ (.A(_09761_),
    .B(_09762_),
    .CON(_01137_),
    .SN(_01133_));
 HAxp5_ASAP7_75t_R _18520_ (.A(_09763_),
    .B(_09764_),
    .CON(_01140_),
    .SN(_01136_));
 HAxp5_ASAP7_75t_R _18521_ (.A(_09765_),
    .B(_09766_),
    .CON(_01143_),
    .SN(_01139_));
 HAxp5_ASAP7_75t_R _18522_ (.A(_09767_),
    .B(_09768_),
    .CON(_01146_),
    .SN(_01142_));
 HAxp5_ASAP7_75t_R _18523_ (.A(_09769_),
    .B(_09770_),
    .CON(_01149_),
    .SN(_01145_));
 HAxp5_ASAP7_75t_R _18524_ (.A(_09771_),
    .B(_09772_),
    .CON(_01152_),
    .SN(_01148_));
 HAxp5_ASAP7_75t_R _18525_ (.A(_09773_),
    .B(_09774_),
    .CON(_01155_),
    .SN(_01151_));
 HAxp5_ASAP7_75t_R _18526_ (.A(_09775_),
    .B(_09776_),
    .CON(_01156_),
    .SN(_01154_));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_0_clk));
 BUFx2_ASAP7_75t_R _18528_ (.A(valid),
    .Y(net97));
 BUFx6f_ASAP7_75t_R \dmem/_153_  (.A(net38),
    .Y(\dmem/_000_ ));
 BUFx3_ASAP7_75t_R \dmem/_154_  (.A(net47),
    .Y(\dmem/_001_ ));
 BUFx6f_ASAP7_75t_R \dmem/_155_  (.A(net56),
    .Y(\dmem/_002_ ));
 OR3x4_ASAP7_75t_R \dmem/_156_  (.A(\dmem/_000_ ),
    .B(\dmem/_001_ ),
    .C(\dmem/_002_ ),
    .Y(\dmem/_003_ ));
 CKINVDCx6p67_ASAP7_75t_R \dmem/_157_  (.A(\dmem/_003_ ),
    .Y(\dmem/ce_mem[0] ));
 BUFx6f_ASAP7_75t_R \dmem/_158_  (.A(\dmem/_000_ ),
    .Y(\dmem/_004_ ));
 BUFx6f_ASAP7_75t_R \dmem/_159_  (.A(\dmem/_001_ ),
    .Y(\dmem/_005_ ));
 NOR2x2_ASAP7_75t_R \dmem/_160_  (.A(\dmem/_005_ ),
    .B(\dmem/_002_ ),
    .Y(\dmem/_006_ ));
 AND2x6_ASAP7_75t_R \dmem/_161_  (.A(\dmem/_004_ ),
    .B(\dmem/_006_ ),
    .Y(\dmem/ce_mem[1] ));
 BUFx6f_ASAP7_75t_R \dmem/_162_  (.A(\dmem/_001_ ),
    .Y(\dmem/_007_ ));
 BUFx6f_ASAP7_75t_R \dmem/_163_  (.A(\dmem/_007_ ),
    .Y(\dmem/_008_ ));
 INVx3_ASAP7_75t_R \dmem/_164_  (.A(\dmem/_002_ ),
    .Y(\dmem/_009_ ));
 BUFx3_ASAP7_75t_R \dmem/_165_  (.A(\dmem/_009_ ),
    .Y(\dmem/_010_ ));
 AND2x6_ASAP7_75t_R \dmem/_166_  (.A(\dmem/_008_ ),
    .B(\dmem/_010_ ),
    .Y(\dmem/ce_mem[2] ));
 BUFx3_ASAP7_75t_R \dmem/_167_  (.A(\dmem/_002_ ),
    .Y(\dmem/_011_ ));
 INVx1_ASAP7_75t_R \dmem/_168_  (.A(\dmem/inter_dmem1[0] ),
    .Y(\dmem/_012_ ));
 NOR2x1_ASAP7_75t_R \dmem/_169_  (.A(\dmem/_005_ ),
    .B(\dmem/inter_dmem2[0] ),
    .Y(\dmem/_013_ ));
 AOI22x1_ASAP7_75t_R \dmem/_170_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_012_ ),
    .B1(\dmem/_013_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_014_ ));
 BUFx6f_ASAP7_75t_R \dmem/_171_  (.A(\dmem/_003_ ),
    .Y(\dmem/_015_ ));
 OA22x2_ASAP7_75t_R \dmem/_172_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[0] ),
    .B1(\dmem/inter_dmem3[0] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_016_ ));
 OA21x2_ASAP7_75t_R \dmem/_173_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_014_ ),
    .B(\dmem/_016_ ),
    .Y(\readdata[0] ));
 INVx1_ASAP7_75t_R \dmem/_174_  (.A(\dmem/inter_dmem1[10] ),
    .Y(\dmem/_017_ ));
 NOR2x1_ASAP7_75t_R \dmem/_175_  (.A(\dmem/_005_ ),
    .B(\dmem/inter_dmem2[10] ),
    .Y(\dmem/_018_ ));
 AOI22x1_ASAP7_75t_R \dmem/_176_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_017_ ),
    .B1(\dmem/_018_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_019_ ));
 OA22x2_ASAP7_75t_R \dmem/_177_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[10] ),
    .B1(\dmem/inter_dmem3[10] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_020_ ));
 OA21x2_ASAP7_75t_R \dmem/_178_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_019_ ),
    .B(\dmem/_020_ ),
    .Y(\readdata[10] ));
 INVx1_ASAP7_75t_R \dmem/_179_  (.A(\dmem/inter_dmem1[11] ),
    .Y(\dmem/_021_ ));
 NOR2x1_ASAP7_75t_R \dmem/_180_  (.A(\dmem/_005_ ),
    .B(\dmem/inter_dmem2[11] ),
    .Y(\dmem/_022_ ));
 AOI22x1_ASAP7_75t_R \dmem/_181_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_021_ ),
    .B1(\dmem/_022_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_023_ ));
 OA22x2_ASAP7_75t_R \dmem/_182_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[11] ),
    .B1(\dmem/inter_dmem3[11] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_024_ ));
 OA21x2_ASAP7_75t_R \dmem/_183_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_023_ ),
    .B(\dmem/_024_ ),
    .Y(\readdata[11] ));
 INVx1_ASAP7_75t_R \dmem/_184_  (.A(\dmem/inter_dmem1[12] ),
    .Y(\dmem/_025_ ));
 NOR2x1_ASAP7_75t_R \dmem/_185_  (.A(\dmem/_005_ ),
    .B(\dmem/inter_dmem2[12] ),
    .Y(\dmem/_026_ ));
 AOI22x1_ASAP7_75t_R \dmem/_186_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_025_ ),
    .B1(\dmem/_026_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_027_ ));
 OA22x2_ASAP7_75t_R \dmem/_187_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[12] ),
    .B1(\dmem/inter_dmem3[12] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_028_ ));
 OA21x2_ASAP7_75t_R \dmem/_188_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_027_ ),
    .B(\dmem/_028_ ),
    .Y(\readdata[12] ));
 INVx1_ASAP7_75t_R \dmem/_189_  (.A(\dmem/inter_dmem1[13] ),
    .Y(\dmem/_029_ ));
 NOR2x1_ASAP7_75t_R \dmem/_190_  (.A(\dmem/_005_ ),
    .B(\dmem/inter_dmem2[13] ),
    .Y(\dmem/_030_ ));
 AOI22x1_ASAP7_75t_R \dmem/_191_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_029_ ),
    .B1(\dmem/_030_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_031_ ));
 OA22x2_ASAP7_75t_R \dmem/_192_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[13] ),
    .B1(\dmem/inter_dmem3[13] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_032_ ));
 OA21x2_ASAP7_75t_R \dmem/_193_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_031_ ),
    .B(\dmem/_032_ ),
    .Y(\readdata[13] ));
 INVx1_ASAP7_75t_R \dmem/_194_  (.A(\dmem/inter_dmem1[14] ),
    .Y(\dmem/_033_ ));
 BUFx6f_ASAP7_75t_R \dmem/_195_  (.A(\dmem/_001_ ),
    .Y(\dmem/_034_ ));
 NOR2x1_ASAP7_75t_R \dmem/_196_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[14] ),
    .Y(\dmem/_035_ ));
 AOI22x1_ASAP7_75t_R \dmem/_197_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_033_ ),
    .B1(\dmem/_035_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_036_ ));
 OA22x2_ASAP7_75t_R \dmem/_198_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[14] ),
    .B1(\dmem/inter_dmem3[14] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_037_ ));
 OA21x2_ASAP7_75t_R \dmem/_199_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_036_ ),
    .B(\dmem/_037_ ),
    .Y(\readdata[14] ));
 INVx1_ASAP7_75t_R \dmem/_200_  (.A(\dmem/inter_dmem1[15] ),
    .Y(\dmem/_038_ ));
 NOR2x1_ASAP7_75t_R \dmem/_201_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[15] ),
    .Y(\dmem/_039_ ));
 AOI22x1_ASAP7_75t_R \dmem/_202_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_038_ ),
    .B1(\dmem/_039_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_040_ ));
 OA22x2_ASAP7_75t_R \dmem/_203_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[15] ),
    .B1(\dmem/inter_dmem3[15] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_041_ ));
 OA21x2_ASAP7_75t_R \dmem/_204_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_040_ ),
    .B(\dmem/_041_ ),
    .Y(\readdata[15] ));
 INVx1_ASAP7_75t_R \dmem/_205_  (.A(\dmem/inter_dmem1[16] ),
    .Y(\dmem/_042_ ));
 NOR2x1_ASAP7_75t_R \dmem/_206_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[16] ),
    .Y(\dmem/_043_ ));
 AOI22x1_ASAP7_75t_R \dmem/_207_  (.A1(\dmem/_008_ ),
    .A2(\dmem/_042_ ),
    .B1(\dmem/_043_ ),
    .B2(\dmem/_004_ ),
    .Y(\dmem/_044_ ));
 OA22x2_ASAP7_75t_R \dmem/_208_  (.A1(\dmem/_010_ ),
    .A2(\dmem/inter_dmem0[16] ),
    .B1(\dmem/inter_dmem3[16] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_045_ ));
 OA21x2_ASAP7_75t_R \dmem/_209_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_044_ ),
    .B(\dmem/_045_ ),
    .Y(\readdata[16] ));
 BUFx6f_ASAP7_75t_R \dmem/_210_  (.A(\dmem/_007_ ),
    .Y(\dmem/_046_ ));
 INVx1_ASAP7_75t_R \dmem/_211_  (.A(\dmem/inter_dmem1[17] ),
    .Y(\dmem/_047_ ));
 NOR2x1_ASAP7_75t_R \dmem/_212_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[17] ),
    .Y(\dmem/_048_ ));
 BUFx6f_ASAP7_75t_R \dmem/_213_  (.A(\dmem/_000_ ),
    .Y(\dmem/_049_ ));
 AOI22x1_ASAP7_75t_R \dmem/_214_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_047_ ),
    .B1(\dmem/_048_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_050_ ));
 BUFx3_ASAP7_75t_R \dmem/_215_  (.A(\dmem/_009_ ),
    .Y(\dmem/_051_ ));
 OA22x2_ASAP7_75t_R \dmem/_216_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[17] ),
    .B1(\dmem/inter_dmem3[17] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_052_ ));
 OA21x2_ASAP7_75t_R \dmem/_217_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_050_ ),
    .B(\dmem/_052_ ),
    .Y(\readdata[17] ));
 INVx1_ASAP7_75t_R \dmem/_218_  (.A(\dmem/inter_dmem1[18] ),
    .Y(\dmem/_053_ ));
 NOR2x1_ASAP7_75t_R \dmem/_219_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[18] ),
    .Y(\dmem/_054_ ));
 AOI22x1_ASAP7_75t_R \dmem/_220_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_053_ ),
    .B1(\dmem/_054_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_055_ ));
 OA22x2_ASAP7_75t_R \dmem/_221_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[18] ),
    .B1(\dmem/inter_dmem3[18] ),
    .B2(\dmem/_015_ ),
    .Y(\dmem/_056_ ));
 OA21x2_ASAP7_75t_R \dmem/_222_  (.A1(\dmem/_011_ ),
    .A2(\dmem/_055_ ),
    .B(\dmem/_056_ ),
    .Y(\readdata[18] ));
 BUFx3_ASAP7_75t_R \dmem/_223_  (.A(\dmem/_002_ ),
    .Y(\dmem/_057_ ));
 INVx1_ASAP7_75t_R \dmem/_224_  (.A(\dmem/inter_dmem1[19] ),
    .Y(\dmem/_058_ ));
 NOR2x1_ASAP7_75t_R \dmem/_225_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[19] ),
    .Y(\dmem/_059_ ));
 AOI22x1_ASAP7_75t_R \dmem/_226_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_058_ ),
    .B1(\dmem/_059_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_060_ ));
 BUFx6f_ASAP7_75t_R \dmem/_227_  (.A(\dmem/_003_ ),
    .Y(\dmem/_061_ ));
 OA22x2_ASAP7_75t_R \dmem/_228_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[19] ),
    .B1(\dmem/inter_dmem3[19] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_062_ ));
 OA21x2_ASAP7_75t_R \dmem/_229_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_060_ ),
    .B(\dmem/_062_ ),
    .Y(\readdata[19] ));
 INVx1_ASAP7_75t_R \dmem/_230_  (.A(\dmem/inter_dmem1[1] ),
    .Y(\dmem/_063_ ));
 NOR2x1_ASAP7_75t_R \dmem/_231_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[1] ),
    .Y(\dmem/_064_ ));
 AOI22x1_ASAP7_75t_R \dmem/_232_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_063_ ),
    .B1(\dmem/_064_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_065_ ));
 OA22x2_ASAP7_75t_R \dmem/_233_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[1] ),
    .B1(\dmem/inter_dmem3[1] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_066_ ));
 OA21x2_ASAP7_75t_R \dmem/_234_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_065_ ),
    .B(\dmem/_066_ ),
    .Y(\readdata[1] ));
 INVx1_ASAP7_75t_R \dmem/_235_  (.A(\dmem/inter_dmem1[20] ),
    .Y(\dmem/_067_ ));
 NOR2x1_ASAP7_75t_R \dmem/_236_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[20] ),
    .Y(\dmem/_068_ ));
 AOI22x1_ASAP7_75t_R \dmem/_237_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_067_ ),
    .B1(\dmem/_068_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_069_ ));
 OA22x2_ASAP7_75t_R \dmem/_238_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[20] ),
    .B1(\dmem/inter_dmem3[20] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_070_ ));
 OA21x2_ASAP7_75t_R \dmem/_239_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_069_ ),
    .B(\dmem/_070_ ),
    .Y(\readdata[20] ));
 INVx1_ASAP7_75t_R \dmem/_240_  (.A(\dmem/inter_dmem1[21] ),
    .Y(\dmem/_071_ ));
 NOR2x1_ASAP7_75t_R \dmem/_241_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[21] ),
    .Y(\dmem/_072_ ));
 AOI22x1_ASAP7_75t_R \dmem/_242_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_071_ ),
    .B1(\dmem/_072_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_073_ ));
 OA22x2_ASAP7_75t_R \dmem/_243_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[21] ),
    .B1(\dmem/inter_dmem3[21] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_074_ ));
 OA21x2_ASAP7_75t_R \dmem/_244_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_073_ ),
    .B(\dmem/_074_ ),
    .Y(\readdata[21] ));
 INVx1_ASAP7_75t_R \dmem/_245_  (.A(\dmem/inter_dmem1[22] ),
    .Y(\dmem/_075_ ));
 NOR2x1_ASAP7_75t_R \dmem/_246_  (.A(\dmem/_034_ ),
    .B(\dmem/inter_dmem2[22] ),
    .Y(\dmem/_076_ ));
 AOI22x1_ASAP7_75t_R \dmem/_247_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_075_ ),
    .B1(\dmem/_076_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_077_ ));
 OA22x2_ASAP7_75t_R \dmem/_248_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[22] ),
    .B1(\dmem/inter_dmem3[22] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_078_ ));
 OA21x2_ASAP7_75t_R \dmem/_249_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_077_ ),
    .B(\dmem/_078_ ),
    .Y(\readdata[22] ));
 INVx1_ASAP7_75t_R \dmem/_250_  (.A(\dmem/inter_dmem1[23] ),
    .Y(\dmem/_079_ ));
 BUFx6f_ASAP7_75t_R \dmem/_251_  (.A(\dmem/_001_ ),
    .Y(\dmem/_080_ ));
 NOR2x1_ASAP7_75t_R \dmem/_252_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[23] ),
    .Y(\dmem/_081_ ));
 AOI22x1_ASAP7_75t_R \dmem/_253_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_079_ ),
    .B1(\dmem/_081_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_082_ ));
 OA22x2_ASAP7_75t_R \dmem/_254_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[23] ),
    .B1(\dmem/inter_dmem3[23] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_083_ ));
 OA21x2_ASAP7_75t_R \dmem/_255_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_082_ ),
    .B(\dmem/_083_ ),
    .Y(\readdata[23] ));
 INVx1_ASAP7_75t_R \dmem/_256_  (.A(\dmem/inter_dmem1[24] ),
    .Y(\dmem/_084_ ));
 NOR2x1_ASAP7_75t_R \dmem/_257_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[24] ),
    .Y(\dmem/_085_ ));
 AOI22x1_ASAP7_75t_R \dmem/_258_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_084_ ),
    .B1(\dmem/_085_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_086_ ));
 OA22x2_ASAP7_75t_R \dmem/_259_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[24] ),
    .B1(\dmem/inter_dmem3[24] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_087_ ));
 OA21x2_ASAP7_75t_R \dmem/_260_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_086_ ),
    .B(\dmem/_087_ ),
    .Y(\readdata[24] ));
 INVx1_ASAP7_75t_R \dmem/_261_  (.A(\dmem/inter_dmem1[25] ),
    .Y(\dmem/_088_ ));
 NOR2x1_ASAP7_75t_R \dmem/_262_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[25] ),
    .Y(\dmem/_089_ ));
 AOI22x1_ASAP7_75t_R \dmem/_263_  (.A1(\dmem/_046_ ),
    .A2(\dmem/_088_ ),
    .B1(\dmem/_089_ ),
    .B2(\dmem/_049_ ),
    .Y(\dmem/_090_ ));
 OA22x2_ASAP7_75t_R \dmem/_264_  (.A1(\dmem/_051_ ),
    .A2(\dmem/inter_dmem0[25] ),
    .B1(\dmem/inter_dmem3[25] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_091_ ));
 OA21x2_ASAP7_75t_R \dmem/_265_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_090_ ),
    .B(\dmem/_091_ ),
    .Y(\readdata[25] ));
 BUFx6f_ASAP7_75t_R \dmem/_266_  (.A(\dmem/_007_ ),
    .Y(\dmem/_092_ ));
 INVx1_ASAP7_75t_R \dmem/_267_  (.A(\dmem/inter_dmem1[26] ),
    .Y(\dmem/_093_ ));
 NOR2x1_ASAP7_75t_R \dmem/_268_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[26] ),
    .Y(\dmem/_094_ ));
 BUFx6f_ASAP7_75t_R \dmem/_269_  (.A(\dmem/_000_ ),
    .Y(\dmem/_095_ ));
 AOI22x1_ASAP7_75t_R \dmem/_270_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_093_ ),
    .B1(\dmem/_094_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_096_ ));
 BUFx3_ASAP7_75t_R \dmem/_271_  (.A(\dmem/_009_ ),
    .Y(\dmem/_097_ ));
 OA22x2_ASAP7_75t_R \dmem/_272_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[26] ),
    .B1(\dmem/inter_dmem3[26] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_098_ ));
 OA21x2_ASAP7_75t_R \dmem/_273_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_096_ ),
    .B(\dmem/_098_ ),
    .Y(\readdata[26] ));
 INVx1_ASAP7_75t_R \dmem/_274_  (.A(\dmem/inter_dmem1[27] ),
    .Y(\dmem/_099_ ));
 NOR2x1_ASAP7_75t_R \dmem/_275_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[27] ),
    .Y(\dmem/_100_ ));
 AOI22x1_ASAP7_75t_R \dmem/_276_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_099_ ),
    .B1(\dmem/_100_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_101_ ));
 OA22x2_ASAP7_75t_R \dmem/_277_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[27] ),
    .B1(\dmem/inter_dmem3[27] ),
    .B2(\dmem/_061_ ),
    .Y(\dmem/_102_ ));
 OA21x2_ASAP7_75t_R \dmem/_278_  (.A1(\dmem/_057_ ),
    .A2(\dmem/_101_ ),
    .B(\dmem/_102_ ),
    .Y(\readdata[27] ));
 BUFx3_ASAP7_75t_R \dmem/_279_  (.A(\dmem/_002_ ),
    .Y(\dmem/_103_ ));
 INVx1_ASAP7_75t_R \dmem/_280_  (.A(\dmem/inter_dmem1[28] ),
    .Y(\dmem/_104_ ));
 NOR2x1_ASAP7_75t_R \dmem/_281_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[28] ),
    .Y(\dmem/_105_ ));
 AOI22x1_ASAP7_75t_R \dmem/_282_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_104_ ),
    .B1(\dmem/_105_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_106_ ));
 BUFx6f_ASAP7_75t_R \dmem/_283_  (.A(\dmem/_003_ ),
    .Y(\dmem/_107_ ));
 OA22x2_ASAP7_75t_R \dmem/_284_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[28] ),
    .B1(\dmem/inter_dmem3[28] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_108_ ));
 OA21x2_ASAP7_75t_R \dmem/_285_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_106_ ),
    .B(\dmem/_108_ ),
    .Y(\readdata[28] ));
 INVx1_ASAP7_75t_R \dmem/_286_  (.A(\dmem/inter_dmem1[29] ),
    .Y(\dmem/_109_ ));
 NOR2x1_ASAP7_75t_R \dmem/_287_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[29] ),
    .Y(\dmem/_110_ ));
 AOI22x1_ASAP7_75t_R \dmem/_288_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_109_ ),
    .B1(\dmem/_110_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_111_ ));
 OA22x2_ASAP7_75t_R \dmem/_289_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[29] ),
    .B1(\dmem/inter_dmem3[29] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_112_ ));
 OA21x2_ASAP7_75t_R \dmem/_290_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_111_ ),
    .B(\dmem/_112_ ),
    .Y(\readdata[29] ));
 INVx1_ASAP7_75t_R \dmem/_291_  (.A(\dmem/inter_dmem1[2] ),
    .Y(\dmem/_113_ ));
 NOR2x1_ASAP7_75t_R \dmem/_292_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[2] ),
    .Y(\dmem/_114_ ));
 AOI22x1_ASAP7_75t_R \dmem/_293_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_113_ ),
    .B1(\dmem/_114_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_115_ ));
 OA22x2_ASAP7_75t_R \dmem/_294_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[2] ),
    .B1(\dmem/inter_dmem3[2] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_116_ ));
 OA21x2_ASAP7_75t_R \dmem/_295_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_115_ ),
    .B(\dmem/_116_ ),
    .Y(\readdata[2] ));
 INVx1_ASAP7_75t_R \dmem/_296_  (.A(\dmem/inter_dmem1[30] ),
    .Y(\dmem/_117_ ));
 NOR2x1_ASAP7_75t_R \dmem/_297_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[30] ),
    .Y(\dmem/_118_ ));
 AOI22x1_ASAP7_75t_R \dmem/_298_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_117_ ),
    .B1(\dmem/_118_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_119_ ));
 OA22x2_ASAP7_75t_R \dmem/_299_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[30] ),
    .B1(\dmem/inter_dmem3[30] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_120_ ));
 OA21x2_ASAP7_75t_R \dmem/_300_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_119_ ),
    .B(\dmem/_120_ ),
    .Y(\readdata[30] ));
 INVx1_ASAP7_75t_R \dmem/_301_  (.A(\dmem/inter_dmem1[31] ),
    .Y(\dmem/_121_ ));
 NOR2x1_ASAP7_75t_R \dmem/_302_  (.A(\dmem/_080_ ),
    .B(\dmem/inter_dmem2[31] ),
    .Y(\dmem/_122_ ));
 AOI22x1_ASAP7_75t_R \dmem/_303_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_121_ ),
    .B1(\dmem/_122_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_123_ ));
 OA22x2_ASAP7_75t_R \dmem/_304_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[31] ),
    .B1(\dmem/inter_dmem3[31] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_124_ ));
 OA21x2_ASAP7_75t_R \dmem/_305_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_123_ ),
    .B(\dmem/_124_ ),
    .Y(\readdata[31] ));
 INVx1_ASAP7_75t_R \dmem/_306_  (.A(\dmem/inter_dmem1[3] ),
    .Y(\dmem/_125_ ));
 NOR2x1_ASAP7_75t_R \dmem/_307_  (.A(\dmem/_007_ ),
    .B(\dmem/inter_dmem2[3] ),
    .Y(\dmem/_126_ ));
 AOI22x1_ASAP7_75t_R \dmem/_308_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_125_ ),
    .B1(\dmem/_126_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_127_ ));
 OA22x2_ASAP7_75t_R \dmem/_309_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[3] ),
    .B1(\dmem/inter_dmem3[3] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_128_ ));
 OA21x2_ASAP7_75t_R \dmem/_310_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_127_ ),
    .B(\dmem/_128_ ),
    .Y(\readdata[3] ));
 INVx1_ASAP7_75t_R \dmem/_311_  (.A(\dmem/inter_dmem1[4] ),
    .Y(\dmem/_129_ ));
 NOR2x1_ASAP7_75t_R \dmem/_312_  (.A(\dmem/_007_ ),
    .B(\dmem/inter_dmem2[4] ),
    .Y(\dmem/_130_ ));
 AOI22x1_ASAP7_75t_R \dmem/_313_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_129_ ),
    .B1(\dmem/_130_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_131_ ));
 OA22x2_ASAP7_75t_R \dmem/_314_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[4] ),
    .B1(\dmem/inter_dmem3[4] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_132_ ));
 OA21x2_ASAP7_75t_R \dmem/_315_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_131_ ),
    .B(\dmem/_132_ ),
    .Y(\readdata[4] ));
 INVx1_ASAP7_75t_R \dmem/_316_  (.A(\dmem/inter_dmem1[5] ),
    .Y(\dmem/_133_ ));
 NOR2x1_ASAP7_75t_R \dmem/_317_  (.A(\dmem/_007_ ),
    .B(\dmem/inter_dmem2[5] ),
    .Y(\dmem/_134_ ));
 AOI22x1_ASAP7_75t_R \dmem/_318_  (.A1(\dmem/_092_ ),
    .A2(\dmem/_133_ ),
    .B1(\dmem/_134_ ),
    .B2(\dmem/_095_ ),
    .Y(\dmem/_135_ ));
 OA22x2_ASAP7_75t_R \dmem/_319_  (.A1(\dmem/_097_ ),
    .A2(\dmem/inter_dmem0[5] ),
    .B1(\dmem/inter_dmem3[5] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_136_ ));
 OA21x2_ASAP7_75t_R \dmem/_320_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_135_ ),
    .B(\dmem/_136_ ),
    .Y(\readdata[5] ));
 INVx1_ASAP7_75t_R \dmem/_321_  (.A(\dmem/inter_dmem1[6] ),
    .Y(\dmem/_137_ ));
 NOR2x1_ASAP7_75t_R \dmem/_322_  (.A(\dmem/_007_ ),
    .B(\dmem/inter_dmem2[6] ),
    .Y(\dmem/_138_ ));
 AOI22x1_ASAP7_75t_R \dmem/_323_  (.A1(\dmem/_005_ ),
    .A2(\dmem/_137_ ),
    .B1(\dmem/_138_ ),
    .B2(\dmem/_000_ ),
    .Y(\dmem/_139_ ));
 OA22x2_ASAP7_75t_R \dmem/_324_  (.A1(\dmem/_009_ ),
    .A2(\dmem/inter_dmem0[6] ),
    .B1(\dmem/inter_dmem3[6] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_140_ ));
 OA21x2_ASAP7_75t_R \dmem/_325_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_139_ ),
    .B(\dmem/_140_ ),
    .Y(\readdata[6] ));
 INVx1_ASAP7_75t_R \dmem/_326_  (.A(\dmem/inter_dmem1[7] ),
    .Y(\dmem/_141_ ));
 NOR2x1_ASAP7_75t_R \dmem/_327_  (.A(\dmem/_007_ ),
    .B(\dmem/inter_dmem2[7] ),
    .Y(\dmem/_142_ ));
 AOI22x1_ASAP7_75t_R \dmem/_328_  (.A1(\dmem/_005_ ),
    .A2(\dmem/_141_ ),
    .B1(\dmem/_142_ ),
    .B2(\dmem/_000_ ),
    .Y(\dmem/_143_ ));
 OA22x2_ASAP7_75t_R \dmem/_329_  (.A1(\dmem/_009_ ),
    .A2(\dmem/inter_dmem0[7] ),
    .B1(\dmem/inter_dmem3[7] ),
    .B2(\dmem/_107_ ),
    .Y(\dmem/_144_ ));
 OA21x2_ASAP7_75t_R \dmem/_330_  (.A1(\dmem/_103_ ),
    .A2(\dmem/_143_ ),
    .B(\dmem/_144_ ),
    .Y(\readdata[7] ));
 INVx1_ASAP7_75t_R \dmem/_331_  (.A(\dmem/inter_dmem1[8] ),
    .Y(\dmem/_145_ ));
 NOR2x1_ASAP7_75t_R \dmem/_332_  (.A(\dmem/_007_ ),
    .B(\dmem/inter_dmem2[8] ),
    .Y(\dmem/_146_ ));
 AOI22x1_ASAP7_75t_R \dmem/_333_  (.A1(\dmem/_005_ ),
    .A2(\dmem/_145_ ),
    .B1(\dmem/_146_ ),
    .B2(\dmem/_000_ ),
    .Y(\dmem/_147_ ));
 OA22x2_ASAP7_75t_R \dmem/_334_  (.A1(\dmem/_009_ ),
    .A2(\dmem/inter_dmem0[8] ),
    .B1(\dmem/inter_dmem3[8] ),
    .B2(\dmem/_003_ ),
    .Y(\dmem/_148_ ));
 OA21x2_ASAP7_75t_R \dmem/_335_  (.A1(\dmem/_002_ ),
    .A2(\dmem/_147_ ),
    .B(\dmem/_148_ ),
    .Y(\readdata[8] ));
 INVx1_ASAP7_75t_R \dmem/_336_  (.A(\dmem/inter_dmem1[9] ),
    .Y(\dmem/_149_ ));
 NOR2x1_ASAP7_75t_R \dmem/_337_  (.A(\dmem/_007_ ),
    .B(\dmem/inter_dmem2[9] ),
    .Y(\dmem/_150_ ));
 AOI22x1_ASAP7_75t_R \dmem/_338_  (.A1(\dmem/_005_ ),
    .A2(\dmem/_149_ ),
    .B1(\dmem/_150_ ),
    .B2(\dmem/_000_ ),
    .Y(\dmem/_151_ ));
 OA22x2_ASAP7_75t_R \dmem/_339_  (.A1(\dmem/_009_ ),
    .A2(\dmem/inter_dmem0[9] ),
    .B1(\dmem/inter_dmem3[9] ),
    .B2(\dmem/_003_ ),
    .Y(\dmem/_152_ ));
 OA21x2_ASAP7_75t_R \dmem/_340_  (.A1(\dmem/_002_ ),
    .A2(\dmem/_151_ ),
    .B(\dmem/_152_ ),
    .Y(\readdata[9] ));
 AND2x2_ASAP7_75t_R \dmem/_341_  (.A(net64),
    .B(\dmem/ce_mem[0] ),
    .Y(\dmem/we_mem[0] ));
 AND3x4_ASAP7_75t_R \dmem/_342_  (.A(\dmem/_004_ ),
    .B(net64),
    .C(\dmem/_006_ ),
    .Y(\dmem/we_mem[1] ));
 AND3x4_ASAP7_75t_R \dmem/_343_  (.A(\dmem/_008_ ),
    .B(\dmem/_010_ ),
    .C(net64),
    .Y(\dmem/we_mem[2] ));
 AND2x6_ASAP7_75t_R \dmem/_344_  (.A(\dmem/_002_ ),
    .B(net64),
    .Y(\dmem/we_mem[3] ));
 fakeram7_256x32 \dmem/dmem0  (.we_in(\dmem/we_mem[0] ),
    .ce_in(\dmem/ce_mem[0] ),
    .clk(clknet_2_2_0_clk),
    .addr_in({net61,
    net60,
    net59,
    net58,
    net57,
    net54,
    net43,
    net32}),
    .rd_out({\dmem/inter_dmem0[31] ,
    \dmem/inter_dmem0[30] ,
    \dmem/inter_dmem0[29] ,
    \dmem/inter_dmem0[28] ,
    \dmem/inter_dmem0[27] ,
    \dmem/inter_dmem0[26] ,
    \dmem/inter_dmem0[25] ,
    \dmem/inter_dmem0[24] ,
    \dmem/inter_dmem0[23] ,
    \dmem/inter_dmem0[22] ,
    \dmem/inter_dmem0[21] ,
    \dmem/inter_dmem0[20] ,
    \dmem/inter_dmem0[19] ,
    \dmem/inter_dmem0[18] ,
    \dmem/inter_dmem0[17] ,
    \dmem/inter_dmem0[16] ,
    \dmem/inter_dmem0[15] ,
    \dmem/inter_dmem0[14] ,
    \dmem/inter_dmem0[13] ,
    \dmem/inter_dmem0[12] ,
    \dmem/inter_dmem0[11] ,
    \dmem/inter_dmem0[10] ,
    \dmem/inter_dmem0[9] ,
    \dmem/inter_dmem0[8] ,
    \dmem/inter_dmem0[7] ,
    \dmem/inter_dmem0[6] ,
    \dmem/inter_dmem0[5] ,
    \dmem/inter_dmem0[4] ,
    \dmem/inter_dmem0[3] ,
    \dmem/inter_dmem0[2] ,
    \dmem/inter_dmem0[1] ,
    \dmem/inter_dmem0[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net4,
    net165,
    net124,
    net121,
    net110,
    net99}));
 fakeram7_256x32 \dmem/dmem1  (.we_in(\dmem/we_mem[1] ),
    .ce_in(\dmem/ce_mem[1] ),
    .clk(clknet_2_2_0_clk),
    .addr_in({net38,
    net37,
    net36,
    net35,
    net34,
    net33,
    net63,
    net62}),
    .rd_out({\dmem/inter_dmem1[31] ,
    \dmem/inter_dmem1[30] ,
    \dmem/inter_dmem1[29] ,
    \dmem/inter_dmem1[28] ,
    \dmem/inter_dmem1[27] ,
    \dmem/inter_dmem1[26] ,
    \dmem/inter_dmem1[25] ,
    \dmem/inter_dmem1[24] ,
    \dmem/inter_dmem1[23] ,
    \dmem/inter_dmem1[22] ,
    \dmem/inter_dmem1[21] ,
    \dmem/inter_dmem1[20] ,
    \dmem/inter_dmem1[19] ,
    \dmem/inter_dmem1[18] ,
    \dmem/inter_dmem1[17] ,
    \dmem/inter_dmem1[16] ,
    \dmem/inter_dmem1[15] ,
    \dmem/inter_dmem1[14] ,
    \dmem/inter_dmem1[13] ,
    \dmem/inter_dmem1[12] ,
    \dmem/inter_dmem1[11] ,
    \dmem/inter_dmem1[10] ,
    \dmem/inter_dmem1[9] ,
    \dmem/inter_dmem1[8] ,
    \dmem/inter_dmem1[7] ,
    \dmem/inter_dmem1[6] ,
    \dmem/inter_dmem1[5] ,
    \dmem/inter_dmem1[4] ,
    \dmem/inter_dmem1[3] ,
    \dmem/inter_dmem1[2] ,
    \dmem/inter_dmem1[1] ,
    \dmem/inter_dmem1[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net126,
    net166,
    net124,
    net121,
    net110,
    net99}));
 fakeram7_256x32 \dmem/dmem2  (.we_in(\dmem/we_mem[2] ),
    .ce_in(\dmem/ce_mem[2] ),
    .clk(clknet_2_2_0_clk),
    .addr_in({net47,
    net46,
    net45,
    net44,
    net42,
    net41,
    net40,
    net39}),
    .rd_out({\dmem/inter_dmem2[31] ,
    \dmem/inter_dmem2[30] ,
    \dmem/inter_dmem2[29] ,
    \dmem/inter_dmem2[28] ,
    \dmem/inter_dmem2[27] ,
    \dmem/inter_dmem2[26] ,
    \dmem/inter_dmem2[25] ,
    \dmem/inter_dmem2[24] ,
    \dmem/inter_dmem2[23] ,
    \dmem/inter_dmem2[22] ,
    \dmem/inter_dmem2[21] ,
    \dmem/inter_dmem2[20] ,
    \dmem/inter_dmem2[19] ,
    \dmem/inter_dmem2[18] ,
    \dmem/inter_dmem2[17] ,
    \dmem/inter_dmem2[16] ,
    \dmem/inter_dmem2[15] ,
    \dmem/inter_dmem2[14] ,
    \dmem/inter_dmem2[13] ,
    \dmem/inter_dmem2[12] ,
    \dmem/inter_dmem2[11] ,
    \dmem/inter_dmem2[10] ,
    \dmem/inter_dmem2[9] ,
    \dmem/inter_dmem2[8] ,
    \dmem/inter_dmem2[7] ,
    \dmem/inter_dmem2[6] ,
    \dmem/inter_dmem2[5] ,
    \dmem/inter_dmem2[4] ,
    \dmem/inter_dmem2[3] ,
    \dmem/inter_dmem2[2] ,
    \dmem/inter_dmem2[1] ,
    \dmem/inter_dmem2[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net4,
    net165,
    net124,
    net121,
    net110,
    net99}));
 fakeram7_256x32 \dmem/dmem3  (.we_in(\dmem/we_mem[3] ),
    .ce_in(net56),
    .clk(clknet_2_2_0_clk),
    .addr_in({net56,
    net55,
    net53,
    net52,
    net51,
    net50,
    net49,
    net48}),
    .rd_out({\dmem/inter_dmem3[31] ,
    \dmem/inter_dmem3[30] ,
    \dmem/inter_dmem3[29] ,
    \dmem/inter_dmem3[28] ,
    \dmem/inter_dmem3[27] ,
    \dmem/inter_dmem3[26] ,
    \dmem/inter_dmem3[25] ,
    \dmem/inter_dmem3[24] ,
    \dmem/inter_dmem3[23] ,
    \dmem/inter_dmem3[22] ,
    \dmem/inter_dmem3[21] ,
    \dmem/inter_dmem3[20] ,
    \dmem/inter_dmem3[19] ,
    \dmem/inter_dmem3[18] ,
    \dmem/inter_dmem3[17] ,
    \dmem/inter_dmem3[16] ,
    \dmem/inter_dmem3[15] ,
    \dmem/inter_dmem3[14] ,
    \dmem/inter_dmem3[13] ,
    \dmem/inter_dmem3[12] ,
    \dmem/inter_dmem3[11] ,
    \dmem/inter_dmem3[10] ,
    \dmem/inter_dmem3[9] ,
    \dmem/inter_dmem3[8] ,
    \dmem/inter_dmem3[7] ,
    \dmem/inter_dmem3[6] ,
    \dmem/inter_dmem3[5] ,
    \dmem/inter_dmem3[4] ,
    \dmem/inter_dmem3[3] ,
    \dmem/inter_dmem3[2] ,
    \dmem/inter_dmem3[1] ,
    \dmem/inter_dmem3[0] }),
    .wd_in({net123,
    net122,
    net120,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net109,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net130,
    net129,
    net128,
    net127,
    net4,
    net166,
    net124,
    net121,
    net110,
    net99}));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[0]$_DFFE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .D(_01220_),
    .QN(_01066_),
    .RESETN(net131),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[10]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[10] ),
    .QN(_01093_),
    .RESETN(net132),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[11]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[11] ),
    .QN(_01096_),
    .RESETN(net133),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[12]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[12] ),
    .QN(_01099_),
    .RESETN(net134),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[13]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[13] ),
    .QN(_01102_),
    .RESETN(net135),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[14]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[14] ),
    .QN(_01105_),
    .RESETN(net136),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[15]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[15] ),
    .QN(_01108_),
    .RESETN(net137),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[16]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[16] ),
    .QN(_01111_),
    .RESETN(net138),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[17]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[17] ),
    .QN(_01114_),
    .RESETN(net139),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[18]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[18] ),
    .QN(_01117_),
    .RESETN(net140),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[19]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[19] ),
    .QN(_01120_),
    .RESETN(net141),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[1]$_DFFE_PP0P_  (.CLK(clknet_leaf_53_clk),
    .D(_01221_),
    .QN(_01068_),
    .RESETN(net142),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[20]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[20] ),
    .QN(_01123_),
    .RESETN(net143),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[21]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[21] ),
    .QN(_01126_),
    .RESETN(net144),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[22]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[22] ),
    .QN(_01129_),
    .RESETN(net145),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[23]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[23] ),
    .QN(_01132_),
    .RESETN(net146),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[24]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[24] ),
    .QN(_01135_),
    .RESETN(net147),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[25]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[25] ),
    .QN(_01138_),
    .RESETN(net148),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[26]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[26] ),
    .QN(_01141_),
    .RESETN(net149),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[27]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[27] ),
    .QN(_01144_),
    .RESETN(net150),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[28]$_DFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .D(\riscv.dp.ISRmux.d0[28] ),
    .QN(_01147_),
    .RESETN(net151),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[29]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[29] ),
    .QN(_01150_),
    .RESETN(net152),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[2]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[2] ),
    .QN(_09717_),
    .RESETN(net153),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[30]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[30] ),
    .QN(_01153_),
    .RESETN(net154),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[31]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[31] ),
    .QN(_01157_),
    .RESETN(net155),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[3]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[3] ),
    .QN(_09718_),
    .RESETN(net156),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[4]$_DFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .D(\riscv.dp.ISRmux.d0[4] ),
    .QN(_01075_),
    .RESETN(net157),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[5]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[5] ),
    .QN(_01078_),
    .RESETN(net158),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[6]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[6] ),
    .QN(_01081_),
    .RESETN(net159),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[7]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[7] ),
    .QN(_01084_),
    .RESETN(net160),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[8]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[8] ),
    .QN(_01087_),
    .RESETN(net161),
    .SETN(_01219_));
 DFFASRHQNx1_ASAP7_75t_R \riscv.dp.pcreg.q[9]$_DFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .D(\riscv.dp.ISRmux.d0[9] ),
    .QN(_01090_),
    .RESETN(net162),
    .SETN(_01219_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01222_),
    .QN(_00000_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01223_),
    .QN(_00732_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01224_),
    .QN(_00699_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01225_),
    .QN(_00666_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01226_),
    .QN(_00633_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01227_),
    .QN(_00600_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01228_),
    .QN(_00566_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01229_),
    .QN(_00533_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01230_),
    .QN(_00500_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01231_),
    .QN(_00467_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01232_),
    .QN(_00434_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01233_),
    .QN(_01032_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01234_),
    .QN(_00401_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01235_),
    .QN(_00368_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01236_),
    .QN(_00335_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01237_),
    .QN(_00301_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01238_),
    .QN(_00268_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01239_),
    .QN(_00235_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01240_),
    .QN(_00201_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01241_),
    .QN(_00168_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01242_),
    .QN(_00134_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01243_),
    .QN(_00101_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01244_),
    .QN(_00999_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01245_),
    .QN(_00067_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01246_),
    .QN(_00035_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01247_),
    .QN(_00966_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01248_),
    .QN(_00933_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01249_),
    .QN(_00899_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01250_),
    .QN(_00866_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01251_),
    .QN(_00832_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01252_),
    .QN(_00799_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01253_),
    .QN(_00765_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01254_),
    .QN(_00010_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01255_),
    .QN(_00742_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01256_),
    .QN(_00709_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][12]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01257_),
    .QN(_00676_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01258_),
    .QN(_00643_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][14]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01259_),
    .QN(_00610_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][15]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01260_),
    .QN(_00576_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][16]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01261_),
    .QN(_00543_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01262_),
    .QN(_00510_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01263_),
    .QN(_00477_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01264_),
    .QN(_00444_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01265_),
    .QN(_01042_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01266_),
    .QN(_00411_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][21]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01267_),
    .QN(_00378_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][22]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01268_),
    .QN(_00345_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01269_),
    .QN(_00311_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][24]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01270_),
    .QN(_00278_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01271_),
    .QN(_00245_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01272_),
    .QN(_00211_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01273_),
    .QN(_00178_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][28]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01274_),
    .QN(_00144_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01275_),
    .QN(_00111_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01276_),
    .QN(_01009_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01277_),
    .QN(_00077_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][31]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01278_),
    .QN(_00045_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01279_),
    .QN(_00976_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01280_),
    .QN(_00943_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01281_),
    .QN(_00909_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01282_),
    .QN(_00876_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01283_),
    .QN(_00842_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01284_),
    .QN(_00809_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01285_),
    .QN(_00775_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01286_),
    .QN(_00011_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01287_),
    .QN(_00743_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01288_),
    .QN(_00710_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01289_),
    .QN(_00677_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01290_),
    .QN(_00644_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01291_),
    .QN(_00611_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][15]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01292_),
    .QN(_00577_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][16]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01293_),
    .QN(_00544_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][17]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01294_),
    .QN(_00511_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][18]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01295_),
    .QN(_00478_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][19]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01296_),
    .QN(_00445_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01297_),
    .QN(_01043_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01298_),
    .QN(_00412_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][21]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01299_),
    .QN(_00379_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][22]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01300_),
    .QN(_00346_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01301_),
    .QN(_00312_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][24]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01302_),
    .QN(_00279_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01303_),
    .QN(_00246_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01304_),
    .QN(_00212_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01305_),
    .QN(_00179_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][28]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01306_),
    .QN(_00145_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01307_),
    .QN(_00112_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01308_),
    .QN(_01010_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01309_),
    .QN(_00078_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][31]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01310_),
    .QN(_00046_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01311_),
    .QN(_00977_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01312_),
    .QN(_00944_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01313_),
    .QN(_00910_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01314_),
    .QN(_00877_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01315_),
    .QN(_00843_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01316_),
    .QN(_00810_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01317_),
    .QN(_00776_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01318_),
    .QN(_00012_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01319_),
    .QN(_00744_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01320_),
    .QN(_00711_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01321_),
    .QN(_00678_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01322_),
    .QN(_00645_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01323_),
    .QN(_00612_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][15]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01324_),
    .QN(_00578_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][16]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01325_),
    .QN(_00545_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01326_),
    .QN(_00512_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01327_),
    .QN(_00479_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01328_),
    .QN(_00446_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01329_),
    .QN(_01044_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][20]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01330_),
    .QN(_00413_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][21]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01331_),
    .QN(_00380_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][22]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01332_),
    .QN(_00347_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][23]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01333_),
    .QN(_00313_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][24]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01334_),
    .QN(_00280_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01335_),
    .QN(_00247_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01336_),
    .QN(_00213_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01337_),
    .QN(_00180_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][28]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01338_),
    .QN(_00146_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][29]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01339_),
    .QN(_00113_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01340_),
    .QN(_01011_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01341_),
    .QN(_00079_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][31]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01342_),
    .QN(_00047_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01343_),
    .QN(_00978_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01344_),
    .QN(_00945_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01345_),
    .QN(_00911_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01346_),
    .QN(_00878_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01347_),
    .QN(_00844_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01348_),
    .QN(_00811_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01349_),
    .QN(_00777_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01350_),
    .QN(_00013_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01351_),
    .QN(_00745_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01352_),
    .QN(_00712_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01353_),
    .QN(_00679_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01354_),
    .QN(_00646_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][14]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01355_),
    .QN(_00613_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][15]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01356_),
    .QN(_00579_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][16]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01357_),
    .QN(_00546_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01358_),
    .QN(_00513_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01359_),
    .QN(_00480_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01360_),
    .QN(_00447_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01361_),
    .QN(_01045_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01362_),
    .QN(_00414_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][21]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01363_),
    .QN(_00381_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][22]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01364_),
    .QN(_00348_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01365_),
    .QN(_00314_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][24]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01366_),
    .QN(_00281_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01367_),
    .QN(_00248_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01368_),
    .QN(_00214_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01369_),
    .QN(_00181_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][28]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01370_),
    .QN(_00147_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][29]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01371_),
    .QN(_00114_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01372_),
    .QN(_01012_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][30]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01373_),
    .QN(_00080_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][31]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01374_),
    .QN(_00048_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01375_),
    .QN(_00979_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01376_),
    .QN(_00946_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01377_),
    .QN(_00912_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01378_),
    .QN(_00879_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01379_),
    .QN(_00845_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01380_),
    .QN(_00812_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01381_),
    .QN(_00778_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01382_),
    .QN(_00014_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01383_),
    .QN(_00746_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01384_),
    .QN(_00713_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][12]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01385_),
    .QN(_00680_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][13]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01386_),
    .QN(_00647_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][14]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01387_),
    .QN(_00614_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][15]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01388_),
    .QN(_00580_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][16]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01389_),
    .QN(_00547_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01390_),
    .QN(_00514_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01391_),
    .QN(_00481_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01392_),
    .QN(_00448_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01393_),
    .QN(_01046_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][20]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01394_),
    .QN(_00415_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][21]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01395_),
    .QN(_00382_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][22]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01396_),
    .QN(_00349_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01397_),
    .QN(_00315_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][24]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01398_),
    .QN(_00282_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01399_),
    .QN(_00249_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01400_),
    .QN(_00215_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01401_),
    .QN(_00182_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][28]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01402_),
    .QN(_00148_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][29]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01403_),
    .QN(_00115_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01404_),
    .QN(_01013_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01405_),
    .QN(_00081_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][31]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01406_),
    .QN(_00049_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01407_),
    .QN(_00980_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01408_),
    .QN(_00947_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01409_),
    .QN(_00913_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01410_),
    .QN(_00880_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01411_),
    .QN(_00846_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01412_),
    .QN(_00813_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01413_),
    .QN(_00779_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01414_),
    .QN(_00015_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01415_),
    .QN(_00747_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01416_),
    .QN(_00714_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][12]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01417_),
    .QN(_00681_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][13]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01418_),
    .QN(_00648_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][14]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01419_),
    .QN(_00615_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][15]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01420_),
    .QN(_00581_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][16]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01421_),
    .QN(_00548_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01422_),
    .QN(_00515_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01423_),
    .QN(_00482_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01424_),
    .QN(_00449_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01425_),
    .QN(_01047_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][20]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01426_),
    .QN(_00416_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][21]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01427_),
    .QN(_00383_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][22]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01428_),
    .QN(_00350_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][23]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01429_),
    .QN(_00316_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][24]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01430_),
    .QN(_00283_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01431_),
    .QN(_00250_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01432_),
    .QN(_00216_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01433_),
    .QN(_00183_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][28]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01434_),
    .QN(_00149_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][29]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01435_),
    .QN(_00116_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01436_),
    .QN(_01014_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][30]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01437_),
    .QN(_00082_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][31]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01438_),
    .QN(_00050_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01439_),
    .QN(_00981_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01440_),
    .QN(_00948_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01441_),
    .QN(_00914_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01442_),
    .QN(_00881_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01443_),
    .QN(_00847_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01444_),
    .QN(_00814_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01445_),
    .QN(_00780_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01446_),
    .QN(_00016_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01447_),
    .QN(_00748_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01448_),
    .QN(_00715_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][12]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01449_),
    .QN(_00682_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][13]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01450_),
    .QN(_00649_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01451_),
    .QN(_00616_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][15]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01452_),
    .QN(_00582_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][16]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01453_),
    .QN(_00549_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01454_),
    .QN(_00516_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01455_),
    .QN(_00483_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01456_),
    .QN(_00450_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01457_),
    .QN(_01048_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01458_),
    .QN(_00417_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][21]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01459_),
    .QN(_00384_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][22]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01460_),
    .QN(_00351_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01461_),
    .QN(_00317_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][24]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01462_),
    .QN(_00284_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01463_),
    .QN(_00251_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01464_),
    .QN(_00217_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01465_),
    .QN(_00184_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][28]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01466_),
    .QN(_00150_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][29]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01467_),
    .QN(_00117_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01468_),
    .QN(_01015_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01469_),
    .QN(_00083_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][31]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01470_),
    .QN(_00051_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01471_),
    .QN(_00982_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01472_),
    .QN(_00949_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01473_),
    .QN(_00915_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01474_),
    .QN(_00882_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01475_),
    .QN(_00848_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01476_),
    .QN(_00815_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01477_),
    .QN(_00781_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01478_),
    .QN(_00017_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01479_),
    .QN(_00749_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01480_),
    .QN(_00716_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][12]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01481_),
    .QN(_00683_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][13]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01482_),
    .QN(_00650_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01483_),
    .QN(_00617_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][15]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01484_),
    .QN(_00583_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][16]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01485_),
    .QN(_00550_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01486_),
    .QN(_00517_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01487_),
    .QN(_00484_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01488_),
    .QN(_00451_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01489_),
    .QN(_01049_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01490_),
    .QN(_00418_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][21]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01491_),
    .QN(_00385_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][22]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01492_),
    .QN(_00352_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01493_),
    .QN(_00318_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][24]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01494_),
    .QN(_00285_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][25]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01495_),
    .QN(_00252_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01496_),
    .QN(_00218_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01497_),
    .QN(_00185_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][28]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01498_),
    .QN(_00151_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01499_),
    .QN(_00118_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01500_),
    .QN(_01016_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01501_),
    .QN(_00084_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][31]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01502_),
    .QN(_00052_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01503_),
    .QN(_00983_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01504_),
    .QN(_00950_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01505_),
    .QN(_00916_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01506_),
    .QN(_00883_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01507_),
    .QN(_00849_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01508_),
    .QN(_00816_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01509_),
    .QN(_00782_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01510_),
    .QN(_00018_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01511_),
    .QN(_00750_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01512_),
    .QN(_00717_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01513_),
    .QN(_00684_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01514_),
    .QN(_00651_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01515_),
    .QN(_00618_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][15]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01516_),
    .QN(_00584_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][16]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01517_),
    .QN(_00551_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01518_),
    .QN(_00518_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01519_),
    .QN(_00485_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01520_),
    .QN(_00452_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01521_),
    .QN(_01050_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01522_),
    .QN(_00419_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][21]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01523_),
    .QN(_00386_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][22]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01524_),
    .QN(_00353_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][23]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01525_),
    .QN(_00319_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][24]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01526_),
    .QN(_00286_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01527_),
    .QN(_00253_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01528_),
    .QN(_00219_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01529_),
    .QN(_00186_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][28]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01530_),
    .QN(_00152_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][29]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01531_),
    .QN(_00119_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01532_),
    .QN(_01017_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01533_),
    .QN(_00085_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][31]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01534_),
    .QN(_00053_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01535_),
    .QN(_00984_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01536_),
    .QN(_00951_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01537_),
    .QN(_00917_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01538_),
    .QN(_00884_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01539_),
    .QN(_00850_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01540_),
    .QN(_00817_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01541_),
    .QN(_00783_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01542_),
    .QN(_00019_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01543_),
    .QN(_00751_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01544_),
    .QN(_00718_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01545_),
    .QN(_00685_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01546_),
    .QN(_00652_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .D(_01547_),
    .QN(_00619_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][15]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01548_),
    .QN(_00585_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][16]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01549_),
    .QN(_00552_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01550_),
    .QN(_00519_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][18]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01551_),
    .QN(_00486_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][19]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01552_),
    .QN(_00453_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01553_),
    .QN(_01051_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01554_),
    .QN(_00420_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][21]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01555_),
    .QN(_00387_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][22]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01556_),
    .QN(_00354_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01557_),
    .QN(_00320_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][24]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01558_),
    .QN(_00287_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01559_),
    .QN(_00254_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01560_),
    .QN(_00220_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01561_),
    .QN(_00187_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][28]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01562_),
    .QN(_00153_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01563_),
    .QN(_00120_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01564_),
    .QN(_01018_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][30]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01565_),
    .QN(_00086_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][31]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01566_),
    .QN(_00054_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01567_),
    .QN(_00985_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01568_),
    .QN(_00952_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01569_),
    .QN(_00918_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .D(_01570_),
    .QN(_00885_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .D(_01571_),
    .QN(_00851_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01572_),
    .QN(_00818_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01573_),
    .QN(_00784_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01574_),
    .QN(_00001_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01575_),
    .QN(_00733_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01576_),
    .QN(_00700_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01577_),
    .QN(_00667_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01578_),
    .QN(_00634_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01579_),
    .QN(_00601_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01580_),
    .QN(_00567_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .D(_01581_),
    .QN(_00534_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .D(_01582_),
    .QN(_00501_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01583_),
    .QN(_00468_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01584_),
    .QN(_00435_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01585_),
    .QN(_01033_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .D(_01586_),
    .QN(_00402_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01587_),
    .QN(_00369_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01588_),
    .QN(_00336_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01589_),
    .QN(_00302_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01590_),
    .QN(_00269_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01591_),
    .QN(_00236_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01592_),
    .QN(_00202_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01593_),
    .QN(_00169_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01594_),
    .QN(_00135_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01595_),
    .QN(_00102_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01596_),
    .QN(_01000_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .D(_01597_),
    .QN(_00068_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01598_),
    .QN(_00036_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01599_),
    .QN(_00967_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01600_),
    .QN(_00934_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .D(_01601_),
    .QN(_00900_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01602_),
    .QN(_00867_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .D(_01603_),
    .QN(_00833_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .D(_01604_),
    .QN(_00800_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .D(_01605_),
    .QN(_00766_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01606_),
    .QN(_00020_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01607_),
    .QN(_00752_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01608_),
    .QN(_00719_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][12]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01609_),
    .QN(_00686_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01610_),
    .QN(_00653_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01611_),
    .QN(_00620_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][15]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01612_),
    .QN(_00586_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][16]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01613_),
    .QN(_00553_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][17]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01614_),
    .QN(_00520_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][18]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01615_),
    .QN(_00487_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][19]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01616_),
    .QN(_00454_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01617_),
    .QN(_01052_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][20]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01618_),
    .QN(_00421_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][21]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01619_),
    .QN(_00388_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01620_),
    .QN(_00355_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][23]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01621_),
    .QN(_00321_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][24]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01622_),
    .QN(_00288_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][25]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01623_),
    .QN(_00255_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][26]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01624_),
    .QN(_00221_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][27]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01625_),
    .QN(_00188_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01626_),
    .QN(_00154_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][29]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01627_),
    .QN(_00121_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01628_),
    .QN(_01019_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][30]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01629_),
    .QN(_00087_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01630_),
    .QN(_00055_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01631_),
    .QN(_00986_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01632_),
    .QN(_00953_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01633_),
    .QN(_00919_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01634_),
    .QN(_00886_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01635_),
    .QN(_00852_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01636_),
    .QN(_00819_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01637_),
    .QN(_00785_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01638_),
    .QN(_00021_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01639_),
    .QN(_00753_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01640_),
    .QN(_00720_));
 DFFHQNx3_ASAP7_75t_R \riscv.dp.rf.rf[21][12]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01641_),
    .QN(_00687_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01642_),
    .QN(_00654_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01643_),
    .QN(_00621_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][15]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01644_),
    .QN(_00587_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][16]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01645_),
    .QN(_00554_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][17]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01646_),
    .QN(_00521_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][18]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01647_),
    .QN(_00488_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][19]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01648_),
    .QN(_00455_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01649_),
    .QN(_01053_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][20]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01650_),
    .QN(_00422_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][21]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01651_),
    .QN(_00389_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][22]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01652_),
    .QN(_00356_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01653_),
    .QN(_00322_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][24]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01654_),
    .QN(_00289_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][25]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01655_),
    .QN(_00256_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][26]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01656_),
    .QN(_00222_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01657_),
    .QN(_00189_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01658_),
    .QN(_00155_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][29]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01659_),
    .QN(_00122_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01660_),
    .QN(_01020_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][30]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01661_),
    .QN(_00088_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01662_),
    .QN(_00056_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01663_),
    .QN(_00987_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01664_),
    .QN(_00954_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01665_),
    .QN(_00920_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01666_),
    .QN(_00887_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01667_),
    .QN(_00853_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01668_),
    .QN(_00820_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01669_),
    .QN(_00786_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01670_),
    .QN(_00022_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01671_),
    .QN(_00754_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01672_),
    .QN(_00721_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01673_),
    .QN(_00688_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01674_),
    .QN(_00655_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01675_),
    .QN(_00622_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][15]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01676_),
    .QN(_00588_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][16]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01677_),
    .QN(_00555_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01678_),
    .QN(_00522_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][18]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01679_),
    .QN(_00489_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][19]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01680_),
    .QN(_00456_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01681_),
    .QN(_01054_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][20]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01682_),
    .QN(_00423_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01683_),
    .QN(_00390_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01684_),
    .QN(_00357_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01685_),
    .QN(_00323_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][24]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01686_),
    .QN(_00290_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][25]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01687_),
    .QN(_00257_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][26]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01688_),
    .QN(_00223_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01689_),
    .QN(_00190_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][28]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01690_),
    .QN(_00156_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][29]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01691_),
    .QN(_00123_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01692_),
    .QN(_01021_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01693_),
    .QN(_00089_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01694_),
    .QN(_00057_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01695_),
    .QN(_00988_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01696_),
    .QN(_00955_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01697_),
    .QN(_00921_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .D(_01698_),
    .QN(_00888_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01699_),
    .QN(_00854_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01700_),
    .QN(_00821_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01701_),
    .QN(_00787_));
 DFFHQNx3_ASAP7_75t_R \riscv.dp.rf.rf[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01702_),
    .QN(_00023_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01703_),
    .QN(_00755_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .D(_01704_),
    .QN(_00722_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][12]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01705_),
    .QN(_00689_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01706_),
    .QN(_00656_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01707_),
    .QN(_00623_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][15]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01708_),
    .QN(_00589_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][16]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01709_),
    .QN(_00556_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01710_),
    .QN(_00523_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][18]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01711_),
    .QN(_00490_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][19]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01712_),
    .QN(_00457_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01713_),
    .QN(_01055_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][20]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01714_),
    .QN(_00424_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01715_),
    .QN(_00391_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][22]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01716_),
    .QN(_00358_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][23]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01717_),
    .QN(_00324_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][24]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01718_),
    .QN(_00291_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][25]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01719_),
    .QN(_00258_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][26]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01720_),
    .QN(_00224_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01721_),
    .QN(_00191_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][28]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01722_),
    .QN(_00157_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][29]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .D(_01723_),
    .QN(_00124_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01724_),
    .QN(_01022_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01725_),
    .QN(_00090_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01726_),
    .QN(_00058_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01727_),
    .QN(_00989_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01728_),
    .QN(_00956_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01729_),
    .QN(_00922_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .D(_01730_),
    .QN(_00889_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01731_),
    .QN(_00855_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01732_),
    .QN(_00822_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01733_),
    .QN(_00788_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01734_),
    .QN(_00024_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01735_),
    .QN(_00756_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01736_),
    .QN(_00723_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01737_),
    .QN(_00690_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01738_),
    .QN(_00657_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][14]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01739_),
    .QN(_00624_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][15]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01740_),
    .QN(_00590_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][16]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .D(_01741_),
    .QN(_00557_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01742_),
    .QN(_00524_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][18]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01743_),
    .QN(_00491_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][19]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01744_),
    .QN(_00458_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01745_),
    .QN(_01056_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][20]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01746_),
    .QN(_00425_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][21]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01747_),
    .QN(_00392_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01748_),
    .QN(_00359_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01749_),
    .QN(_00325_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01750_),
    .QN(_00292_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01751_),
    .QN(_00259_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][26]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01752_),
    .QN(_00225_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][27]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01753_),
    .QN(_00192_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][28]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01754_),
    .QN(_00158_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][29]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01755_),
    .QN(_00125_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01756_),
    .QN(_01023_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01757_),
    .QN(_00091_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01758_),
    .QN(_00059_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01759_),
    .QN(_00990_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01760_),
    .QN(_00957_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01761_),
    .QN(_00923_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01762_),
    .QN(_00890_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01763_),
    .QN(_00856_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01764_),
    .QN(_00823_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01765_),
    .QN(_00789_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01766_),
    .QN(_00025_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01767_),
    .QN(_00757_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01768_),
    .QN(_00724_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01769_),
    .QN(_00691_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01770_),
    .QN(_00658_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][14]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01771_),
    .QN(_00625_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][15]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01772_),
    .QN(_00591_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][16]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01773_),
    .QN(_00558_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01774_),
    .QN(_00525_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][18]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01775_),
    .QN(_00492_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][19]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .D(_01776_),
    .QN(_00459_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01777_),
    .QN(_01057_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][20]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01778_),
    .QN(_00426_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01779_),
    .QN(_00393_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01780_),
    .QN(_00360_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01781_),
    .QN(_00326_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01782_),
    .QN(_00293_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01783_),
    .QN(_00260_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][26]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01784_),
    .QN(_00226_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][27]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01785_),
    .QN(_00193_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][28]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01786_),
    .QN(_00159_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01787_),
    .QN(_00126_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01788_),
    .QN(_01024_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01789_),
    .QN(_00092_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01790_),
    .QN(_00060_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01791_),
    .QN(_00991_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01792_),
    .QN(_00958_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01793_),
    .QN(_00924_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01794_),
    .QN(_00891_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01795_),
    .QN(_00857_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01796_),
    .QN(_00824_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01797_),
    .QN(_00790_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01798_),
    .QN(_00026_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01799_),
    .QN(_00758_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01800_),
    .QN(_00725_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01801_),
    .QN(_00692_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01802_),
    .QN(_00659_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][14]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01803_),
    .QN(_00626_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][15]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01804_),
    .QN(_00592_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][16]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01805_),
    .QN(_00559_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][17]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01806_),
    .QN(_00526_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][18]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01807_),
    .QN(_00493_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][19]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01808_),
    .QN(_00460_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01809_),
    .QN(_01058_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][20]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01810_),
    .QN(_00427_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01811_),
    .QN(_00394_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01812_),
    .QN(_00361_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01813_),
    .QN(_00327_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01814_),
    .QN(_00294_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01815_),
    .QN(_00261_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][26]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01816_),
    .QN(_00227_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][27]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01817_),
    .QN(_00194_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][28]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01818_),
    .QN(_00160_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][29]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01819_),
    .QN(_00127_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01820_),
    .QN(_01025_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01821_),
    .QN(_00093_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01822_),
    .QN(_00061_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01823_),
    .QN(_00992_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01824_),
    .QN(_00959_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01825_),
    .QN(_00925_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01826_),
    .QN(_00892_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01827_),
    .QN(_00858_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01828_),
    .QN(_00825_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01829_),
    .QN(_00791_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01830_),
    .QN(_00027_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01831_),
    .QN(_00759_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01832_),
    .QN(_00726_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01833_),
    .QN(_00693_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01834_),
    .QN(_00660_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][14]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01835_),
    .QN(_00627_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][15]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01836_),
    .QN(_00593_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][16]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .D(_01837_),
    .QN(_00560_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][17]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01838_),
    .QN(_00527_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01839_),
    .QN(_00494_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][19]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01840_),
    .QN(_00461_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01841_),
    .QN(_01059_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][20]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01842_),
    .QN(_00428_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][21]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01843_),
    .QN(_00395_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01844_),
    .QN(_00362_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][23]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01845_),
    .QN(_00328_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01846_),
    .QN(_00295_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01847_),
    .QN(_00262_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][26]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01848_),
    .QN(_00228_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][27]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01849_),
    .QN(_00195_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][28]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01850_),
    .QN(_00161_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01851_),
    .QN(_00128_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01852_),
    .QN(_01026_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01853_),
    .QN(_00094_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01854_),
    .QN(_00062_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01855_),
    .QN(_00993_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01856_),
    .QN(_00960_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01857_),
    .QN(_00926_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01858_),
    .QN(_00893_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01859_),
    .QN(_00859_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01860_),
    .QN(_00826_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01861_),
    .QN(_00792_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01862_),
    .QN(_00028_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01863_),
    .QN(_00760_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01864_),
    .QN(_00727_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][12]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01865_),
    .QN(_00694_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01866_),
    .QN(_00661_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][14]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01867_),
    .QN(_00628_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][15]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01868_),
    .QN(_00594_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][16]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01869_),
    .QN(_00561_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01870_),
    .QN(_00528_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01871_),
    .QN(_00495_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][19]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01872_),
    .QN(_00462_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01873_),
    .QN(_01060_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][20]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01874_),
    .QN(_00429_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][21]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01875_),
    .QN(_00396_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01876_),
    .QN(_00363_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01877_),
    .QN(_00329_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01878_),
    .QN(_00296_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01879_),
    .QN(_00263_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][26]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .D(_01880_),
    .QN(_00229_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01881_),
    .QN(_00196_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_01882_),
    .QN(_00162_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01883_),
    .QN(_00129_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01884_),
    .QN(_01027_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01885_),
    .QN(_00095_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01886_),
    .QN(_00063_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01887_),
    .QN(_00994_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01888_),
    .QN(_00961_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01889_),
    .QN(_00927_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .D(_01890_),
    .QN(_00894_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .D(_01891_),
    .QN(_00860_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01892_),
    .QN(_00827_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .D(_01893_),
    .QN(_00793_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01894_),
    .QN(_00029_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01895_),
    .QN(_00761_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01896_),
    .QN(_00728_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_01897_),
    .QN(_00695_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01898_),
    .QN(_00662_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][14]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01899_),
    .QN(_00629_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][15]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .D(_01900_),
    .QN(_00595_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][16]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01901_),
    .QN(_00562_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01902_),
    .QN(_00529_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01903_),
    .QN(_00496_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][19]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01904_),
    .QN(_00463_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01905_),
    .QN(_01061_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][20]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01906_),
    .QN(_00430_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01907_),
    .QN(_00397_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01908_),
    .QN(_00364_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][23]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01909_),
    .QN(_00330_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][24]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01910_),
    .QN(_00297_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01911_),
    .QN(_00264_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][26]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01912_),
    .QN(_00230_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][27]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01913_),
    .QN(_00197_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_01914_),
    .QN(_00163_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][29]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01915_),
    .QN(_00130_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01916_),
    .QN(_01028_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01917_),
    .QN(_00096_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01918_),
    .QN(_00064_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01919_),
    .QN(_00995_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01920_),
    .QN(_00962_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01921_),
    .QN(_00928_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01922_),
    .QN(_00895_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01923_),
    .QN(_00861_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01924_),
    .QN(_00828_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_01925_),
    .QN(_00794_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01926_),
    .QN(_00002_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01927_),
    .QN(_00734_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01928_),
    .QN(_00701_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01929_),
    .QN(_00668_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_01930_),
    .QN(_00635_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01931_),
    .QN(_00602_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01932_),
    .QN(_00568_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01933_),
    .QN(_00535_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01934_),
    .QN(_00502_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01935_),
    .QN(_00469_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_01936_),
    .QN(_00436_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01937_),
    .QN(_01034_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01938_),
    .QN(_00403_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01939_),
    .QN(_00370_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01940_),
    .QN(_00337_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01941_),
    .QN(_00303_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01942_),
    .QN(_00270_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01943_),
    .QN(_00237_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01944_),
    .QN(_00203_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01945_),
    .QN(_00170_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_01946_),
    .QN(_00136_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01947_),
    .QN(_00103_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01948_),
    .QN(_01001_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01949_),
    .QN(_00069_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01950_),
    .QN(_00037_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01951_),
    .QN(_00968_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01952_),
    .QN(_00935_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01953_),
    .QN(_00901_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01954_),
    .QN(_00868_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01955_),
    .QN(_00834_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01956_),
    .QN(_00801_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01957_),
    .QN(_00767_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01958_),
    .QN(_00030_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01959_),
    .QN(_00762_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01960_),
    .QN(_00729_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][12]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01961_),
    .QN(_00696_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][13]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01962_),
    .QN(_00663_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][14]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01963_),
    .QN(_00630_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][15]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01964_),
    .QN(_00596_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01965_),
    .QN(_00563_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01966_),
    .QN(_00530_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01967_),
    .QN(_00497_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][19]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01968_),
    .QN(_00464_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01969_),
    .QN(_01062_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][20]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01970_),
    .QN(_00431_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][21]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01971_),
    .QN(_00398_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01972_),
    .QN(_00365_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01973_),
    .QN(_00331_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01974_),
    .QN(_00298_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01975_),
    .QN(_00265_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][26]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01976_),
    .QN(_00231_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01977_),
    .QN(_00198_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][28]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01978_),
    .QN(_00164_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01979_),
    .QN(_00131_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_01980_),
    .QN(_01029_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][30]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01981_),
    .QN(_00097_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01982_),
    .QN(_00065_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01983_),
    .QN(_00996_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01984_),
    .QN(_00963_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01985_),
    .QN(_00929_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01986_),
    .QN(_00896_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01987_),
    .QN(_00862_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01988_),
    .QN(_00829_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01989_),
    .QN(_00795_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01990_),
    .QN(_00031_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01991_),
    .QN(_00763_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_01992_),
    .QN(_00730_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_01993_),
    .QN(_00697_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][13]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_01994_),
    .QN(_00664_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][14]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01995_),
    .QN(_00631_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][15]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_01996_),
    .QN(_00597_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01997_),
    .QN(_00564_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_01998_),
    .QN(_00531_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_01999_),
    .QN(_00498_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][19]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_02000_),
    .QN(_00465_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02001_),
    .QN(_01063_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][20]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_02002_),
    .QN(_00432_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][21]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02003_),
    .QN(_00399_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02004_),
    .QN(_00366_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02005_),
    .QN(_00332_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02006_),
    .QN(_00299_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02007_),
    .QN(_00266_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][26]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02008_),
    .QN(_00232_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][27]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02009_),
    .QN(_00199_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][28]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_02010_),
    .QN(_00165_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][29]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02011_),
    .QN(_00132_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_02012_),
    .QN(_01030_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][30]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02013_),
    .QN(_00098_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02014_),
    .QN(_00066_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02015_),
    .QN(_00997_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02016_),
    .QN(_00964_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02017_),
    .QN(_00930_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02018_),
    .QN(_00897_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02019_),
    .QN(_00863_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02020_),
    .QN(_00830_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02021_),
    .QN(_00796_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02022_),
    .QN(_00003_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02023_),
    .QN(_00735_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02024_),
    .QN(_00702_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_02025_),
    .QN(_00669_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02026_),
    .QN(_00636_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02027_),
    .QN(_00603_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02028_),
    .QN(_00569_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02029_),
    .QN(_00536_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02030_),
    .QN(_00503_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02031_),
    .QN(_00470_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_02032_),
    .QN(_00437_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_02033_),
    .QN(_01035_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02034_),
    .QN(_00404_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02035_),
    .QN(_00371_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02036_),
    .QN(_00338_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02037_),
    .QN(_00304_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02038_),
    .QN(_00271_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02039_),
    .QN(_00238_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02040_),
    .QN(_00204_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02041_),
    .QN(_00171_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02042_),
    .QN(_00137_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02043_),
    .QN(_00104_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_02044_),
    .QN(_01002_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02045_),
    .QN(_00070_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02046_),
    .QN(_00038_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02047_),
    .QN(_00969_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02048_),
    .QN(_00936_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_02049_),
    .QN(_00902_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02050_),
    .QN(_00869_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02051_),
    .QN(_00835_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02052_),
    .QN(_00802_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02053_),
    .QN(_00768_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02054_),
    .QN(_00004_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02055_),
    .QN(_00736_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02056_),
    .QN(_00703_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02057_),
    .QN(_00670_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02058_),
    .QN(_00637_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02059_),
    .QN(_00604_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02060_),
    .QN(_00570_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02061_),
    .QN(_00537_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02062_),
    .QN(_00504_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02063_),
    .QN(_00471_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02064_),
    .QN(_00438_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02065_),
    .QN(_01036_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02066_),
    .QN(_00405_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02067_),
    .QN(_00372_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02068_),
    .QN(_00339_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02069_),
    .QN(_00305_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02070_),
    .QN(_00272_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02071_),
    .QN(_00239_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02072_),
    .QN(_00205_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02073_),
    .QN(_00172_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02074_),
    .QN(_00138_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02075_),
    .QN(_00105_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_02076_),
    .QN(_01003_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_02077_),
    .QN(_00071_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02078_),
    .QN(_00039_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02079_),
    .QN(_00970_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02080_),
    .QN(_00937_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02081_),
    .QN(_00903_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02082_),
    .QN(_00870_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02083_),
    .QN(_00836_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02084_),
    .QN(_00803_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02085_),
    .QN(_00769_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02086_),
    .QN(_00005_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02087_),
    .QN(_00737_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02088_),
    .QN(_00704_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02089_),
    .QN(_00671_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02090_),
    .QN(_00638_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02091_),
    .QN(_00605_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02092_),
    .QN(_00571_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02093_),
    .QN(_00538_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_02094_),
    .QN(_00505_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02095_),
    .QN(_00472_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_02096_),
    .QN(_00439_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02097_),
    .QN(_01037_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02098_),
    .QN(_00406_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02099_),
    .QN(_00373_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02100_),
    .QN(_00340_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02101_),
    .QN(_00306_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02102_),
    .QN(_00273_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02103_),
    .QN(_00240_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02104_),
    .QN(_00206_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02105_),
    .QN(_00173_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02106_),
    .QN(_00139_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02107_),
    .QN(_00106_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02108_),
    .QN(_01004_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02109_),
    .QN(_00072_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02110_),
    .QN(_00040_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02111_),
    .QN(_00971_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02112_),
    .QN(_00938_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02113_),
    .QN(_00904_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02114_),
    .QN(_00871_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02115_),
    .QN(_00837_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02116_),
    .QN(_00804_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02117_),
    .QN(_00770_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_02118_),
    .QN(_00006_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02119_),
    .QN(_00738_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02120_),
    .QN(_00705_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02121_),
    .QN(_00672_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_02122_),
    .QN(_00639_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02123_),
    .QN(_00606_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02124_),
    .QN(_00572_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02125_),
    .QN(_00539_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02126_),
    .QN(_00506_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02127_),
    .QN(_00473_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_02128_),
    .QN(_00440_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02129_),
    .QN(_01038_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02130_),
    .QN(_00407_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02131_),
    .QN(_00374_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02132_),
    .QN(_00341_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02133_),
    .QN(_00307_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02134_),
    .QN(_00274_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02135_),
    .QN(_00241_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02136_),
    .QN(_00207_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02137_),
    .QN(_00174_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02138_),
    .QN(_00140_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02139_),
    .QN(_00107_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_02140_),
    .QN(_01005_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02141_),
    .QN(_00073_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02142_),
    .QN(_00041_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02143_),
    .QN(_00972_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02144_),
    .QN(_00939_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02145_),
    .QN(_00905_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02146_),
    .QN(_00872_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02147_),
    .QN(_00838_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02148_),
    .QN(_00805_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02149_),
    .QN(_00771_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_02150_),
    .QN(_00007_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02151_),
    .QN(_00739_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02152_),
    .QN(_00706_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_02153_),
    .QN(_00673_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_02154_),
    .QN(_00640_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02155_),
    .QN(_00607_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02156_),
    .QN(_00573_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02157_),
    .QN(_00540_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02158_),
    .QN(_00507_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02159_),
    .QN(_00474_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_02160_),
    .QN(_00441_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02161_),
    .QN(_01039_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02162_),
    .QN(_00408_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02163_),
    .QN(_00375_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02164_),
    .QN(_00342_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02165_),
    .QN(_00308_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02166_),
    .QN(_00275_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02167_),
    .QN(_00242_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02168_),
    .QN(_00208_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02169_),
    .QN(_00175_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_02170_),
    .QN(_00141_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02171_),
    .QN(_00108_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .D(_02172_),
    .QN(_01006_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02173_),
    .QN(_00074_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02174_),
    .QN(_00042_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02175_),
    .QN(_00973_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02176_),
    .QN(_00940_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02177_),
    .QN(_00906_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02178_),
    .QN(_00873_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02179_),
    .QN(_00839_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_02180_),
    .QN(_00806_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02181_),
    .QN(_00772_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02182_),
    .QN(_00008_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02183_),
    .QN(_00740_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02184_),
    .QN(_00707_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][12]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02185_),
    .QN(_00674_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][13]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02186_),
    .QN(_00641_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][14]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02187_),
    .QN(_00608_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][15]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_02188_),
    .QN(_00574_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02189_),
    .QN(_00541_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .D(_02190_),
    .QN(_00508_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_02191_),
    .QN(_00475_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][19]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_02192_),
    .QN(_00442_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02193_),
    .QN(_01040_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][20]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02194_),
    .QN(_00409_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][21]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02195_),
    .QN(_00376_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][22]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02196_),
    .QN(_00343_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02197_),
    .QN(_00309_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][24]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02198_),
    .QN(_00276_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][25]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_02199_),
    .QN(_00243_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][26]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02200_),
    .QN(_00209_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][27]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02201_),
    .QN(_00176_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][28]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02202_),
    .QN(_00142_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][29]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_02203_),
    .QN(_00109_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .D(_02204_),
    .QN(_01007_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][30]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02205_),
    .QN(_00075_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][31]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .D(_02206_),
    .QN(_00043_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02207_),
    .QN(_00974_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02208_),
    .QN(_00941_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_02209_),
    .QN(_00907_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02210_),
    .QN(_00874_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02211_),
    .QN(_00840_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02212_),
    .QN(_00807_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .D(_02213_),
    .QN(_00773_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02214_),
    .QN(_00009_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02215_),
    .QN(_00741_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02216_),
    .QN(_00708_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][12]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02217_),
    .QN(_00675_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02218_),
    .QN(_00642_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][14]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02219_),
    .QN(_00609_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][15]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .D(_02220_),
    .QN(_00575_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02221_),
    .QN(_00542_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][17]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_02222_),
    .QN(_00509_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][18]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .D(_02223_),
    .QN(_00476_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][19]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .D(_02224_),
    .QN(_00443_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02225_),
    .QN(_01041_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][20]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_02226_),
    .QN(_00410_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][21]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_02227_),
    .QN(_00377_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][22]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_02228_),
    .QN(_00344_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][23]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02229_),
    .QN(_00310_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][24]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_02230_),
    .QN(_00277_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][25]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_02231_),
    .QN(_00244_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][26]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_02232_),
    .QN(_00210_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][27]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_02233_),
    .QN(_00177_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][28]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02234_),
    .QN(_00143_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][29]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_02235_),
    .QN(_00110_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02236_),
    .QN(_01008_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_02237_),
    .QN(_00076_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][31]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_02238_),
    .QN(_00044_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02239_),
    .QN(_00975_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_02240_),
    .QN(_00942_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02241_),
    .QN(_00908_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02242_),
    .QN(_00875_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_02243_),
    .QN(_00841_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .D(_02244_),
    .QN(_00808_));
 DFFHQNx2_ASAP7_75t_R \riscv.dp.rf.rf[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_02245_),
    .QN(_00774_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Left_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Left_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Left_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Left_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Left_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Left_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Left_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Left_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Left_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Left_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Left_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Left_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Left_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Left_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Left_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Right_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Right_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Right_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Right_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Right_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Right_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Right_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Right_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_5_Right_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_5_Right_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_5_Right_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_5_Right_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_5_Right_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_5_Right_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_5_Right_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_5_Right_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_5_Right_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_5_Right_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_5_Right_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_5_Right_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_5_Right_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_5_Right_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_5_Right_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_5_Right_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_5_Right_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_5_Right_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_5_Right_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_5_Right_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_5_Right_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_5_Right_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_5_Right_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_5_Right_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_5_Right_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_5_Right_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_5_Right_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_5_Right_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_5_Right_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_5_Right_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_5_Right_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_5_Right_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_5_Right_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_5_Right_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_5_Right_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_5_Right_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_5_Right_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_5_Right_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_5_Right_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_5_Right_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_5_Right_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_5_Right_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_5_Right_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_5_Right_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_5_Right_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_5_Right_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_5_Right_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_5_Right_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_5_Right_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_5_Right_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_5_Right_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_5_Right_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_5_Right_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_5_Right_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_5_Right_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_5_Right_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_5_Right_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_5_Right_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_5_Right_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_5_Right_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_5_Right_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_5_Right_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_5_Right_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_5_Right_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_5_Right_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_5_Right_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_5_Right_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_5_Right_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_5_Right_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_5_Right_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_5_Right_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_5_Right_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_5_Right_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_5_Right_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_5_Right_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_5_Right_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_5_Right_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_5_Right_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_5_Right_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_5_Right_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_5_Right_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_5_Right_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_5_Right_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_5_Right_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_5_Right_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_5_Right_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_5_Right_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_5_Right_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_5_Right_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_5_Right_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_5_Right_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_5_Right_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_5_Right_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_5_Right_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_5_Right_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_5_Right_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_5_Right_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_5_Right_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_5_Right_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_5_Right_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_5_Right_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_5_Right_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_5_Right_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_5_Right_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_5_Right_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_5_Right_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_5_Right_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_5_Right_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_5_Right_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_5_Right_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_5_Right_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_5_Right_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_5_Right_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_5_Right_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_5_Right_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_5_Right_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_5_Right_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_5_Right_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_5_Right_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_5_Right_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_5_Right_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_5_Right_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_5_Right_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_5_Right_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_5_Right_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_5_Right_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_5_Right_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_5_Right_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_5_Right_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_5_Right_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_5_Right_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_5_Right_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_5_Right_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_5_Right_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_5_Right_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_5_Right_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_5_Right_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_5_Right_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_5_Right_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_5_Right_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_5_Right_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_5_Right_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_5_Right_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_5_Right_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_5_Right_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_5_Right_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_5_Right_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_5_Right_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_5_Right_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_5_Right_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_5_Right_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_5_Right_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_5_Right_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_5_Right_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_5_Right_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_5_Right_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_5_Right_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_5_Right_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_5_Right_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_5_Right_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_5_Right_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_5_Right_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_5_Right_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_5_Right_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_5_Right_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_5_Right_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_5_Right_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_5_Right_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_5_Right_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_5_Right_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_5_Right_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_5_Left_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_5_Left_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_5_Left_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_5_Left_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_5_Left_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_5_Left_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_5_Left_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_5_Left_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_5_Left_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_5_Left_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_5_Left_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_5_Left_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_5_Left_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_5_Left_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_5_Left_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_5_Left_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_5_Left_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_5_Left_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_5_Left_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_5_Left_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_5_Left_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_5_Left_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_5_Left_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_5_Left_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_5_Left_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_5_Left_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_5_Left_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_5_Left_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_5_Left_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_5_Left_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_5_Left_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_5_Left_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_5_Left_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_5_Left_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_5_Left_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_5_Left_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_5_Left_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_5_Left_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_5_Left_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_5_Left_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_5_Left_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_5_Left_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_5_Left_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_5_Left_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_5_Left_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_5_Left_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_5_Left_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_5_Left_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_5_Left_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_5_Left_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_5_Left_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_5_Left_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_5_Left_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_5_Left_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_5_Left_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_5_Left_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_5_Left_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_5_Left_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_5_Left_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_5_Left_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_5_Left_479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_5_Left_480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_5_Left_481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_5_Left_482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_5_Left_483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_5_Left_484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_5_Left_485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_5_Left_486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_5_Left_487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_5_Left_488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_5_Left_489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_5_Left_490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_5_Left_491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_5_Left_492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_5_Left_493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_5_Left_494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_5_Left_495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_5_Left_496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_5_Left_497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_5_Left_498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_5_Left_499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_5_Left_500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_5_Left_501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_5_Left_502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_5_Left_503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_5_Left_504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_5_Left_505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_5_Left_506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_5_Left_507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_5_Left_508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_5_Left_509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_5_Left_510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_5_Left_511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_5_Left_512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_5_Left_513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_5_Left_514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_5_Left_515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_5_Left_516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_5_Left_517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_5_Left_518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_5_Left_519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_5_Left_520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_5_Left_521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_5_Left_522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_5_Left_523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_5_Left_524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_5_Left_525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_5_Left_526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_5_Left_527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_5_Left_528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_5_Left_529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_5_Left_530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_5_Left_531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_5_Left_532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_5_Left_533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_5_Left_534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_5_Left_535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_5_Left_536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_5_Left_537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_5_Left_538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_5_Left_539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_5_Left_540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_5_Left_541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_5_Left_542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_5_Left_543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_5_Left_544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_5_Left_545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_5_Left_546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_5_Left_547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_5_Left_548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_5_Left_549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_5_Left_550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_5_Left_551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_5_Left_552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_5_Left_553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_5_Left_554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_5_Left_555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_5_Left_556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_5_Left_557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_5_Left_558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_5_Left_559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_5_Left_560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_5_Left_561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_5_Left_562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_5_Left_563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_5_Left_564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_5_Left_565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_5_Left_566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_5_Left_567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_5_Left_568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_5_Left_569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_5_Left_570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_5_Left_571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_5_Left_572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_5_Left_573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_5_Left_574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_5_Left_575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_5_Left_576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_5_Left_577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_5_Left_578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_5_Left_579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_5_Left_580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_5_Left_581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_5_Left_582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_5_Left_583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_5_Left_584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_5_Left_585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_5_Left_586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_5_Left_587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_5_Left_588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_5_Left_589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_15_606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_17_608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_19_610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_21_612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_23_614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_25_616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_27_618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_29_620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_31_622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_33_624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_35_626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_37_628 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_629 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_39_630 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_631 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_41_632 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_633 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_43_634 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_635 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_45_636 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_637 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_47_638 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_639 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_49_640 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_641 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_51_642 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_643 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_53_644 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_645 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_55_646 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_647 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_57_648 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_649 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_59_650 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_651 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_61_652 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_653 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_63_654 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_655 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_65_656 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_657 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_67_658 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_659 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_69_660 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_661 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_71_662 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_663 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_73_664 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_665 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_75_666 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_667 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_77_668 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_669 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_79_670 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_671 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_81_672 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_673 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_83_674 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_675 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_85_676 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_677 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_87_678 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_679 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_89_680 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_681 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_91_682 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_683 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_684 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_685 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_95_686 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_687 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_97_688 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_689 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_99_690 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_691 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_101_692 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_693 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_103_694 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_695 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_105_696 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_697 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_107_698 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_699 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_109_700 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_701 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_111_702 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_703 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_113_704 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_705 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_115_706 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_707 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_117_708 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_709 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_119_710 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_711 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_121_712 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_713 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_123_714 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_123_715 ();
 BUFx12f_ASAP7_75t_R max_cap3 (.A(net4),
    .Y(net126));
 BUFx16f_ASAP7_75t_R wire4 (.A(net3),
    .Y(net4));
 BUFx2_ASAP7_75t_R input1 (.A(instr[0]),
    .Y(net1));
 BUFx4f_ASAP7_75t_R input2 (.A(instr[10]),
    .Y(net2));
 BUFx4f_ASAP7_75t_R input3 (.A(instr[11]),
    .Y(net5));
 BUFx3_ASAP7_75t_R input4 (.A(instr[14]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input5 (.A(instr[16]),
    .Y(net7));
 BUFx2_ASAP7_75t_R input6 (.A(instr[17]),
    .Y(net8));
 BUFx10_ASAP7_75t_R input7 (.A(instr[18]),
    .Y(net9));
 BUFx2_ASAP7_75t_R input8 (.A(instr[19]),
    .Y(net10));
 BUFx2_ASAP7_75t_R input9 (.A(instr[1]),
    .Y(net11));
 BUFx6f_ASAP7_75t_R input10 (.A(instr[21]),
    .Y(net12));
 BUFx6f_ASAP7_75t_R input11 (.A(instr[22]),
    .Y(net13));
 BUFx4f_ASAP7_75t_R input12 (.A(instr[23]),
    .Y(net14));
 BUFx4f_ASAP7_75t_R input13 (.A(instr[24]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input14 (.A(instr[25]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input15 (.A(instr[26]),
    .Y(net17));
 BUFx2_ASAP7_75t_R input16 (.A(instr[27]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input17 (.A(instr[28]),
    .Y(net19));
 BUFx2_ASAP7_75t_R input18 (.A(instr[29]),
    .Y(net20));
 BUFx3_ASAP7_75t_R input19 (.A(instr[2]),
    .Y(net21));
 BUFx4f_ASAP7_75t_R input20 (.A(instr[30]),
    .Y(net22));
 BUFx2_ASAP7_75t_R input21 (.A(instr[31]),
    .Y(net23));
 BUFx12f_ASAP7_75t_R input22 (.A(instr[3]),
    .Y(net24));
 BUFx3_ASAP7_75t_R input23 (.A(instr[4]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input24 (.A(instr[5]),
    .Y(net26));
 BUFx4f_ASAP7_75t_R input25 (.A(instr[6]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input26 (.A(instr[7]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input27 (.A(instr[8]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input28 (.A(instr[9]),
    .Y(net30));
 BUFx6f_ASAP7_75t_R input29 (.A(reset),
    .Y(net31));
 BUFx2_ASAP7_75t_R output30 (.A(net32),
    .Y(dataadr[0]));
 BUFx2_ASAP7_75t_R output31 (.A(net33),
    .Y(dataadr[10]));
 BUFx2_ASAP7_75t_R output32 (.A(net34),
    .Y(dataadr[11]));
 BUFx2_ASAP7_75t_R output33 (.A(net35),
    .Y(dataadr[12]));
 BUFx2_ASAP7_75t_R output34 (.A(net36),
    .Y(dataadr[13]));
 BUFx2_ASAP7_75t_R output35 (.A(net37),
    .Y(dataadr[14]));
 BUFx2_ASAP7_75t_R output36 (.A(net38),
    .Y(dataadr[15]));
 BUFx2_ASAP7_75t_R output37 (.A(net39),
    .Y(dataadr[16]));
 BUFx2_ASAP7_75t_R output38 (.A(net40),
    .Y(dataadr[17]));
 BUFx2_ASAP7_75t_R output39 (.A(net41),
    .Y(dataadr[18]));
 BUFx2_ASAP7_75t_R output40 (.A(net42),
    .Y(dataadr[19]));
 BUFx2_ASAP7_75t_R output41 (.A(net43),
    .Y(dataadr[1]));
 BUFx2_ASAP7_75t_R output42 (.A(net44),
    .Y(dataadr[20]));
 BUFx2_ASAP7_75t_R output43 (.A(net45),
    .Y(dataadr[21]));
 BUFx2_ASAP7_75t_R output44 (.A(net46),
    .Y(dataadr[22]));
 BUFx2_ASAP7_75t_R output45 (.A(net47),
    .Y(dataadr[23]));
 BUFx2_ASAP7_75t_R output46 (.A(net48),
    .Y(dataadr[24]));
 BUFx2_ASAP7_75t_R output47 (.A(net49),
    .Y(dataadr[25]));
 BUFx2_ASAP7_75t_R output48 (.A(net50),
    .Y(dataadr[26]));
 BUFx2_ASAP7_75t_R output49 (.A(net51),
    .Y(dataadr[27]));
 BUFx2_ASAP7_75t_R output50 (.A(net52),
    .Y(dataadr[28]));
 BUFx2_ASAP7_75t_R output51 (.A(net53),
    .Y(dataadr[29]));
 BUFx2_ASAP7_75t_R output52 (.A(net54),
    .Y(dataadr[2]));
 BUFx2_ASAP7_75t_R output53 (.A(net55),
    .Y(dataadr[30]));
 BUFx2_ASAP7_75t_R output54 (.A(net56),
    .Y(dataadr[31]));
 BUFx2_ASAP7_75t_R output55 (.A(net57),
    .Y(dataadr[3]));
 BUFx2_ASAP7_75t_R output56 (.A(net58),
    .Y(dataadr[4]));
 BUFx2_ASAP7_75t_R output57 (.A(net59),
    .Y(dataadr[5]));
 BUFx2_ASAP7_75t_R output58 (.A(net60),
    .Y(dataadr[6]));
 BUFx2_ASAP7_75t_R output59 (.A(net61),
    .Y(dataadr[7]));
 BUFx2_ASAP7_75t_R output60 (.A(net62),
    .Y(dataadr[8]));
 BUFx2_ASAP7_75t_R output61 (.A(net63),
    .Y(dataadr[9]));
 BUFx2_ASAP7_75t_R output62 (.A(net64),
    .Y(memwrite));
 BUFx2_ASAP7_75t_R output63 (.A(net65),
    .Y(pc[0]));
 BUFx2_ASAP7_75t_R output64 (.A(net66),
    .Y(pc[10]));
 BUFx2_ASAP7_75t_R output65 (.A(net67),
    .Y(pc[11]));
 BUFx2_ASAP7_75t_R output66 (.A(net68),
    .Y(pc[12]));
 BUFx2_ASAP7_75t_R output67 (.A(net69),
    .Y(pc[13]));
 BUFx2_ASAP7_75t_R output68 (.A(net70),
    .Y(pc[14]));
 BUFx2_ASAP7_75t_R output69 (.A(net71),
    .Y(pc[15]));
 BUFx2_ASAP7_75t_R output70 (.A(net72),
    .Y(pc[16]));
 BUFx2_ASAP7_75t_R output71 (.A(net73),
    .Y(pc[17]));
 BUFx2_ASAP7_75t_R output72 (.A(net74),
    .Y(pc[18]));
 BUFx2_ASAP7_75t_R output73 (.A(net75),
    .Y(pc[19]));
 BUFx2_ASAP7_75t_R output74 (.A(net76),
    .Y(pc[1]));
 BUFx2_ASAP7_75t_R output75 (.A(net77),
    .Y(pc[20]));
 BUFx2_ASAP7_75t_R output76 (.A(net78),
    .Y(pc[21]));
 BUFx2_ASAP7_75t_R output77 (.A(net79),
    .Y(pc[22]));
 BUFx2_ASAP7_75t_R output78 (.A(net80),
    .Y(pc[23]));
 BUFx2_ASAP7_75t_R output79 (.A(net81),
    .Y(pc[24]));
 BUFx2_ASAP7_75t_R output80 (.A(net82),
    .Y(pc[25]));
 BUFx2_ASAP7_75t_R output81 (.A(net83),
    .Y(pc[26]));
 BUFx2_ASAP7_75t_R output82 (.A(net84),
    .Y(pc[27]));
 BUFx2_ASAP7_75t_R output83 (.A(net85),
    .Y(pc[28]));
 BUFx2_ASAP7_75t_R output84 (.A(net86),
    .Y(pc[29]));
 BUFx2_ASAP7_75t_R output85 (.A(net87),
    .Y(pc[2]));
 BUFx2_ASAP7_75t_R output86 (.A(net88),
    .Y(pc[30]));
 BUFx2_ASAP7_75t_R output87 (.A(net89),
    .Y(pc[31]));
 BUFx2_ASAP7_75t_R output88 (.A(net90),
    .Y(pc[3]));
 BUFx2_ASAP7_75t_R output89 (.A(net91),
    .Y(pc[4]));
 BUFx2_ASAP7_75t_R output90 (.A(net92),
    .Y(pc[5]));
 BUFx2_ASAP7_75t_R output91 (.A(net93),
    .Y(pc[6]));
 BUFx2_ASAP7_75t_R output92 (.A(net94),
    .Y(pc[7]));
 BUFx2_ASAP7_75t_R output93 (.A(net95),
    .Y(pc[8]));
 BUFx2_ASAP7_75t_R output94 (.A(net96),
    .Y(pc[9]));
 BUFx2_ASAP7_75t_R output95 (.A(net97),
    .Y(ready));
 BUFx2_ASAP7_75t_R output96 (.A(net98),
    .Y(suspend));
 BUFx2_ASAP7_75t_R output97 (.A(net99),
    .Y(writedata[0]));
 BUFx2_ASAP7_75t_R output98 (.A(net100),
    .Y(writedata[10]));
 BUFx2_ASAP7_75t_R output99 (.A(net101),
    .Y(writedata[11]));
 BUFx2_ASAP7_75t_R output100 (.A(net102),
    .Y(writedata[12]));
 BUFx2_ASAP7_75t_R output101 (.A(net103),
    .Y(writedata[13]));
 BUFx2_ASAP7_75t_R output102 (.A(net104),
    .Y(writedata[14]));
 BUFx2_ASAP7_75t_R output103 (.A(net105),
    .Y(writedata[15]));
 BUFx2_ASAP7_75t_R output104 (.A(net106),
    .Y(writedata[16]));
 BUFx2_ASAP7_75t_R output105 (.A(net107),
    .Y(writedata[17]));
 BUFx2_ASAP7_75t_R output106 (.A(net108),
    .Y(writedata[18]));
 BUFx2_ASAP7_75t_R output107 (.A(net109),
    .Y(writedata[19]));
 BUFx2_ASAP7_75t_R output108 (.A(net110),
    .Y(writedata[1]));
 BUFx2_ASAP7_75t_R output109 (.A(net111),
    .Y(writedata[20]));
 BUFx2_ASAP7_75t_R output110 (.A(net112),
    .Y(writedata[21]));
 BUFx2_ASAP7_75t_R output111 (.A(net113),
    .Y(writedata[22]));
 BUFx2_ASAP7_75t_R output112 (.A(net114),
    .Y(writedata[23]));
 BUFx2_ASAP7_75t_R output113 (.A(net115),
    .Y(writedata[24]));
 BUFx2_ASAP7_75t_R output114 (.A(net116),
    .Y(writedata[25]));
 BUFx2_ASAP7_75t_R output115 (.A(net117),
    .Y(writedata[26]));
 BUFx2_ASAP7_75t_R output116 (.A(net118),
    .Y(writedata[27]));
 BUFx2_ASAP7_75t_R output117 (.A(net119),
    .Y(writedata[28]));
 BUFx2_ASAP7_75t_R output118 (.A(net120),
    .Y(writedata[29]));
 BUFx2_ASAP7_75t_R output119 (.A(net121),
    .Y(writedata[2]));
 BUFx2_ASAP7_75t_R output120 (.A(net122),
    .Y(writedata[30]));
 BUFx2_ASAP7_75t_R output121 (.A(net123),
    .Y(writedata[31]));
 BUFx2_ASAP7_75t_R output122 (.A(net124),
    .Y(writedata[3]));
 BUFx2_ASAP7_75t_R output123 (.A(net167),
    .Y(writedata[4]));
 BUFx2_ASAP7_75t_R output124 (.A(net126),
    .Y(writedata[5]));
 BUFx2_ASAP7_75t_R output125 (.A(net127),
    .Y(writedata[6]));
 BUFx2_ASAP7_75t_R output126 (.A(net128),
    .Y(writedata[7]));
 BUFx2_ASAP7_75t_R output127 (.A(net129),
    .Y(writedata[8]));
 BUFx2_ASAP7_75t_R output128 (.A(net130),
    .Y(writedata[9]));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[0]$_DFFE_PP0P__129  (.H(net131));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[10]$_DFF_PP0__130  (.H(net132));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[11]$_DFF_PP0__131  (.H(net133));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[12]$_DFF_PP0__132  (.H(net134));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[13]$_DFF_PP0__133  (.H(net135));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[14]$_DFF_PP0__134  (.H(net136));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[15]$_DFF_PP0__135  (.H(net137));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[16]$_DFF_PP0__136  (.H(net138));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[17]$_DFF_PP0__137  (.H(net139));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[18]$_DFF_PP0__138  (.H(net140));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[19]$_DFF_PP0__139  (.H(net141));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[1]$_DFFE_PP0P__140  (.H(net142));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[20]$_DFF_PP0__141  (.H(net143));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[21]$_DFF_PP0__142  (.H(net144));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[22]$_DFF_PP0__143  (.H(net145));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[23]$_DFF_PP0__144  (.H(net146));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[24]$_DFF_PP0__145  (.H(net147));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[25]$_DFF_PP0__146  (.H(net148));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[26]$_DFF_PP0__147  (.H(net149));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[27]$_DFF_PP0__148  (.H(net150));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[28]$_DFF_PP0__149  (.H(net151));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[29]$_DFF_PP0__150  (.H(net152));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[2]$_DFF_PP0__151  (.H(net153));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[30]$_DFF_PP0__152  (.H(net154));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[31]$_DFF_PP0__153  (.H(net155));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[3]$_DFF_PP0__154  (.H(net156));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[4]$_DFF_PP0__155  (.H(net157));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[5]$_DFF_PP0__156  (.H(net158));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[6]$_DFF_PP0__157  (.H(net159));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[7]$_DFF_PP0__158  (.H(net160));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[8]$_DFF_PP0__159  (.H(net161));
 TIEHIx1_ASAP7_75t_R \riscv.dp.pcreg.q[9]$_DFF_PP0__160  (.H(net162));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_1_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_2_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_3_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_4_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_8_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_11_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_14_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_15_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_18_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_19_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_21_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_23_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_24_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_25_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_26_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_27_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_28_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_28_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_29_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_29_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_30_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_30_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_31_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_31_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_32_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_32_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_33_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_33_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_34_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_34_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_35_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_35_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_36_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_36_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_37_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_37_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_38_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_38_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_39_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_39_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_40_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_40_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_41_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_41_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_42_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_42_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_43_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_43_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_44_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_44_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_45_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_45_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_46_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_46_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_47_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_47_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_48_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_48_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_49_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_49_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_50_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_50_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_51_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_51_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_52_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_52_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_53_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_53_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_54_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_54_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_55_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_55_clk));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_0_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_1_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_2_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_3_0_clk));
 CKINVDCx20_ASAP7_75t_R clkload0 (.A(clknet_2_0_0_clk));
 CKINVDCx20_ASAP7_75t_R clkload1 (.A(clknet_2_1_0_clk));
 CKINVDCx20_ASAP7_75t_R clkload2 (.A(clknet_2_3_0_clk));
 CKINVDCx10_ASAP7_75t_R clkload3 (.A(clknet_leaf_0_clk));
 BUFx4f_ASAP7_75t_R clkload4 (.A(clknet_leaf_1_clk));
 BUFx4f_ASAP7_75t_R clkload5 (.A(clknet_leaf_2_clk));
 BUFx24_ASAP7_75t_R clkload6 (.A(clknet_leaf_3_clk));
 CKINVDCx20_ASAP7_75t_R clkload7 (.A(clknet_leaf_4_clk));
 INVx8_ASAP7_75t_R clkload8 (.A(clknet_leaf_43_clk));
 BUFx24_ASAP7_75t_R clkload9 (.A(clknet_leaf_44_clk));
 INVx3_ASAP7_75t_R clkload10 (.A(clknet_leaf_45_clk));
 CKINVDCx9p33_ASAP7_75t_R clkload11 (.A(clknet_leaf_46_clk));
 BUFx24_ASAP7_75t_R clkload12 (.A(clknet_leaf_47_clk));
 BUFx12_ASAP7_75t_R clkload13 (.A(clknet_leaf_48_clk));
 INVxp67_ASAP7_75t_R clkload14 (.A(clknet_leaf_50_clk));
 BUFx12_ASAP7_75t_R clkload15 (.A(clknet_leaf_51_clk));
 INVx3_ASAP7_75t_R clkload16 (.A(clknet_leaf_52_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload17 (.A(clknet_leaf_53_clk));
 CKINVDCx11_ASAP7_75t_R clkload18 (.A(clknet_leaf_54_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload19 (.A(clknet_leaf_55_clk));
 BUFx4f_ASAP7_75t_R clkload20 (.A(clknet_leaf_28_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload21 (.A(clknet_leaf_29_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload22 (.A(clknet_leaf_30_clk));
 BUFx24_ASAP7_75t_R clkload23 (.A(clknet_leaf_31_clk));
 BUFx4f_ASAP7_75t_R clkload24 (.A(clknet_leaf_32_clk));
 INVxp67_ASAP7_75t_R clkload25 (.A(clknet_leaf_34_clk));
 BUFx24_ASAP7_75t_R clkload26 (.A(clknet_leaf_35_clk));
 INVx5_ASAP7_75t_R clkload27 (.A(clknet_leaf_36_clk));
 INVx3_ASAP7_75t_R clkload28 (.A(clknet_leaf_37_clk));
 BUFx24_ASAP7_75t_R clkload29 (.A(clknet_leaf_38_clk));
 INVx3_ASAP7_75t_R clkload30 (.A(clknet_leaf_39_clk));
 INVx3_ASAP7_75t_R clkload31 (.A(clknet_leaf_40_clk));
 BUFx4f_ASAP7_75t_R clkload32 (.A(clknet_leaf_41_clk));
 CKINVDCx8_ASAP7_75t_R clkload33 (.A(clknet_leaf_42_clk));
 CKINVDCx14_ASAP7_75t_R clkload34 (.A(clknet_leaf_8_clk));
 BUFx12_ASAP7_75t_R clkload35 (.A(clknet_leaf_10_clk));
 INVx5_ASAP7_75t_R clkload36 (.A(clknet_leaf_11_clk));
 BUFx4f_ASAP7_75t_R clkload37 (.A(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkload38 (.A(clknet_leaf_22_clk));
 INVxp67_ASAP7_75t_R clkload39 (.A(clknet_leaf_12_clk));
 BUFx12_ASAP7_75t_R clkload40 (.A(clknet_leaf_15_clk));
 INVx3_ASAP7_75t_R clkload41 (.A(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkload42 (.A(clknet_leaf_18_clk));
 INVx6_ASAP7_75t_R clkload43 (.A(clknet_leaf_19_clk));
 INVx3_ASAP7_75t_R clkload44 (.A(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkload45 (.A(clknet_leaf_21_clk));
 INVx5_ASAP7_75t_R clkload46 (.A(clknet_leaf_23_clk));
 CKINVDCx11_ASAP7_75t_R clkload47 (.A(clknet_leaf_24_clk));
 BUFx24_ASAP7_75t_R clkload48 (.A(clknet_leaf_25_clk));
 INVx8_ASAP7_75t_R clkload49 (.A(clknet_leaf_26_clk));
 BUFx4f_ASAP7_75t_R clkload50 (.A(clknet_leaf_27_clk));
 BUFx3_ASAP7_75t_R rebuffer1 (.A(_01031_),
    .Y(net163));
 BUFx2_ASAP7_75t_R rebuffer2 (.A(net163),
    .Y(net164));
 BUFx2_ASAP7_75t_R rebuffer3 (.A(net125),
    .Y(net165));
 BUFx6f_ASAP7_75t_R rebuffer4 (.A(net165),
    .Y(net166));
 BUFx2_ASAP7_75t_R rebuffer5 (.A(net125),
    .Y(net167));
 BUFx6f_ASAP7_75t_R rebuffer6 (.A(_01157_),
    .Y(net168));
 BUFx2_ASAP7_75t_R rebuffer7 (.A(net168),
    .Y(net169));
 BUFx2_ASAP7_75t_R rebuffer8 (.A(net169),
    .Y(net170));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144 ();
 DECAPx6_ASAP7_75t_R FILLER_0_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186 ();
 DECAPx6_ASAP7_75t_R FILLER_0_192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212 ();
 FILLER_ASAP7_75t_R FILLER_0_376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_428 ();
 DECAPx2_ASAP7_75t_R FILLER_0_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_575 ();
 DECAPx1_ASAP7_75t_R FILLER_0_591 ();
 DECAPx4_ASAP7_75t_R FILLER_0_616 ();
 FILLER_ASAP7_75t_R FILLER_0_626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_651 ();
 DECAPx10_ASAP7_75t_R FILLER_0_673 ();
 DECAPx10_ASAP7_75t_R FILLER_0_695 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_755 ();
 DECAPx1_ASAP7_75t_R FILLER_0_777 ();
 DECAPx4_ASAP7_75t_R FILLER_0_795 ();
 FILLER_ASAP7_75t_R FILLER_0_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_816 ();
 DECAPx2_ASAP7_75t_R FILLER_0_838 ();
 FILLER_ASAP7_75t_R FILLER_0_844 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851 ();
 DECAPx2_ASAP7_75t_R FILLER_0_873 ();
 FILLER_ASAP7_75t_R FILLER_0_879 ();
 DECAPx6_ASAP7_75t_R FILLER_0_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_909 ();
 DECAPx1_ASAP7_75t_R FILLER_0_920 ();
 DECAPx6_ASAP7_75t_R FILLER_0_926 ();
 DECAPx1_ASAP7_75t_R FILLER_0_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_944 ();
 DECAPx10_ASAP7_75t_R FILLER_0_958 ();
 DECAPx10_ASAP7_75t_R FILLER_0_980 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1189 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx4_ASAP7_75t_R FILLER_1_178 ();
 FILLER_ASAP7_75t_R FILLER_1_188 ();
 FILLER_ASAP7_75t_R FILLER_1_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_392 ();
 FILLER_ASAP7_75t_R FILLER_1_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_571 ();
 FILLER_ASAP7_75t_R FILLER_1_593 ();
 DECAPx6_ASAP7_75t_R FILLER_1_602 ();
 DECAPx10_ASAP7_75t_R FILLER_1_637 ();
 DECAPx10_ASAP7_75t_R FILLER_1_659 ();
 DECAPx10_ASAP7_75t_R FILLER_1_681 ();
 DECAPx10_ASAP7_75t_R FILLER_1_703 ();
 DECAPx4_ASAP7_75t_R FILLER_1_746 ();
 FILLER_ASAP7_75t_R FILLER_1_756 ();
 DECAPx4_ASAP7_75t_R FILLER_1_765 ();
 FILLER_ASAP7_75t_R FILLER_1_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_777 ();
 FILLER_ASAP7_75t_R FILLER_1_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_801 ();
 DECAPx2_ASAP7_75t_R FILLER_1_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_857 ();
 DECAPx1_ASAP7_75t_R FILLER_1_868 ();
 DECAPx10_ASAP7_75t_R FILLER_1_888 ();
 FILLER_ASAP7_75t_R FILLER_1_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_912 ();
 FILLER_ASAP7_75t_R FILLER_1_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_992 ();
 FILLER_ASAP7_75t_R FILLER_1_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1037 ();
 FILLER_ASAP7_75t_R FILLER_1_1043 ();
 FILLER_ASAP7_75t_R FILLER_1_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1120 ();
 FILLER_ASAP7_75t_R FILLER_1_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_1_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1168 ();
 DECAPx1_ASAP7_75t_R FILLER_1_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 FILLER_ASAP7_75t_R FILLER_2_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_316 ();
 FILLER_ASAP7_75t_R FILLER_2_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_396 ();
 FILLER_ASAP7_75t_R FILLER_2_402 ();
 FILLER_ASAP7_75t_R FILLER_2_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_421 ();
 FILLER_ASAP7_75t_R FILLER_2_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_434 ();
 FILLER_ASAP7_75t_R FILLER_2_457 ();
 DECAPx4_ASAP7_75t_R FILLER_2_492 ();
 FILLER_ASAP7_75t_R FILLER_2_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_504 ();
 FILLER_ASAP7_75t_R FILLER_2_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_542 ();
 FILLER_ASAP7_75t_R FILLER_2_548 ();
 FILLER_ASAP7_75t_R FILLER_2_557 ();
 FILLER_ASAP7_75t_R FILLER_2_569 ();
 DECAPx4_ASAP7_75t_R FILLER_2_578 ();
 FILLER_ASAP7_75t_R FILLER_2_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_590 ();
 DECAPx1_ASAP7_75t_R FILLER_2_601 ();
 DECAPx1_ASAP7_75t_R FILLER_2_626 ();
 DECAPx10_ASAP7_75t_R FILLER_2_651 ();
 DECAPx10_ASAP7_75t_R FILLER_2_673 ();
 DECAPx10_ASAP7_75t_R FILLER_2_695 ();
 DECAPx4_ASAP7_75t_R FILLER_2_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_727 ();
 DECAPx4_ASAP7_75t_R FILLER_2_745 ();
 FILLER_ASAP7_75t_R FILLER_2_755 ();
 FILLER_ASAP7_75t_R FILLER_2_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_769 ();
 DECAPx2_ASAP7_75t_R FILLER_2_784 ();
 FILLER_ASAP7_75t_R FILLER_2_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_798 ();
 DECAPx1_ASAP7_75t_R FILLER_2_844 ();
 DECAPx10_ASAP7_75t_R FILLER_2_879 ();
 DECAPx6_ASAP7_75t_R FILLER_2_901 ();
 FILLER_ASAP7_75t_R FILLER_2_915 ();
 DECAPx10_ASAP7_75t_R FILLER_2_938 ();
 FILLER_ASAP7_75t_R FILLER_2_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_984 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_2_1019 ();
 FILLER_ASAP7_75t_R FILLER_2_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1031 ();
 FILLER_ASAP7_75t_R FILLER_2_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1192 ();
 FILLER_ASAP7_75t_R FILLER_2_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_2_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx2_ASAP7_75t_R FILLER_3_134 ();
 FILLER_ASAP7_75t_R FILLER_3_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_142 ();
 DECAPx2_ASAP7_75t_R FILLER_3_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_349 ();
 FILLER_ASAP7_75t_R FILLER_3_399 ();
 FILLER_ASAP7_75t_R FILLER_3_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_423 ();
 DECAPx1_ASAP7_75t_R FILLER_3_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_438 ();
 DECAPx1_ASAP7_75t_R FILLER_3_477 ();
 FILLER_ASAP7_75t_R FILLER_3_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_530 ();
 FILLER_ASAP7_75t_R FILLER_3_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_550 ();
 DECAPx6_ASAP7_75t_R FILLER_3_566 ();
 FILLER_ASAP7_75t_R FILLER_3_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_582 ();
 DECAPx10_ASAP7_75t_R FILLER_3_610 ();
 FILLER_ASAP7_75t_R FILLER_3_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_634 ();
 DECAPx10_ASAP7_75t_R FILLER_3_642 ();
 DECAPx1_ASAP7_75t_R FILLER_3_664 ();
 DECAPx10_ASAP7_75t_R FILLER_3_682 ();
 DECAPx10_ASAP7_75t_R FILLER_3_704 ();
 DECAPx1_ASAP7_75t_R FILLER_3_726 ();
 DECAPx4_ASAP7_75t_R FILLER_3_758 ();
 FILLER_ASAP7_75t_R FILLER_3_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_794 ();
 DECAPx6_ASAP7_75t_R FILLER_3_811 ();
 FILLER_ASAP7_75t_R FILLER_3_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_868 ();
 DECAPx10_ASAP7_75t_R FILLER_3_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_926 ();
 DECAPx2_ASAP7_75t_R FILLER_3_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_943 ();
 DECAPx4_ASAP7_75t_R FILLER_3_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1032 ();
 FILLER_ASAP7_75t_R FILLER_3_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1086 ();
 FILLER_ASAP7_75t_R FILLER_3_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1125 ();
 FILLER_ASAP7_75t_R FILLER_3_1139 ();
 FILLER_ASAP7_75t_R FILLER_3_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1167 ();
 FILLER_ASAP7_75t_R FILLER_3_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1205 ();
 FILLER_ASAP7_75t_R FILLER_3_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx4_ASAP7_75t_R FILLER_4_112 ();
 FILLER_ASAP7_75t_R FILLER_4_122 ();
 DECAPx10_ASAP7_75t_R FILLER_4_127 ();
 DECAPx2_ASAP7_75t_R FILLER_4_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_155 ();
 FILLER_ASAP7_75t_R FILLER_4_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_161 ();
 FILLER_ASAP7_75t_R FILLER_4_196 ();
 FILLER_ASAP7_75t_R FILLER_4_210 ();
 FILLER_ASAP7_75t_R FILLER_4_243 ();
 FILLER_ASAP7_75t_R FILLER_4_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_296 ();
 FILLER_ASAP7_75t_R FILLER_4_334 ();
 FILLER_ASAP7_75t_R FILLER_4_365 ();
 FILLER_ASAP7_75t_R FILLER_4_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_417 ();
 FILLER_ASAP7_75t_R FILLER_4_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_441 ();
 DECAPx4_ASAP7_75t_R FILLER_4_452 ();
 DECAPx4_ASAP7_75t_R FILLER_4_464 ();
 FILLER_ASAP7_75t_R FILLER_4_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_476 ();
 DECAPx6_ASAP7_75t_R FILLER_4_484 ();
 DECAPx1_ASAP7_75t_R FILLER_4_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_523 ();
 DECAPx4_ASAP7_75t_R FILLER_4_608 ();
 DECAPx10_ASAP7_75t_R FILLER_4_645 ();
 DECAPx10_ASAP7_75t_R FILLER_4_667 ();
 DECAPx10_ASAP7_75t_R FILLER_4_689 ();
 DECAPx2_ASAP7_75t_R FILLER_4_711 ();
 FILLER_ASAP7_75t_R FILLER_4_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_719 ();
 DECAPx6_ASAP7_75t_R FILLER_4_730 ();
 DECAPx1_ASAP7_75t_R FILLER_4_744 ();
 DECAPx6_ASAP7_75t_R FILLER_4_758 ();
 DECAPx1_ASAP7_75t_R FILLER_4_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_776 ();
 DECAPx6_ASAP7_75t_R FILLER_4_798 ();
 FILLER_ASAP7_75t_R FILLER_4_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_814 ();
 DECAPx10_ASAP7_75t_R FILLER_4_829 ();
 DECAPx10_ASAP7_75t_R FILLER_4_851 ();
 DECAPx6_ASAP7_75t_R FILLER_4_873 ();
 FILLER_ASAP7_75t_R FILLER_4_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_889 ();
 DECAPx10_ASAP7_75t_R FILLER_4_897 ();
 DECAPx6_ASAP7_75t_R FILLER_4_919 ();
 DECAPx1_ASAP7_75t_R FILLER_4_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_974 ();
 DECAPx10_ASAP7_75t_R FILLER_4_981 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1165 ();
 FILLER_ASAP7_75t_R FILLER_4_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx6_ASAP7_75t_R FILLER_5_90 ();
 DECAPx2_ASAP7_75t_R FILLER_5_104 ();
 DECAPx6_ASAP7_75t_R FILLER_5_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_150 ();
 DECAPx6_ASAP7_75t_R FILLER_5_156 ();
 FILLER_ASAP7_75t_R FILLER_5_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_172 ();
 DECAPx2_ASAP7_75t_R FILLER_5_176 ();
 FILLER_ASAP7_75t_R FILLER_5_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_189 ();
 FILLER_ASAP7_75t_R FILLER_5_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_226 ();
 FILLER_ASAP7_75t_R FILLER_5_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_257 ();
 FILLER_ASAP7_75t_R FILLER_5_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_360 ();
 FILLER_ASAP7_75t_R FILLER_5_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_408 ();
 DECAPx2_ASAP7_75t_R FILLER_5_414 ();
 FILLER_ASAP7_75t_R FILLER_5_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_437 ();
 DECAPx1_ASAP7_75t_R FILLER_5_445 ();
 DECAPx1_ASAP7_75t_R FILLER_5_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_502 ();
 DECAPx1_ASAP7_75t_R FILLER_5_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_514 ();
 DECAPx2_ASAP7_75t_R FILLER_5_525 ();
 FILLER_ASAP7_75t_R FILLER_5_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_533 ();
 DECAPx1_ASAP7_75t_R FILLER_5_544 ();
 DECAPx2_ASAP7_75t_R FILLER_5_555 ();
 FILLER_ASAP7_75t_R FILLER_5_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_563 ();
 DECAPx2_ASAP7_75t_R FILLER_5_581 ();
 FILLER_ASAP7_75t_R FILLER_5_587 ();
 DECAPx2_ASAP7_75t_R FILLER_5_596 ();
 FILLER_ASAP7_75t_R FILLER_5_602 ();
 DECAPx10_ASAP7_75t_R FILLER_5_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_636 ();
 DECAPx10_ASAP7_75t_R FILLER_5_644 ();
 DECAPx10_ASAP7_75t_R FILLER_5_666 ();
 DECAPx4_ASAP7_75t_R FILLER_5_688 ();
 FILLER_ASAP7_75t_R FILLER_5_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_700 ();
 DECAPx6_ASAP7_75t_R FILLER_5_711 ();
 FILLER_ASAP7_75t_R FILLER_5_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_727 ();
 DECAPx6_ASAP7_75t_R FILLER_5_738 ();
 DECAPx1_ASAP7_75t_R FILLER_5_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_756 ();
 DECAPx2_ASAP7_75t_R FILLER_5_778 ();
 FILLER_ASAP7_75t_R FILLER_5_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_786 ();
 DECAPx1_ASAP7_75t_R FILLER_5_794 ();
 FILLER_ASAP7_75t_R FILLER_5_811 ();
 DECAPx10_ASAP7_75t_R FILLER_5_848 ();
 DECAPx10_ASAP7_75t_R FILLER_5_870 ();
 DECAPx10_ASAP7_75t_R FILLER_5_892 ();
 DECAPx4_ASAP7_75t_R FILLER_5_914 ();
 DECAPx4_ASAP7_75t_R FILLER_5_926 ();
 FILLER_ASAP7_75t_R FILLER_5_936 ();
 DECAPx2_ASAP7_75t_R FILLER_5_955 ();
 DECAPx1_ASAP7_75t_R FILLER_5_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_995 ();
 FILLER_ASAP7_75t_R FILLER_5_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1018 ();
 FILLER_ASAP7_75t_R FILLER_5_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_5_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1126 ();
 FILLER_ASAP7_75t_R FILLER_5_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1134 ();
 FILLER_ASAP7_75t_R FILLER_5_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_5_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx6_ASAP7_75t_R FILLER_6_90 ();
 DECAPx2_ASAP7_75t_R FILLER_6_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_147 ();
 FILLER_ASAP7_75t_R FILLER_6_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_156 ();
 DECAPx2_ASAP7_75t_R FILLER_6_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_177 ();
 DECAPx2_ASAP7_75t_R FILLER_6_190 ();
 FILLER_ASAP7_75t_R FILLER_6_196 ();
 DECAPx4_ASAP7_75t_R FILLER_6_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_224 ();
 FILLER_ASAP7_75t_R FILLER_6_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_291 ();
 FILLER_ASAP7_75t_R FILLER_6_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_322 ();
 FILLER_ASAP7_75t_R FILLER_6_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_384 ();
 FILLER_ASAP7_75t_R FILLER_6_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_407 ();
 FILLER_ASAP7_75t_R FILLER_6_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_451 ();
 DECAPx10_ASAP7_75t_R FILLER_6_464 ();
 DECAPx6_ASAP7_75t_R FILLER_6_486 ();
 DECAPx1_ASAP7_75t_R FILLER_6_500 ();
 DECAPx10_ASAP7_75t_R FILLER_6_525 ();
 DECAPx6_ASAP7_75t_R FILLER_6_568 ();
 FILLER_ASAP7_75t_R FILLER_6_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_595 ();
 DECAPx4_ASAP7_75t_R FILLER_6_624 ();
 FILLER_ASAP7_75t_R FILLER_6_634 ();
 DECAPx10_ASAP7_75t_R FILLER_6_657 ();
 DECAPx10_ASAP7_75t_R FILLER_6_679 ();
 DECAPx2_ASAP7_75t_R FILLER_6_701 ();
 FILLER_ASAP7_75t_R FILLER_6_707 ();
 DECAPx4_ASAP7_75t_R FILLER_6_737 ();
 DECAPx10_ASAP7_75t_R FILLER_6_764 ();
 DECAPx2_ASAP7_75t_R FILLER_6_786 ();
 DECAPx2_ASAP7_75t_R FILLER_6_813 ();
 FILLER_ASAP7_75t_R FILLER_6_819 ();
 FILLER_ASAP7_75t_R FILLER_6_860 ();
 DECAPx10_ASAP7_75t_R FILLER_6_876 ();
 DECAPx4_ASAP7_75t_R FILLER_6_898 ();
 FILLER_ASAP7_75t_R FILLER_6_908 ();
 DECAPx4_ASAP7_75t_R FILLER_6_948 ();
 DECAPx1_ASAP7_75t_R FILLER_6_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_983 ();
 FILLER_ASAP7_75t_R FILLER_6_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1038 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1066 ();
 FILLER_ASAP7_75t_R FILLER_6_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1078 ();
 FILLER_ASAP7_75t_R FILLER_6_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1171 ();
 FILLER_ASAP7_75t_R FILLER_6_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1280 ();
 FILLER_ASAP7_75t_R FILLER_6_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx4_ASAP7_75t_R FILLER_7_112 ();
 FILLER_ASAP7_75t_R FILLER_7_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_132 ();
 FILLER_ASAP7_75t_R FILLER_7_154 ();
 DECAPx6_ASAP7_75t_R FILLER_7_168 ();
 DECAPx2_ASAP7_75t_R FILLER_7_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_196 ();
 DECAPx2_ASAP7_75t_R FILLER_7_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_217 ();
 DECAPx1_ASAP7_75t_R FILLER_7_225 ();
 DECAPx2_ASAP7_75t_R FILLER_7_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_242 ();
 FILLER_ASAP7_75t_R FILLER_7_283 ();
 DECAPx1_ASAP7_75t_R FILLER_7_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_301 ();
 DECAPx2_ASAP7_75t_R FILLER_7_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_337 ();
 DECAPx1_ASAP7_75t_R FILLER_7_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_347 ();
 FILLER_ASAP7_75t_R FILLER_7_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_358 ();
 FILLER_ASAP7_75t_R FILLER_7_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_374 ();
 DECAPx10_ASAP7_75t_R FILLER_7_396 ();
 DECAPx4_ASAP7_75t_R FILLER_7_418 ();
 DECAPx4_ASAP7_75t_R FILLER_7_456 ();
 DECAPx2_ASAP7_75t_R FILLER_7_497 ();
 FILLER_ASAP7_75t_R FILLER_7_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_520 ();
 DECAPx6_ASAP7_75t_R FILLER_7_531 ();
 FILLER_ASAP7_75t_R FILLER_7_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_547 ();
 FILLER_ASAP7_75t_R FILLER_7_558 ();
 DECAPx6_ASAP7_75t_R FILLER_7_581 ();
 DECAPx2_ASAP7_75t_R FILLER_7_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_640 ();
 DECAPx10_ASAP7_75t_R FILLER_7_651 ();
 DECAPx10_ASAP7_75t_R FILLER_7_673 ();
 DECAPx10_ASAP7_75t_R FILLER_7_695 ();
 FILLER_ASAP7_75t_R FILLER_7_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_741 ();
 DECAPx2_ASAP7_75t_R FILLER_7_749 ();
 FILLER_ASAP7_75t_R FILLER_7_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_757 ();
 DECAPx6_ASAP7_75t_R FILLER_7_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_798 ();
 FILLER_ASAP7_75t_R FILLER_7_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_822 ();
 DECAPx4_ASAP7_75t_R FILLER_7_844 ();
 FILLER_ASAP7_75t_R FILLER_7_854 ();
 FILLER_ASAP7_75t_R FILLER_7_862 ();
 DECAPx10_ASAP7_75t_R FILLER_7_880 ();
 DECAPx6_ASAP7_75t_R FILLER_7_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_923 ();
 FILLER_ASAP7_75t_R FILLER_7_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_949 ();
 DECAPx1_ASAP7_75t_R FILLER_7_971 ();
 DECAPx2_ASAP7_75t_R FILLER_7_989 ();
 DECAPx1_ASAP7_75t_R FILLER_7_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_7_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1123 ();
 FILLER_ASAP7_75t_R FILLER_7_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_7_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1186 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_7_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx4_ASAP7_75t_R FILLER_8_112 ();
 FILLER_ASAP7_75t_R FILLER_8_122 ();
 DECAPx1_ASAP7_75t_R FILLER_8_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_140 ();
 FILLER_ASAP7_75t_R FILLER_8_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_155 ();
 DECAPx2_ASAP7_75t_R FILLER_8_182 ();
 DECAPx2_ASAP7_75t_R FILLER_8_200 ();
 DECAPx6_ASAP7_75t_R FILLER_8_212 ();
 DECAPx1_ASAP7_75t_R FILLER_8_226 ();
 DECAPx2_ASAP7_75t_R FILLER_8_236 ();
 FILLER_ASAP7_75t_R FILLER_8_242 ();
 DECAPx1_ASAP7_75t_R FILLER_8_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_255 ();
 FILLER_ASAP7_75t_R FILLER_8_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_265 ();
 DECAPx1_ASAP7_75t_R FILLER_8_269 ();
 FILLER_ASAP7_75t_R FILLER_8_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_292 ();
 DECAPx1_ASAP7_75t_R FILLER_8_299 ();
 FILLER_ASAP7_75t_R FILLER_8_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_318 ();
 DECAPx2_ASAP7_75t_R FILLER_8_351 ();
 FILLER_ASAP7_75t_R FILLER_8_357 ();
 DECAPx6_ASAP7_75t_R FILLER_8_365 ();
 DECAPx1_ASAP7_75t_R FILLER_8_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_383 ();
 DECAPx6_ASAP7_75t_R FILLER_8_422 ();
 FILLER_ASAP7_75t_R FILLER_8_436 ();
 DECAPx1_ASAP7_75t_R FILLER_8_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_464 ();
 FILLER_ASAP7_75t_R FILLER_8_472 ();
 FILLER_ASAP7_75t_R FILLER_8_484 ();
 FILLER_ASAP7_75t_R FILLER_8_514 ();
 DECAPx1_ASAP7_75t_R FILLER_8_526 ();
 DECAPx4_ASAP7_75t_R FILLER_8_537 ();
 DECAPx2_ASAP7_75t_R FILLER_8_554 ();
 FILLER_ASAP7_75t_R FILLER_8_560 ();
 DECAPx1_ASAP7_75t_R FILLER_8_569 ();
 DECAPx2_ASAP7_75t_R FILLER_8_594 ();
 FILLER_ASAP7_75t_R FILLER_8_600 ();
 DECAPx4_ASAP7_75t_R FILLER_8_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_622 ();
 DECAPx10_ASAP7_75t_R FILLER_8_644 ();
 DECAPx4_ASAP7_75t_R FILLER_8_666 ();
 DECAPx6_ASAP7_75t_R FILLER_8_683 ();
 FILLER_ASAP7_75t_R FILLER_8_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_699 ();
 DECAPx10_ASAP7_75t_R FILLER_8_714 ();
 DECAPx6_ASAP7_75t_R FILLER_8_736 ();
 FILLER_ASAP7_75t_R FILLER_8_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_790 ();
 FILLER_ASAP7_75t_R FILLER_8_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_815 ();
 DECAPx4_ASAP7_75t_R FILLER_8_844 ();
 FILLER_ASAP7_75t_R FILLER_8_854 ();
 DECAPx4_ASAP7_75t_R FILLER_8_863 ();
 FILLER_ASAP7_75t_R FILLER_8_873 ();
 DECAPx2_ASAP7_75t_R FILLER_8_885 ();
 DECAPx4_ASAP7_75t_R FILLER_8_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_915 ();
 DECAPx2_ASAP7_75t_R FILLER_8_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_974 ();
 DECAPx2_ASAP7_75t_R FILLER_8_989 ();
 DECAPx4_ASAP7_75t_R FILLER_8_1015 ();
 FILLER_ASAP7_75t_R FILLER_8_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1044 ();
 FILLER_ASAP7_75t_R FILLER_8_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1140 ();
 FILLER_ASAP7_75t_R FILLER_8_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx6_ASAP7_75t_R FILLER_9_90 ();
 FILLER_ASAP7_75t_R FILLER_9_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_106 ();
 DECAPx2_ASAP7_75t_R FILLER_9_121 ();
 FILLER_ASAP7_75t_R FILLER_9_127 ();
 DECAPx1_ASAP7_75t_R FILLER_9_176 ();
 FILLER_ASAP7_75t_R FILLER_9_204 ();
 DECAPx2_ASAP7_75t_R FILLER_9_212 ();
 DECAPx1_ASAP7_75t_R FILLER_9_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_240 ();
 DECAPx4_ASAP7_75t_R FILLER_9_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_257 ();
 FILLER_ASAP7_75t_R FILLER_9_265 ();
 DECAPx2_ASAP7_75t_R FILLER_9_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_292 ();
 FILLER_ASAP7_75t_R FILLER_9_299 ();
 FILLER_ASAP7_75t_R FILLER_9_320 ();
 FILLER_ASAP7_75t_R FILLER_9_326 ();
 DECAPx6_ASAP7_75t_R FILLER_9_340 ();
 DECAPx1_ASAP7_75t_R FILLER_9_354 ();
 DECAPx10_ASAP7_75t_R FILLER_9_367 ();
 DECAPx2_ASAP7_75t_R FILLER_9_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_395 ();
 DECAPx4_ASAP7_75t_R FILLER_9_424 ();
 DECAPx2_ASAP7_75t_R FILLER_9_441 ();
 FILLER_ASAP7_75t_R FILLER_9_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_449 ();
 DECAPx10_ASAP7_75t_R FILLER_9_471 ();
 DECAPx4_ASAP7_75t_R FILLER_9_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_503 ();
 DECAPx2_ASAP7_75t_R FILLER_9_556 ();
 FILLER_ASAP7_75t_R FILLER_9_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_564 ();
 DECAPx6_ASAP7_75t_R FILLER_9_582 ();
 DECAPx2_ASAP7_75t_R FILLER_9_596 ();
 DECAPx6_ASAP7_75t_R FILLER_9_609 ();
 DECAPx2_ASAP7_75t_R FILLER_9_623 ();
 DECAPx10_ASAP7_75t_R FILLER_9_650 ();
 DECAPx10_ASAP7_75t_R FILLER_9_672 ();
 DECAPx6_ASAP7_75t_R FILLER_9_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_708 ();
 DECAPx4_ASAP7_75t_R FILLER_9_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_747 ();
 FILLER_ASAP7_75t_R FILLER_9_755 ();
 DECAPx2_ASAP7_75t_R FILLER_9_767 ();
 FILLER_ASAP7_75t_R FILLER_9_773 ();
 DECAPx1_ASAP7_75t_R FILLER_9_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_810 ();
 DECAPx1_ASAP7_75t_R FILLER_9_817 ();
 DECAPx2_ASAP7_75t_R FILLER_9_828 ();
 FILLER_ASAP7_75t_R FILLER_9_834 ();
 DECAPx4_ASAP7_75t_R FILLER_9_849 ();
 DECAPx1_ASAP7_75t_R FILLER_9_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_969 ();
 DECAPx6_ASAP7_75t_R FILLER_9_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_991 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_9_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_9_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1080 ();
 FILLER_ASAP7_75t_R FILLER_9_1094 ();
 FILLER_ASAP7_75t_R FILLER_9_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1111 ();
 FILLER_ASAP7_75t_R FILLER_9_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_9_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_9_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1218 ();
 FILLER_ASAP7_75t_R FILLER_9_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_9_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx6_ASAP7_75t_R FILLER_10_90 ();
 FILLER_ASAP7_75t_R FILLER_10_104 ();
 DECAPx1_ASAP7_75t_R FILLER_10_136 ();
 DECAPx6_ASAP7_75t_R FILLER_10_170 ();
 DECAPx4_ASAP7_75t_R FILLER_10_190 ();
 FILLER_ASAP7_75t_R FILLER_10_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_202 ();
 DECAPx2_ASAP7_75t_R FILLER_10_271 ();
 FILLER_ASAP7_75t_R FILLER_10_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_279 ();
 DECAPx2_ASAP7_75t_R FILLER_10_286 ();
 DECAPx2_ASAP7_75t_R FILLER_10_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_350 ();
 DECAPx10_ASAP7_75t_R FILLER_10_360 ();
 DECAPx10_ASAP7_75t_R FILLER_10_382 ();
 DECAPx2_ASAP7_75t_R FILLER_10_404 ();
 DECAPx1_ASAP7_75t_R FILLER_10_427 ();
 FILLER_ASAP7_75t_R FILLER_10_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_461 ();
 DECAPx2_ASAP7_75t_R FILLER_10_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_470 ();
 FILLER_ASAP7_75t_R FILLER_10_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_501 ();
 DECAPx1_ASAP7_75t_R FILLER_10_509 ();
 FILLER_ASAP7_75t_R FILLER_10_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_545 ();
 DECAPx2_ASAP7_75t_R FILLER_10_553 ();
 DECAPx1_ASAP7_75t_R FILLER_10_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_573 ();
 DECAPx1_ASAP7_75t_R FILLER_10_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_619 ();
 FILLER_ASAP7_75t_R FILLER_10_644 ();
 DECAPx10_ASAP7_75t_R FILLER_10_656 ();
 DECAPx10_ASAP7_75t_R FILLER_10_678 ();
 DECAPx10_ASAP7_75t_R FILLER_10_700 ();
 DECAPx2_ASAP7_75t_R FILLER_10_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_738 ();
 FILLER_ASAP7_75t_R FILLER_10_770 ();
 DECAPx4_ASAP7_75t_R FILLER_10_785 ();
 FILLER_ASAP7_75t_R FILLER_10_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_797 ();
 DECAPx6_ASAP7_75t_R FILLER_10_829 ();
 FILLER_ASAP7_75t_R FILLER_10_843 ();
 DECAPx2_ASAP7_75t_R FILLER_10_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_858 ();
 DECAPx10_ASAP7_75t_R FILLER_10_869 ();
 DECAPx6_ASAP7_75t_R FILLER_10_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_905 ();
 FILLER_ASAP7_75t_R FILLER_10_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_922 ();
 DECAPx1_ASAP7_75t_R FILLER_10_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_937 ();
 DECAPx10_ASAP7_75t_R FILLER_10_948 ();
 DECAPx10_ASAP7_75t_R FILLER_10_970 ();
 FILLER_ASAP7_75t_R FILLER_10_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1026 ();
 FILLER_ASAP7_75t_R FILLER_10_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_10_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1075 ();
 FILLER_ASAP7_75t_R FILLER_10_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1121 ();
 FILLER_ASAP7_75t_R FILLER_10_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1183 ();
 FILLER_ASAP7_75t_R FILLER_10_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_10_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx6_ASAP7_75t_R FILLER_11_90 ();
 DECAPx1_ASAP7_75t_R FILLER_11_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_108 ();
 DECAPx1_ASAP7_75t_R FILLER_11_135 ();
 FILLER_ASAP7_75t_R FILLER_11_161 ();
 DECAPx6_ASAP7_75t_R FILLER_11_172 ();
 DECAPx1_ASAP7_75t_R FILLER_11_198 ();
 DECAPx1_ASAP7_75t_R FILLER_11_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_226 ();
 FILLER_ASAP7_75t_R FILLER_11_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_245 ();
 FILLER_ASAP7_75t_R FILLER_11_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_257 ();
 FILLER_ASAP7_75t_R FILLER_11_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_303 ();
 FILLER_ASAP7_75t_R FILLER_11_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_380 ();
 FILLER_ASAP7_75t_R FILLER_11_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_391 ();
 DECAPx6_ASAP7_75t_R FILLER_11_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_414 ();
 DECAPx4_ASAP7_75t_R FILLER_11_422 ();
 FILLER_ASAP7_75t_R FILLER_11_432 ();
 DECAPx6_ASAP7_75t_R FILLER_11_467 ();
 FILLER_ASAP7_75t_R FILLER_11_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_483 ();
 DECAPx1_ASAP7_75t_R FILLER_11_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_498 ();
 DECAPx6_ASAP7_75t_R FILLER_11_530 ();
 FILLER_ASAP7_75t_R FILLER_11_544 ();
 DECAPx6_ASAP7_75t_R FILLER_11_567 ();
 DECAPx1_ASAP7_75t_R FILLER_11_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_585 ();
 DECAPx2_ASAP7_75t_R FILLER_11_593 ();
 DECAPx2_ASAP7_75t_R FILLER_11_609 ();
 FILLER_ASAP7_75t_R FILLER_11_615 ();
 DECAPx10_ASAP7_75t_R FILLER_11_668 ();
 DECAPx6_ASAP7_75t_R FILLER_11_690 ();
 FILLER_ASAP7_75t_R FILLER_11_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_706 ();
 DECAPx4_ASAP7_75t_R FILLER_11_745 ();
 FILLER_ASAP7_75t_R FILLER_11_755 ();
 FILLER_ASAP7_75t_R FILLER_11_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_780 ();
 DECAPx6_ASAP7_75t_R FILLER_11_788 ();
 FILLER_ASAP7_75t_R FILLER_11_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_812 ();
 DECAPx6_ASAP7_75t_R FILLER_11_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_842 ();
 DECAPx2_ASAP7_75t_R FILLER_11_850 ();
 FILLER_ASAP7_75t_R FILLER_11_862 ();
 DECAPx4_ASAP7_75t_R FILLER_11_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_884 ();
 DECAPx2_ASAP7_75t_R FILLER_11_918 ();
 DECAPx6_ASAP7_75t_R FILLER_11_933 ();
 DECAPx1_ASAP7_75t_R FILLER_11_947 ();
 DECAPx1_ASAP7_75t_R FILLER_11_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_971 ();
 FILLER_ASAP7_75t_R FILLER_11_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1005 ();
 FILLER_ASAP7_75t_R FILLER_11_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1065 ();
 FILLER_ASAP7_75t_R FILLER_11_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1095 ();
 FILLER_ASAP7_75t_R FILLER_11_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_11_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_11_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_12_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_112 ();
 DECAPx6_ASAP7_75t_R FILLER_12_123 ();
 DECAPx2_ASAP7_75t_R FILLER_12_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_169 ();
 DECAPx2_ASAP7_75t_R FILLER_12_196 ();
 DECAPx2_ASAP7_75t_R FILLER_12_233 ();
 DECAPx2_ASAP7_75t_R FILLER_12_245 ();
 DECAPx2_ASAP7_75t_R FILLER_12_279 ();
 FILLER_ASAP7_75t_R FILLER_12_291 ();
 DECAPx1_ASAP7_75t_R FILLER_12_300 ();
 DECAPx2_ASAP7_75t_R FILLER_12_323 ();
 FILLER_ASAP7_75t_R FILLER_12_329 ();
 DECAPx4_ASAP7_75t_R FILLER_12_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_353 ();
 FILLER_ASAP7_75t_R FILLER_12_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_401 ();
 FILLER_ASAP7_75t_R FILLER_12_433 ();
 DECAPx2_ASAP7_75t_R FILLER_12_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_471 ();
 DECAPx2_ASAP7_75t_R FILLER_12_482 ();
 DECAPx6_ASAP7_75t_R FILLER_12_496 ();
 FILLER_ASAP7_75t_R FILLER_12_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_512 ();
 DECAPx2_ASAP7_75t_R FILLER_12_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_526 ();
 DECAPx1_ASAP7_75t_R FILLER_12_555 ();
 DECAPx4_ASAP7_75t_R FILLER_12_580 ();
 FILLER_ASAP7_75t_R FILLER_12_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_592 ();
 DECAPx1_ASAP7_75t_R FILLER_12_621 ();
 FILLER_ASAP7_75t_R FILLER_12_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_637 ();
 DECAPx10_ASAP7_75t_R FILLER_12_668 ();
 DECAPx6_ASAP7_75t_R FILLER_12_690 ();
 DECAPx1_ASAP7_75t_R FILLER_12_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_708 ();
 DECAPx4_ASAP7_75t_R FILLER_12_733 ();
 DECAPx10_ASAP7_75t_R FILLER_12_760 ();
 DECAPx6_ASAP7_75t_R FILLER_12_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_796 ();
 DECAPx2_ASAP7_75t_R FILLER_12_811 ();
 DECAPx1_ASAP7_75t_R FILLER_12_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_873 ();
 DECAPx6_ASAP7_75t_R FILLER_12_904 ();
 FILLER_ASAP7_75t_R FILLER_12_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_920 ();
 FILLER_ASAP7_75t_R FILLER_12_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_944 ();
 DECAPx6_ASAP7_75t_R FILLER_12_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_986 ();
 DECAPx6_ASAP7_75t_R FILLER_12_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1022 ();
 FILLER_ASAP7_75t_R FILLER_12_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_12_1091 ();
 FILLER_ASAP7_75t_R FILLER_12_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_12_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1158 ();
 FILLER_ASAP7_75t_R FILLER_12_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_12_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1268 ();
 FILLER_ASAP7_75t_R FILLER_12_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_13_68 ();
 DECAPx6_ASAP7_75t_R FILLER_13_90 ();
 DECAPx2_ASAP7_75t_R FILLER_13_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_110 ();
 DECAPx4_ASAP7_75t_R FILLER_13_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_145 ();
 FILLER_ASAP7_75t_R FILLER_13_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_161 ();
 DECAPx4_ASAP7_75t_R FILLER_13_188 ();
 FILLER_ASAP7_75t_R FILLER_13_198 ();
 FILLER_ASAP7_75t_R FILLER_13_212 ();
 FILLER_ASAP7_75t_R FILLER_13_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_222 ();
 DECAPx10_ASAP7_75t_R FILLER_13_230 ();
 DECAPx2_ASAP7_75t_R FILLER_13_252 ();
 FILLER_ASAP7_75t_R FILLER_13_258 ();
 DECAPx4_ASAP7_75t_R FILLER_13_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_283 ();
 DECAPx4_ASAP7_75t_R FILLER_13_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_312 ();
 FILLER_ASAP7_75t_R FILLER_13_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_487 ();
 FILLER_ASAP7_75t_R FILLER_13_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_497 ();
 FILLER_ASAP7_75t_R FILLER_13_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_510 ();
 DECAPx2_ASAP7_75t_R FILLER_13_532 ();
 FILLER_ASAP7_75t_R FILLER_13_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_540 ();
 DECAPx1_ASAP7_75t_R FILLER_13_569 ();
 DECAPx10_ASAP7_75t_R FILLER_13_604 ();
 DECAPx4_ASAP7_75t_R FILLER_13_626 ();
 FILLER_ASAP7_75t_R FILLER_13_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_638 ();
 DECAPx4_ASAP7_75t_R FILLER_13_660 ();
 FILLER_ASAP7_75t_R FILLER_13_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_672 ();
 DECAPx6_ASAP7_75t_R FILLER_13_683 ();
 FILLER_ASAP7_75t_R FILLER_13_697 ();
 DECAPx1_ASAP7_75t_R FILLER_13_705 ();
 DECAPx1_ASAP7_75t_R FILLER_13_735 ();
 DECAPx4_ASAP7_75t_R FILLER_13_767 ();
 FILLER_ASAP7_75t_R FILLER_13_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_793 ();
 DECAPx2_ASAP7_75t_R FILLER_13_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_832 ();
 DECAPx2_ASAP7_75t_R FILLER_13_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_850 ();
 DECAPx1_ASAP7_75t_R FILLER_13_864 ();
 FILLER_ASAP7_75t_R FILLER_13_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_891 ();
 DECAPx4_ASAP7_75t_R FILLER_13_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_923 ();
 DECAPx6_ASAP7_75t_R FILLER_13_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_940 ();
 FILLER_ASAP7_75t_R FILLER_13_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_964 ();
 DECAPx4_ASAP7_75t_R FILLER_13_986 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1024 ();
 FILLER_ASAP7_75t_R FILLER_13_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_13_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_13_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1154 ();
 FILLER_ASAP7_75t_R FILLER_13_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_14_68 ();
 DECAPx10_ASAP7_75t_R FILLER_14_90 ();
 DECAPx4_ASAP7_75t_R FILLER_14_112 ();
 DECAPx6_ASAP7_75t_R FILLER_14_125 ();
 DECAPx1_ASAP7_75t_R FILLER_14_139 ();
 FILLER_ASAP7_75t_R FILLER_14_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_156 ();
 FILLER_ASAP7_75t_R FILLER_14_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_165 ();
 FILLER_ASAP7_75t_R FILLER_14_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_187 ();
 FILLER_ASAP7_75t_R FILLER_14_200 ();
 DECAPx4_ASAP7_75t_R FILLER_14_210 ();
 DECAPx4_ASAP7_75t_R FILLER_14_226 ();
 FILLER_ASAP7_75t_R FILLER_14_236 ();
 DECAPx2_ASAP7_75t_R FILLER_14_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_250 ();
 DECAPx6_ASAP7_75t_R FILLER_14_257 ();
 DECAPx10_ASAP7_75t_R FILLER_14_277 ();
 DECAPx1_ASAP7_75t_R FILLER_14_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_303 ();
 DECAPx1_ASAP7_75t_R FILLER_14_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_314 ();
 DECAPx4_ASAP7_75t_R FILLER_14_321 ();
 FILLER_ASAP7_75t_R FILLER_14_331 ();
 DECAPx10_ASAP7_75t_R FILLER_14_336 ();
 DECAPx2_ASAP7_75t_R FILLER_14_358 ();
 FILLER_ASAP7_75t_R FILLER_14_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_387 ();
 DECAPx2_ASAP7_75t_R FILLER_14_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_432 ();
 DECAPx4_ASAP7_75t_R FILLER_14_450 ();
 FILLER_ASAP7_75t_R FILLER_14_460 ();
 DECAPx2_ASAP7_75t_R FILLER_14_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_487 ();
 DECAPx4_ASAP7_75t_R FILLER_14_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_519 ();
 DECAPx4_ASAP7_75t_R FILLER_14_536 ();
 FILLER_ASAP7_75t_R FILLER_14_546 ();
 FILLER_ASAP7_75t_R FILLER_14_558 ();
 DECAPx1_ASAP7_75t_R FILLER_14_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_582 ();
 DECAPx4_ASAP7_75t_R FILLER_14_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_621 ();
 DECAPx2_ASAP7_75t_R FILLER_14_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_638 ();
 DECAPx6_ASAP7_75t_R FILLER_14_646 ();
 FILLER_ASAP7_75t_R FILLER_14_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_662 ();
 DECAPx1_ASAP7_75t_R FILLER_14_747 ();
 DECAPx1_ASAP7_75t_R FILLER_14_772 ();
 DECAPx4_ASAP7_75t_R FILLER_14_797 ();
 FILLER_ASAP7_75t_R FILLER_14_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_829 ();
 FILLER_ASAP7_75t_R FILLER_14_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_848 ();
 DECAPx2_ASAP7_75t_R FILLER_14_870 ();
 FILLER_ASAP7_75t_R FILLER_14_876 ();
 DECAPx4_ASAP7_75t_R FILLER_14_893 ();
 FILLER_ASAP7_75t_R FILLER_14_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_905 ();
 FILLER_ASAP7_75t_R FILLER_14_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_939 ();
 DECAPx4_ASAP7_75t_R FILLER_14_957 ();
 FILLER_ASAP7_75t_R FILLER_14_967 ();
 DECAPx10_ASAP7_75t_R FILLER_14_979 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_14_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1079 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1109 ();
 FILLER_ASAP7_75t_R FILLER_14_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1143 ();
 FILLER_ASAP7_75t_R FILLER_14_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1269 ();
 FILLER_ASAP7_75t_R FILLER_14_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_15_68 ();
 DECAPx6_ASAP7_75t_R FILLER_15_90 ();
 DECAPx1_ASAP7_75t_R FILLER_15_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_157 ();
 DECAPx1_ASAP7_75t_R FILLER_15_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_174 ();
 FILLER_ASAP7_75t_R FILLER_15_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_201 ();
 FILLER_ASAP7_75t_R FILLER_15_223 ();
 DECAPx4_ASAP7_75t_R FILLER_15_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_274 ();
 DECAPx1_ASAP7_75t_R FILLER_15_284 ();
 FILLER_ASAP7_75t_R FILLER_15_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_302 ();
 DECAPx1_ASAP7_75t_R FILLER_15_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_313 ();
 DECAPx1_ASAP7_75t_R FILLER_15_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_337 ();
 DECAPx10_ASAP7_75t_R FILLER_15_345 ();
 DECAPx2_ASAP7_75t_R FILLER_15_367 ();
 DECAPx10_ASAP7_75t_R FILLER_15_408 ();
 DECAPx10_ASAP7_75t_R FILLER_15_458 ();
 DECAPx1_ASAP7_75t_R FILLER_15_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_484 ();
 DECAPx10_ASAP7_75t_R FILLER_15_488 ();
 DECAPx4_ASAP7_75t_R FILLER_15_510 ();
 FILLER_ASAP7_75t_R FILLER_15_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_527 ();
 DECAPx6_ASAP7_75t_R FILLER_15_545 ();
 DECAPx1_ASAP7_75t_R FILLER_15_559 ();
 DECAPx4_ASAP7_75t_R FILLER_15_584 ();
 FILLER_ASAP7_75t_R FILLER_15_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_602 ();
 DECAPx2_ASAP7_75t_R FILLER_15_609 ();
 DECAPx10_ASAP7_75t_R FILLER_15_636 ();
 DECAPx6_ASAP7_75t_R FILLER_15_658 ();
 DECAPx2_ASAP7_75t_R FILLER_15_672 ();
 DECAPx2_ASAP7_75t_R FILLER_15_690 ();
 DECAPx6_ASAP7_75t_R FILLER_15_702 ();
 FILLER_ASAP7_75t_R FILLER_15_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_718 ();
 DECAPx6_ASAP7_75t_R FILLER_15_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_757 ();
 DECAPx4_ASAP7_75t_R FILLER_15_768 ();
 DECAPx2_ASAP7_75t_R FILLER_15_792 ();
 FILLER_ASAP7_75t_R FILLER_15_798 ();
 FILLER_ASAP7_75t_R FILLER_15_849 ();
 DECAPx1_ASAP7_75t_R FILLER_15_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_865 ();
 FILLER_ASAP7_75t_R FILLER_15_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_901 ();
 DECAPx4_ASAP7_75t_R FILLER_15_950 ();
 FILLER_ASAP7_75t_R FILLER_15_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_986 ();
 FILLER_ASAP7_75t_R FILLER_15_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1061 ();
 FILLER_ASAP7_75t_R FILLER_15_1067 ();
 FILLER_ASAP7_75t_R FILLER_15_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_15_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1214 ();
 FILLER_ASAP7_75t_R FILLER_15_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1285 ();
 FILLER_ASAP7_75t_R FILLER_15_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_16_68 ();
 DECAPx4_ASAP7_75t_R FILLER_16_90 ();
 FILLER_ASAP7_75t_R FILLER_16_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_152 ();
 DECAPx2_ASAP7_75t_R FILLER_16_196 ();
 DECAPx2_ASAP7_75t_R FILLER_16_218 ();
 FILLER_ASAP7_75t_R FILLER_16_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_243 ();
 FILLER_ASAP7_75t_R FILLER_16_284 ();
 FILLER_ASAP7_75t_R FILLER_16_296 ();
 FILLER_ASAP7_75t_R FILLER_16_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_307 ();
 FILLER_ASAP7_75t_R FILLER_16_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_317 ();
 FILLER_ASAP7_75t_R FILLER_16_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_326 ();
 FILLER_ASAP7_75t_R FILLER_16_353 ();
 DECAPx10_ASAP7_75t_R FILLER_16_361 ();
 DECAPx2_ASAP7_75t_R FILLER_16_383 ();
 DECAPx4_ASAP7_75t_R FILLER_16_431 ();
 DECAPx4_ASAP7_75t_R FILLER_16_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_474 ();
 DECAPx6_ASAP7_75t_R FILLER_16_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_517 ();
 DECAPx6_ASAP7_75t_R FILLER_16_528 ();
 DECAPx1_ASAP7_75t_R FILLER_16_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_546 ();
 DECAPx6_ASAP7_75t_R FILLER_16_554 ();
 FILLER_ASAP7_75t_R FILLER_16_568 ();
 DECAPx10_ASAP7_75t_R FILLER_16_627 ();
 DECAPx10_ASAP7_75t_R FILLER_16_649 ();
 DECAPx1_ASAP7_75t_R FILLER_16_671 ();
 DECAPx10_ASAP7_75t_R FILLER_16_696 ();
 DECAPx10_ASAP7_75t_R FILLER_16_718 ();
 DECAPx6_ASAP7_75t_R FILLER_16_740 ();
 FILLER_ASAP7_75t_R FILLER_16_754 ();
 FILLER_ASAP7_75t_R FILLER_16_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_768 ();
 DECAPx2_ASAP7_75t_R FILLER_16_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_806 ();
 DECAPx6_ASAP7_75t_R FILLER_16_814 ();
 DECAPx1_ASAP7_75t_R FILLER_16_828 ();
 DECAPx10_ASAP7_75t_R FILLER_16_839 ();
 DECAPx1_ASAP7_75t_R FILLER_16_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_865 ();
 DECAPx4_ASAP7_75t_R FILLER_16_881 ();
 DECAPx2_ASAP7_75t_R FILLER_16_894 ();
 FILLER_ASAP7_75t_R FILLER_16_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_902 ();
 DECAPx2_ASAP7_75t_R FILLER_16_915 ();
 FILLER_ASAP7_75t_R FILLER_16_921 ();
 DECAPx4_ASAP7_75t_R FILLER_16_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_945 ();
 DECAPx4_ASAP7_75t_R FILLER_16_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_16_1129 ();
 FILLER_ASAP7_75t_R FILLER_16_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1152 ();
 FILLER_ASAP7_75t_R FILLER_16_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1183 ();
 FILLER_ASAP7_75t_R FILLER_16_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_16_1216 ();
 FILLER_ASAP7_75t_R FILLER_16_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1228 ();
 FILLER_ASAP7_75t_R FILLER_16_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_16_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_17_68 ();
 DECAPx6_ASAP7_75t_R FILLER_17_90 ();
 DECAPx2_ASAP7_75t_R FILLER_17_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_110 ();
 FILLER_ASAP7_75t_R FILLER_17_117 ();
 FILLER_ASAP7_75t_R FILLER_17_126 ();
 DECAPx1_ASAP7_75t_R FILLER_17_131 ();
 FILLER_ASAP7_75t_R FILLER_17_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_149 ();
 DECAPx1_ASAP7_75t_R FILLER_17_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_167 ();
 DECAPx6_ASAP7_75t_R FILLER_17_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_208 ();
 DECAPx2_ASAP7_75t_R FILLER_17_216 ();
 FILLER_ASAP7_75t_R FILLER_17_222 ();
 DECAPx2_ASAP7_75t_R FILLER_17_265 ();
 FILLER_ASAP7_75t_R FILLER_17_278 ();
 DECAPx1_ASAP7_75t_R FILLER_17_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_305 ();
 DECAPx2_ASAP7_75t_R FILLER_17_312 ();
 FILLER_ASAP7_75t_R FILLER_17_333 ();
 DECAPx10_ASAP7_75t_R FILLER_17_341 ();
 DECAPx1_ASAP7_75t_R FILLER_17_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_367 ();
 DECAPx2_ASAP7_75t_R FILLER_17_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_381 ();
 DECAPx4_ASAP7_75t_R FILLER_17_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_409 ();
 DECAPx2_ASAP7_75t_R FILLER_17_417 ();
 FILLER_ASAP7_75t_R FILLER_17_423 ();
 FILLER_ASAP7_75t_R FILLER_17_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_437 ();
 DECAPx2_ASAP7_75t_R FILLER_17_445 ();
 DECAPx2_ASAP7_75t_R FILLER_17_461 ();
 DECAPx1_ASAP7_75t_R FILLER_17_488 ();
 DECAPx1_ASAP7_75t_R FILLER_17_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_604 ();
 FILLER_ASAP7_75t_R FILLER_17_615 ();
 FILLER_ASAP7_75t_R FILLER_17_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_653 ();
 DECAPx2_ASAP7_75t_R FILLER_17_672 ();
 FILLER_ASAP7_75t_R FILLER_17_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_687 ();
 DECAPx6_ASAP7_75t_R FILLER_17_700 ();
 DECAPx2_ASAP7_75t_R FILLER_17_714 ();
 DECAPx10_ASAP7_75t_R FILLER_17_726 ();
 DECAPx4_ASAP7_75t_R FILLER_17_748 ();
 DECAPx10_ASAP7_75t_R FILLER_17_786 ();
 DECAPx10_ASAP7_75t_R FILLER_17_808 ();
 DECAPx2_ASAP7_75t_R FILLER_17_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_864 ();
 DECAPx2_ASAP7_75t_R FILLER_17_873 ();
 FILLER_ASAP7_75t_R FILLER_17_879 ();
 DECAPx6_ASAP7_75t_R FILLER_17_899 ();
 DECAPx1_ASAP7_75t_R FILLER_17_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_917 ();
 FILLER_ASAP7_75t_R FILLER_17_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_928 ();
 DECAPx2_ASAP7_75t_R FILLER_17_941 ();
 FILLER_ASAP7_75t_R FILLER_17_947 ();
 DECAPx6_ASAP7_75t_R FILLER_17_952 ();
 FILLER_ASAP7_75t_R FILLER_17_966 ();
 FILLER_ASAP7_75t_R FILLER_17_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_999 ();
 FILLER_ASAP7_75t_R FILLER_17_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_17_1097 ();
 FILLER_ASAP7_75t_R FILLER_17_1113 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_17_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_18_90 ();
 DECAPx2_ASAP7_75t_R FILLER_18_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_118 ();
 DECAPx10_ASAP7_75t_R FILLER_18_125 ();
 DECAPx1_ASAP7_75t_R FILLER_18_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_151 ();
 FILLER_ASAP7_75t_R FILLER_18_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_160 ();
 FILLER_ASAP7_75t_R FILLER_18_167 ();
 FILLER_ASAP7_75t_R FILLER_18_172 ();
 DECAPx1_ASAP7_75t_R FILLER_18_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_182 ();
 DECAPx10_ASAP7_75t_R FILLER_18_213 ();
 DECAPx10_ASAP7_75t_R FILLER_18_235 ();
 DECAPx6_ASAP7_75t_R FILLER_18_263 ();
 DECAPx2_ASAP7_75t_R FILLER_18_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_283 ();
 DECAPx1_ASAP7_75t_R FILLER_18_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_308 ();
 DECAPx2_ASAP7_75t_R FILLER_18_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_331 ();
 DECAPx10_ASAP7_75t_R FILLER_18_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_368 ();
 FILLER_ASAP7_75t_R FILLER_18_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_392 ();
 DECAPx4_ASAP7_75t_R FILLER_18_403 ();
 FILLER_ASAP7_75t_R FILLER_18_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_415 ();
 DECAPx1_ASAP7_75t_R FILLER_18_458 ();
 FILLER_ASAP7_75t_R FILLER_18_464 ();
 DECAPx4_ASAP7_75t_R FILLER_18_473 ();
 DECAPx2_ASAP7_75t_R FILLER_18_525 ();
 DECAPx2_ASAP7_75t_R FILLER_18_562 ();
 FILLER_ASAP7_75t_R FILLER_18_568 ();
 DECAPx2_ASAP7_75t_R FILLER_18_596 ();
 FILLER_ASAP7_75t_R FILLER_18_602 ();
 DECAPx1_ASAP7_75t_R FILLER_18_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_618 ();
 FILLER_ASAP7_75t_R FILLER_18_640 ();
 DECAPx6_ASAP7_75t_R FILLER_18_663 ();
 DECAPx2_ASAP7_75t_R FILLER_18_677 ();
 DECAPx10_ASAP7_75t_R FILLER_18_689 ();
 DECAPx1_ASAP7_75t_R FILLER_18_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_715 ();
 FILLER_ASAP7_75t_R FILLER_18_737 ();
 DECAPx10_ASAP7_75t_R FILLER_18_760 ();
 DECAPx4_ASAP7_75t_R FILLER_18_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_864 ();
 FILLER_ASAP7_75t_R FILLER_18_881 ();
 FILLER_ASAP7_75t_R FILLER_18_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_906 ();
 FILLER_ASAP7_75t_R FILLER_18_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_959 ();
 DECAPx2_ASAP7_75t_R FILLER_18_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_976 ();
 FILLER_ASAP7_75t_R FILLER_18_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_991 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_18_1094 ();
 FILLER_ASAP7_75t_R FILLER_18_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_18_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1158 ();
 DECAPx4_ASAP7_75t_R FILLER_18_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1216 ();
 FILLER_ASAP7_75t_R FILLER_18_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1269 ();
 FILLER_ASAP7_75t_R FILLER_18_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_19_68 ();
 DECAPx10_ASAP7_75t_R FILLER_19_90 ();
 DECAPx1_ASAP7_75t_R FILLER_19_112 ();
 DECAPx2_ASAP7_75t_R FILLER_19_132 ();
 DECAPx10_ASAP7_75t_R FILLER_19_144 ();
 DECAPx2_ASAP7_75t_R FILLER_19_166 ();
 FILLER_ASAP7_75t_R FILLER_19_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_174 ();
 FILLER_ASAP7_75t_R FILLER_19_193 ();
 FILLER_ASAP7_75t_R FILLER_19_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_215 ();
 DECAPx2_ASAP7_75t_R FILLER_19_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_236 ();
 DECAPx2_ASAP7_75t_R FILLER_19_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_250 ();
 DECAPx2_ASAP7_75t_R FILLER_19_265 ();
 FILLER_ASAP7_75t_R FILLER_19_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_279 ();
 DECAPx2_ASAP7_75t_R FILLER_19_286 ();
 DECAPx1_ASAP7_75t_R FILLER_19_310 ();
 DECAPx4_ASAP7_75t_R FILLER_19_321 ();
 FILLER_ASAP7_75t_R FILLER_19_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_333 ();
 FILLER_ASAP7_75t_R FILLER_19_354 ();
 DECAPx2_ASAP7_75t_R FILLER_19_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_386 ();
 DECAPx2_ASAP7_75t_R FILLER_19_408 ();
 FILLER_ASAP7_75t_R FILLER_19_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_416 ();
 DECAPx2_ASAP7_75t_R FILLER_19_434 ();
 FILLER_ASAP7_75t_R FILLER_19_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_442 ();
 DECAPx6_ASAP7_75t_R FILLER_19_453 ();
 DECAPx6_ASAP7_75t_R FILLER_19_477 ();
 FILLER_ASAP7_75t_R FILLER_19_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_493 ();
 FILLER_ASAP7_75t_R FILLER_19_501 ();
 FILLER_ASAP7_75t_R FILLER_19_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_518 ();
 DECAPx10_ASAP7_75t_R FILLER_19_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_551 ();
 DECAPx2_ASAP7_75t_R FILLER_19_558 ();
 FILLER_ASAP7_75t_R FILLER_19_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_576 ();
 DECAPx2_ASAP7_75t_R FILLER_19_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_590 ();
 DECAPx1_ASAP7_75t_R FILLER_19_597 ();
 DECAPx4_ASAP7_75t_R FILLER_19_608 ();
 FILLER_ASAP7_75t_R FILLER_19_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_620 ();
 DECAPx10_ASAP7_75t_R FILLER_19_631 ();
 FILLER_ASAP7_75t_R FILLER_19_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_655 ();
 DECAPx6_ASAP7_75t_R FILLER_19_668 ();
 DECAPx1_ASAP7_75t_R FILLER_19_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_686 ();
 FILLER_ASAP7_75t_R FILLER_19_720 ();
 DECAPx2_ASAP7_75t_R FILLER_19_739 ();
 FILLER_ASAP7_75t_R FILLER_19_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_747 ();
 DECAPx6_ASAP7_75t_R FILLER_19_792 ();
 FILLER_ASAP7_75t_R FILLER_19_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_808 ();
 FILLER_ASAP7_75t_R FILLER_19_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_833 ();
 FILLER_ASAP7_75t_R FILLER_19_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_911 ();
 DECAPx10_ASAP7_75t_R FILLER_19_926 ();
 FILLER_ASAP7_75t_R FILLER_19_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_950 ();
 DECAPx1_ASAP7_75t_R FILLER_19_977 ();
 DECAPx1_ASAP7_75t_R FILLER_19_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_19_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1108 ();
 FILLER_ASAP7_75t_R FILLER_19_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1179 ();
 FILLER_ASAP7_75t_R FILLER_19_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_20_90 ();
 FILLER_ASAP7_75t_R FILLER_20_140 ();
 DECAPx1_ASAP7_75t_R FILLER_20_161 ();
 DECAPx1_ASAP7_75t_R FILLER_20_178 ();
 DECAPx10_ASAP7_75t_R FILLER_20_186 ();
 FILLER_ASAP7_75t_R FILLER_20_254 ();
 FILLER_ASAP7_75t_R FILLER_20_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_266 ();
 FILLER_ASAP7_75t_R FILLER_20_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_275 ();
 FILLER_ASAP7_75t_R FILLER_20_286 ();
 DECAPx2_ASAP7_75t_R FILLER_20_304 ();
 FILLER_ASAP7_75t_R FILLER_20_310 ();
 DECAPx2_ASAP7_75t_R FILLER_20_321 ();
 DECAPx2_ASAP7_75t_R FILLER_20_335 ();
 FILLER_ASAP7_75t_R FILLER_20_341 ();
 DECAPx1_ASAP7_75t_R FILLER_20_381 ();
 DECAPx1_ASAP7_75t_R FILLER_20_392 ();
 DECAPx1_ASAP7_75t_R FILLER_20_406 ();
 DECAPx10_ASAP7_75t_R FILLER_20_427 ();
 DECAPx4_ASAP7_75t_R FILLER_20_449 ();
 FILLER_ASAP7_75t_R FILLER_20_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_461 ();
 DECAPx10_ASAP7_75t_R FILLER_20_464 ();
 DECAPx4_ASAP7_75t_R FILLER_20_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_506 ();
 DECAPx6_ASAP7_75t_R FILLER_20_514 ();
 FILLER_ASAP7_75t_R FILLER_20_528 ();
 DECAPx2_ASAP7_75t_R FILLER_20_540 ();
 FILLER_ASAP7_75t_R FILLER_20_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_548 ();
 DECAPx4_ASAP7_75t_R FILLER_20_566 ();
 DECAPx1_ASAP7_75t_R FILLER_20_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_601 ();
 DECAPx6_ASAP7_75t_R FILLER_20_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_637 ();
 DECAPx6_ASAP7_75t_R FILLER_20_645 ();
 DECAPx1_ASAP7_75t_R FILLER_20_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_663 ();
 DECAPx10_ASAP7_75t_R FILLER_20_671 ();
 DECAPx10_ASAP7_75t_R FILLER_20_693 ();
 DECAPx10_ASAP7_75t_R FILLER_20_715 ();
 DECAPx2_ASAP7_75t_R FILLER_20_737 ();
 FILLER_ASAP7_75t_R FILLER_20_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_745 ();
 DECAPx4_ASAP7_75t_R FILLER_20_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_787 ();
 FILLER_ASAP7_75t_R FILLER_20_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_797 ();
 DECAPx2_ASAP7_75t_R FILLER_20_806 ();
 FILLER_ASAP7_75t_R FILLER_20_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_814 ();
 FILLER_ASAP7_75t_R FILLER_20_832 ();
 FILLER_ASAP7_75t_R FILLER_20_841 ();
 FILLER_ASAP7_75t_R FILLER_20_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_866 ();
 DECAPx4_ASAP7_75t_R FILLER_20_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_889 ();
 FILLER_ASAP7_75t_R FILLER_20_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_912 ();
 FILLER_ASAP7_75t_R FILLER_20_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_918 ();
 DECAPx2_ASAP7_75t_R FILLER_20_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_967 ();
 DECAPx1_ASAP7_75t_R FILLER_20_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_982 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_20_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_20_1196 ();
 FILLER_ASAP7_75t_R FILLER_20_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1269 ();
 FILLER_ASAP7_75t_R FILLER_20_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_21_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_146 ();
 FILLER_ASAP7_75t_R FILLER_21_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_193 ();
 DECAPx1_ASAP7_75t_R FILLER_21_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_210 ();
 FILLER_ASAP7_75t_R FILLER_21_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_226 ();
 FILLER_ASAP7_75t_R FILLER_21_239 ();
 FILLER_ASAP7_75t_R FILLER_21_247 ();
 FILLER_ASAP7_75t_R FILLER_21_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_310 ();
 FILLER_ASAP7_75t_R FILLER_21_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_320 ();
 DECAPx10_ASAP7_75t_R FILLER_21_329 ();
 DECAPx6_ASAP7_75t_R FILLER_21_351 ();
 DECAPx2_ASAP7_75t_R FILLER_21_365 ();
 DECAPx2_ASAP7_75t_R FILLER_21_397 ();
 FILLER_ASAP7_75t_R FILLER_21_403 ();
 DECAPx4_ASAP7_75t_R FILLER_21_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_436 ();
 DECAPx4_ASAP7_75t_R FILLER_21_454 ();
 DECAPx1_ASAP7_75t_R FILLER_21_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_502 ();
 DECAPx1_ASAP7_75t_R FILLER_21_513 ();
 DECAPx2_ASAP7_75t_R FILLER_21_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_550 ();
 DECAPx4_ASAP7_75t_R FILLER_21_579 ();
 FILLER_ASAP7_75t_R FILLER_21_589 ();
 DECAPx10_ASAP7_75t_R FILLER_21_597 ();
 FILLER_ASAP7_75t_R FILLER_21_619 ();
 DECAPx4_ASAP7_75t_R FILLER_21_629 ();
 FILLER_ASAP7_75t_R FILLER_21_639 ();
 DECAPx10_ASAP7_75t_R FILLER_21_662 ();
 DECAPx10_ASAP7_75t_R FILLER_21_684 ();
 DECAPx10_ASAP7_75t_R FILLER_21_706 ();
 DECAPx1_ASAP7_75t_R FILLER_21_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_732 ();
 FILLER_ASAP7_75t_R FILLER_21_743 ();
 DECAPx6_ASAP7_75t_R FILLER_21_773 ();
 DECAPx2_ASAP7_75t_R FILLER_21_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_793 ();
 DECAPx6_ASAP7_75t_R FILLER_21_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_815 ();
 DECAPx6_ASAP7_75t_R FILLER_21_872 ();
 DECAPx2_ASAP7_75t_R FILLER_21_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_892 ();
 DECAPx6_ASAP7_75t_R FILLER_21_903 ();
 DECAPx1_ASAP7_75t_R FILLER_21_917 ();
 DECAPx2_ASAP7_75t_R FILLER_21_926 ();
 FILLER_ASAP7_75t_R FILLER_21_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_934 ();
 DECAPx4_ASAP7_75t_R FILLER_21_942 ();
 FILLER_ASAP7_75t_R FILLER_21_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_954 ();
 FILLER_ASAP7_75t_R FILLER_21_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_21_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_21_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_21_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_21_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1127 ();
 FILLER_ASAP7_75t_R FILLER_21_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_21_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_21_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1268 ();
 FILLER_ASAP7_75t_R FILLER_21_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx6_ASAP7_75t_R FILLER_22_112 ();
 DECAPx2_ASAP7_75t_R FILLER_22_126 ();
 DECAPx4_ASAP7_75t_R FILLER_22_139 ();
 DECAPx2_ASAP7_75t_R FILLER_22_155 ();
 FILLER_ASAP7_75t_R FILLER_22_161 ();
 DECAPx2_ASAP7_75t_R FILLER_22_175 ();
 DECAPx10_ASAP7_75t_R FILLER_22_193 ();
 DECAPx6_ASAP7_75t_R FILLER_22_215 ();
 DECAPx10_ASAP7_75t_R FILLER_22_241 ();
 DECAPx10_ASAP7_75t_R FILLER_22_263 ();
 DECAPx1_ASAP7_75t_R FILLER_22_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_289 ();
 FILLER_ASAP7_75t_R FILLER_22_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_313 ();
 DECAPx1_ASAP7_75t_R FILLER_22_321 ();
 DECAPx10_ASAP7_75t_R FILLER_22_331 ();
 DECAPx1_ASAP7_75t_R FILLER_22_353 ();
 FILLER_ASAP7_75t_R FILLER_22_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_377 ();
 DECAPx6_ASAP7_75t_R FILLER_22_395 ();
 DECAPx2_ASAP7_75t_R FILLER_22_409 ();
 DECAPx1_ASAP7_75t_R FILLER_22_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_461 ();
 DECAPx10_ASAP7_75t_R FILLER_22_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_529 ();
 DECAPx2_ASAP7_75t_R FILLER_22_561 ();
 FILLER_ASAP7_75t_R FILLER_22_567 ();
 DECAPx1_ASAP7_75t_R FILLER_22_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_594 ();
 FILLER_ASAP7_75t_R FILLER_22_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_618 ();
 FILLER_ASAP7_75t_R FILLER_22_641 ();
 DECAPx6_ASAP7_75t_R FILLER_22_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_667 ();
 FILLER_ASAP7_75t_R FILLER_22_675 ();
 DECAPx10_ASAP7_75t_R FILLER_22_689 ();
 DECAPx2_ASAP7_75t_R FILLER_22_711 ();
 FILLER_ASAP7_75t_R FILLER_22_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_719 ();
 DECAPx1_ASAP7_75t_R FILLER_22_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_730 ();
 DECAPx4_ASAP7_75t_R FILLER_22_738 ();
 FILLER_ASAP7_75t_R FILLER_22_748 ();
 DECAPx6_ASAP7_75t_R FILLER_22_771 ();
 DECAPx4_ASAP7_75t_R FILLER_22_814 ();
 FILLER_ASAP7_75t_R FILLER_22_824 ();
 DECAPx10_ASAP7_75t_R FILLER_22_840 ();
 DECAPx6_ASAP7_75t_R FILLER_22_865 ();
 DECAPx2_ASAP7_75t_R FILLER_22_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_885 ();
 DECAPx4_ASAP7_75t_R FILLER_22_898 ();
 FILLER_ASAP7_75t_R FILLER_22_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_910 ();
 DECAPx1_ASAP7_75t_R FILLER_22_932 ();
 DECAPx2_ASAP7_75t_R FILLER_22_946 ();
 FILLER_ASAP7_75t_R FILLER_22_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_954 ();
 FILLER_ASAP7_75t_R FILLER_22_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_997 ();
 FILLER_ASAP7_75t_R FILLER_22_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1080 ();
 FILLER_ASAP7_75t_R FILLER_22_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1131 ();
 FILLER_ASAP7_75t_R FILLER_22_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1151 ();
 FILLER_ASAP7_75t_R FILLER_22_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1171 ();
 FILLER_ASAP7_75t_R FILLER_22_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1202 ();
 FILLER_ASAP7_75t_R FILLER_22_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_23_68 ();
 DECAPx6_ASAP7_75t_R FILLER_23_90 ();
 DECAPx1_ASAP7_75t_R FILLER_23_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_108 ();
 DECAPx2_ASAP7_75t_R FILLER_23_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_143 ();
 DECAPx1_ASAP7_75t_R FILLER_23_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_167 ();
 DECAPx2_ASAP7_75t_R FILLER_23_175 ();
 FILLER_ASAP7_75t_R FILLER_23_181 ();
 FILLER_ASAP7_75t_R FILLER_23_188 ();
 FILLER_ASAP7_75t_R FILLER_23_212 ();
 FILLER_ASAP7_75t_R FILLER_23_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_230 ();
 DECAPx4_ASAP7_75t_R FILLER_23_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_248 ();
 FILLER_ASAP7_75t_R FILLER_23_281 ();
 DECAPx2_ASAP7_75t_R FILLER_23_299 ();
 DECAPx6_ASAP7_75t_R FILLER_23_320 ();
 DECAPx1_ASAP7_75t_R FILLER_23_413 ();
 DECAPx4_ASAP7_75t_R FILLER_23_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_454 ();
 DECAPx10_ASAP7_75t_R FILLER_23_461 ();
 DECAPx4_ASAP7_75t_R FILLER_23_483 ();
 FILLER_ASAP7_75t_R FILLER_23_493 ();
 DECAPx10_ASAP7_75t_R FILLER_23_541 ();
 DECAPx2_ASAP7_75t_R FILLER_23_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_569 ();
 FILLER_ASAP7_75t_R FILLER_23_580 ();
 DECAPx2_ASAP7_75t_R FILLER_23_603 ();
 DECAPx2_ASAP7_75t_R FILLER_23_621 ();
 DECAPx10_ASAP7_75t_R FILLER_23_649 ();
 DECAPx4_ASAP7_75t_R FILLER_23_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_681 ();
 DECAPx2_ASAP7_75t_R FILLER_23_698 ();
 FILLER_ASAP7_75t_R FILLER_23_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_713 ();
 FILLER_ASAP7_75t_R FILLER_23_749 ();
 DECAPx1_ASAP7_75t_R FILLER_23_768 ();
 FILLER_ASAP7_75t_R FILLER_23_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_789 ();
 DECAPx2_ASAP7_75t_R FILLER_23_804 ();
 FILLER_ASAP7_75t_R FILLER_23_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_818 ();
 DECAPx4_ASAP7_75t_R FILLER_23_836 ();
 FILLER_ASAP7_75t_R FILLER_23_846 ();
 DECAPx6_ASAP7_75t_R FILLER_23_855 ();
 DECAPx1_ASAP7_75t_R FILLER_23_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_885 ();
 FILLER_ASAP7_75t_R FILLER_23_922 ();
 FILLER_ASAP7_75t_R FILLER_23_935 ();
 DECAPx1_ASAP7_75t_R FILLER_23_958 ();
 DECAPx2_ASAP7_75t_R FILLER_23_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_23_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1072 ();
 FILLER_ASAP7_75t_R FILLER_23_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_23_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1200 ();
 DECAPx6_ASAP7_75t_R FILLER_23_1222 ();
 FILLER_ASAP7_75t_R FILLER_23_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_23_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx2_ASAP7_75t_R FILLER_24_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_118 ();
 FILLER_ASAP7_75t_R FILLER_24_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_166 ();
 FILLER_ASAP7_75t_R FILLER_24_189 ();
 DECAPx6_ASAP7_75t_R FILLER_24_219 ();
 DECAPx2_ASAP7_75t_R FILLER_24_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_247 ();
 FILLER_ASAP7_75t_R FILLER_24_260 ();
 DECAPx2_ASAP7_75t_R FILLER_24_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_288 ();
 DECAPx6_ASAP7_75t_R FILLER_24_297 ();
 FILLER_ASAP7_75t_R FILLER_24_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_313 ();
 DECAPx10_ASAP7_75t_R FILLER_24_320 ();
 DECAPx10_ASAP7_75t_R FILLER_24_342 ();
 DECAPx2_ASAP7_75t_R FILLER_24_364 ();
 FILLER_ASAP7_75t_R FILLER_24_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_372 ();
 DECAPx10_ASAP7_75t_R FILLER_24_387 ();
 DECAPx2_ASAP7_75t_R FILLER_24_409 ();
 FILLER_ASAP7_75t_R FILLER_24_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_435 ();
 DECAPx1_ASAP7_75t_R FILLER_24_458 ();
 DECAPx2_ASAP7_75t_R FILLER_24_472 ();
 FILLER_ASAP7_75t_R FILLER_24_478 ();
 DECAPx4_ASAP7_75t_R FILLER_24_512 ();
 DECAPx10_ASAP7_75t_R FILLER_24_532 ();
 DECAPx4_ASAP7_75t_R FILLER_24_575 ();
 FILLER_ASAP7_75t_R FILLER_24_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_587 ();
 DECAPx10_ASAP7_75t_R FILLER_24_600 ();
 DECAPx10_ASAP7_75t_R FILLER_24_622 ();
 DECAPx10_ASAP7_75t_R FILLER_24_644 ();
 DECAPx10_ASAP7_75t_R FILLER_24_666 ();
 DECAPx6_ASAP7_75t_R FILLER_24_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_702 ();
 DECAPx4_ASAP7_75t_R FILLER_24_724 ();
 FILLER_ASAP7_75t_R FILLER_24_734 ();
 DECAPx6_ASAP7_75t_R FILLER_24_748 ();
 FILLER_ASAP7_75t_R FILLER_24_762 ();
 DECAPx10_ASAP7_75t_R FILLER_24_791 ();
 DECAPx6_ASAP7_75t_R FILLER_24_813 ();
 FILLER_ASAP7_75t_R FILLER_24_827 ();
 DECAPx2_ASAP7_75t_R FILLER_24_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_901 ();
 DECAPx2_ASAP7_75t_R FILLER_24_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_918 ();
 DECAPx4_ASAP7_75t_R FILLER_24_925 ();
 FILLER_ASAP7_75t_R FILLER_24_935 ();
 DECAPx10_ASAP7_75t_R FILLER_24_947 ();
 DECAPx2_ASAP7_75t_R FILLER_24_969 ();
 FILLER_ASAP7_75t_R FILLER_24_975 ();
 FILLER_ASAP7_75t_R FILLER_24_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_985 ();
 DECAPx4_ASAP7_75t_R FILLER_24_996 ();
 DECAPx6_ASAP7_75t_R FILLER_24_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1063 ();
 FILLER_ASAP7_75t_R FILLER_24_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1094 ();
 FILLER_ASAP7_75t_R FILLER_24_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_24_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1169 ();
 FILLER_ASAP7_75t_R FILLER_24_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_24_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_25_90 ();
 FILLER_ASAP7_75t_R FILLER_25_112 ();
 DECAPx4_ASAP7_75t_R FILLER_25_145 ();
 DECAPx1_ASAP7_75t_R FILLER_25_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_168 ();
 DECAPx10_ASAP7_75t_R FILLER_25_184 ();
 DECAPx4_ASAP7_75t_R FILLER_25_206 ();
 DECAPx6_ASAP7_75t_R FILLER_25_224 ();
 FILLER_ASAP7_75t_R FILLER_25_238 ();
 DECAPx1_ASAP7_75t_R FILLER_25_252 ();
 DECAPx2_ASAP7_75t_R FILLER_25_275 ();
 FILLER_ASAP7_75t_R FILLER_25_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_283 ();
 FILLER_ASAP7_75t_R FILLER_25_307 ();
 DECAPx4_ASAP7_75t_R FILLER_25_339 ();
 FILLER_ASAP7_75t_R FILLER_25_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_351 ();
 FILLER_ASAP7_75t_R FILLER_25_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_376 ();
 DECAPx4_ASAP7_75t_R FILLER_25_398 ();
 DECAPx6_ASAP7_75t_R FILLER_25_429 ();
 FILLER_ASAP7_75t_R FILLER_25_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_445 ();
 FILLER_ASAP7_75t_R FILLER_25_458 ();
 DECAPx10_ASAP7_75t_R FILLER_25_466 ();
 DECAPx2_ASAP7_75t_R FILLER_25_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_494 ();
 DECAPx10_ASAP7_75t_R FILLER_25_517 ();
 DECAPx6_ASAP7_75t_R FILLER_25_539 ();
 DECAPx1_ASAP7_75t_R FILLER_25_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_557 ();
 DECAPx10_ASAP7_75t_R FILLER_25_561 ();
 DECAPx10_ASAP7_75t_R FILLER_25_583 ();
 DECAPx10_ASAP7_75t_R FILLER_25_605 ();
 DECAPx10_ASAP7_75t_R FILLER_25_627 ();
 DECAPx6_ASAP7_75t_R FILLER_25_649 ();
 DECAPx1_ASAP7_75t_R FILLER_25_663 ();
 DECAPx6_ASAP7_75t_R FILLER_25_673 ();
 FILLER_ASAP7_75t_R FILLER_25_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_689 ();
 DECAPx10_ASAP7_75t_R FILLER_25_711 ();
 DECAPx4_ASAP7_75t_R FILLER_25_733 ();
 FILLER_ASAP7_75t_R FILLER_25_743 ();
 DECAPx1_ASAP7_75t_R FILLER_25_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_770 ();
 DECAPx1_ASAP7_75t_R FILLER_25_792 ();
 FILLER_ASAP7_75t_R FILLER_25_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_828 ();
 DECAPx2_ASAP7_75t_R FILLER_25_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_859 ();
 DECAPx10_ASAP7_75t_R FILLER_25_873 ();
 DECAPx1_ASAP7_75t_R FILLER_25_895 ();
 DECAPx6_ASAP7_75t_R FILLER_25_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_923 ();
 DECAPx1_ASAP7_75t_R FILLER_25_926 ();
 DECAPx4_ASAP7_75t_R FILLER_25_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_968 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1005 ();
 FILLER_ASAP7_75t_R FILLER_25_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1041 ();
 FILLER_ASAP7_75t_R FILLER_25_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1068 ();
 FILLER_ASAP7_75t_R FILLER_25_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1102 ();
 FILLER_ASAP7_75t_R FILLER_25_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1137 ();
 FILLER_ASAP7_75t_R FILLER_25_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_25_1163 ();
 FILLER_ASAP7_75t_R FILLER_25_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1203 ();
 FILLER_ASAP7_75t_R FILLER_25_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 DECAPx6_ASAP7_75t_R FILLER_26_112 ();
 DECAPx2_ASAP7_75t_R FILLER_26_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_132 ();
 DECAPx10_ASAP7_75t_R FILLER_26_140 ();
 DECAPx10_ASAP7_75t_R FILLER_26_162 ();
 DECAPx10_ASAP7_75t_R FILLER_26_184 ();
 DECAPx4_ASAP7_75t_R FILLER_26_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_216 ();
 FILLER_ASAP7_75t_R FILLER_26_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_238 ();
 DECAPx6_ASAP7_75t_R FILLER_26_274 ();
 DECAPx1_ASAP7_75t_R FILLER_26_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_310 ();
 DECAPx10_ASAP7_75t_R FILLER_26_333 ();
 DECAPx10_ASAP7_75t_R FILLER_26_355 ();
 DECAPx1_ASAP7_75t_R FILLER_26_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_381 ();
 DECAPx6_ASAP7_75t_R FILLER_26_399 ();
 FILLER_ASAP7_75t_R FILLER_26_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_415 ();
 DECAPx2_ASAP7_75t_R FILLER_26_419 ();
 FILLER_ASAP7_75t_R FILLER_26_425 ();
 FILLER_ASAP7_75t_R FILLER_26_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_439 ();
 DECAPx4_ASAP7_75t_R FILLER_26_450 ();
 FILLER_ASAP7_75t_R FILLER_26_460 ();
 DECAPx6_ASAP7_75t_R FILLER_26_464 ();
 FILLER_ASAP7_75t_R FILLER_26_478 ();
 DECAPx1_ASAP7_75t_R FILLER_26_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_498 ();
 DECAPx10_ASAP7_75t_R FILLER_26_513 ();
 DECAPx1_ASAP7_75t_R FILLER_26_535 ();
 DECAPx10_ASAP7_75t_R FILLER_26_566 ();
 DECAPx4_ASAP7_75t_R FILLER_26_588 ();
 FILLER_ASAP7_75t_R FILLER_26_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_600 ();
 DECAPx10_ASAP7_75t_R FILLER_26_609 ();
 DECAPx1_ASAP7_75t_R FILLER_26_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_635 ();
 DECAPx6_ASAP7_75t_R FILLER_26_642 ();
 DECAPx1_ASAP7_75t_R FILLER_26_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_660 ();
 DECAPx10_ASAP7_75t_R FILLER_26_669 ();
 DECAPx2_ASAP7_75t_R FILLER_26_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_704 ();
 DECAPx10_ASAP7_75t_R FILLER_26_717 ();
 DECAPx1_ASAP7_75t_R FILLER_26_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_770 ();
 DECAPx10_ASAP7_75t_R FILLER_26_792 ();
 DECAPx4_ASAP7_75t_R FILLER_26_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_861 ();
 DECAPx1_ASAP7_75t_R FILLER_26_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_880 ();
 DECAPx2_ASAP7_75t_R FILLER_26_893 ();
 FILLER_ASAP7_75t_R FILLER_26_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_901 ();
 DECAPx4_ASAP7_75t_R FILLER_26_935 ();
 FILLER_ASAP7_75t_R FILLER_26_945 ();
 DECAPx4_ASAP7_75t_R FILLER_26_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_979 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1098 ();
 FILLER_ASAP7_75t_R FILLER_26_1172 ();
 FILLER_ASAP7_75t_R FILLER_26_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1245 ();
 FILLER_ASAP7_75t_R FILLER_26_1267 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_27_90 ();
 DECAPx10_ASAP7_75t_R FILLER_27_112 ();
 DECAPx10_ASAP7_75t_R FILLER_27_134 ();
 DECAPx6_ASAP7_75t_R FILLER_27_156 ();
 DECAPx2_ASAP7_75t_R FILLER_27_170 ();
 FILLER_ASAP7_75t_R FILLER_27_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_189 ();
 DECAPx2_ASAP7_75t_R FILLER_27_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_214 ();
 FILLER_ASAP7_75t_R FILLER_27_227 ();
 DECAPx1_ASAP7_75t_R FILLER_27_236 ();
 FILLER_ASAP7_75t_R FILLER_27_247 ();
 FILLER_ASAP7_75t_R FILLER_27_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_260 ();
 DECAPx2_ASAP7_75t_R FILLER_27_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_274 ();
 FILLER_ASAP7_75t_R FILLER_27_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_306 ();
 FILLER_ASAP7_75t_R FILLER_27_322 ();
 DECAPx4_ASAP7_75t_R FILLER_27_332 ();
 FILLER_ASAP7_75t_R FILLER_27_342 ();
 DECAPx10_ASAP7_75t_R FILLER_27_386 ();
 DECAPx4_ASAP7_75t_R FILLER_27_408 ();
 FILLER_ASAP7_75t_R FILLER_27_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_426 ();
 DECAPx2_ASAP7_75t_R FILLER_27_434 ();
 FILLER_ASAP7_75t_R FILLER_27_440 ();
 DECAPx2_ASAP7_75t_R FILLER_27_454 ();
 DECAPx10_ASAP7_75t_R FILLER_27_466 ();
 DECAPx2_ASAP7_75t_R FILLER_27_488 ();
 DECAPx10_ASAP7_75t_R FILLER_27_512 ();
 DECAPx1_ASAP7_75t_R FILLER_27_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_538 ();
 DECAPx6_ASAP7_75t_R FILLER_27_555 ();
 DECAPx2_ASAP7_75t_R FILLER_27_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_575 ();
 DECAPx2_ASAP7_75t_R FILLER_27_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_600 ();
 DECAPx10_ASAP7_75t_R FILLER_27_607 ();
 DECAPx10_ASAP7_75t_R FILLER_27_629 ();
 DECAPx1_ASAP7_75t_R FILLER_27_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_655 ();
 DECAPx4_ASAP7_75t_R FILLER_27_662 ();
 FILLER_ASAP7_75t_R FILLER_27_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_674 ();
 DECAPx4_ASAP7_75t_R FILLER_27_681 ();
 DECAPx4_ASAP7_75t_R FILLER_27_718 ();
 DECAPx2_ASAP7_75t_R FILLER_27_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_744 ();
 DECAPx10_ASAP7_75t_R FILLER_27_784 ();
 DECAPx4_ASAP7_75t_R FILLER_27_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_816 ();
 DECAPx1_ASAP7_75t_R FILLER_27_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_827 ();
 DECAPx2_ASAP7_75t_R FILLER_27_844 ();
 DECAPx2_ASAP7_75t_R FILLER_27_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_878 ();
 FILLER_ASAP7_75t_R FILLER_27_903 ();
 FILLER_ASAP7_75t_R FILLER_27_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_923 ();
 DECAPx10_ASAP7_75t_R FILLER_27_926 ();
 DECAPx10_ASAP7_75t_R FILLER_27_948 ();
 DECAPx4_ASAP7_75t_R FILLER_27_970 ();
 DECAPx1_ASAP7_75t_R FILLER_27_996 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1096 ();
 FILLER_ASAP7_75t_R FILLER_27_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1165 ();
 FILLER_ASAP7_75t_R FILLER_27_1175 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1207 ();
 FILLER_ASAP7_75t_R FILLER_27_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1226 ();
 FILLER_ASAP7_75t_R FILLER_27_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_27_1277 ();
 FILLER_ASAP7_75t_R FILLER_27_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_28_68 ();
 DECAPx10_ASAP7_75t_R FILLER_28_90 ();
 DECAPx6_ASAP7_75t_R FILLER_28_130 ();
 FILLER_ASAP7_75t_R FILLER_28_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_146 ();
 FILLER_ASAP7_75t_R FILLER_28_178 ();
 FILLER_ASAP7_75t_R FILLER_28_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_197 ();
 FILLER_ASAP7_75t_R FILLER_28_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_248 ();
 FILLER_ASAP7_75t_R FILLER_28_256 ();
 DECAPx2_ASAP7_75t_R FILLER_28_266 ();
 DECAPx2_ASAP7_75t_R FILLER_28_279 ();
 FILLER_ASAP7_75t_R FILLER_28_285 ();
 DECAPx10_ASAP7_75t_R FILLER_28_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_351 ();
 FILLER_ASAP7_75t_R FILLER_28_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_359 ();
 DECAPx6_ASAP7_75t_R FILLER_28_366 ();
 DECAPx4_ASAP7_75t_R FILLER_28_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_408 ();
 DECAPx6_ASAP7_75t_R FILLER_28_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_461 ();
 DECAPx2_ASAP7_75t_R FILLER_28_470 ();
 DECAPx2_ASAP7_75t_R FILLER_28_498 ();
 FILLER_ASAP7_75t_R FILLER_28_504 ();
 DECAPx1_ASAP7_75t_R FILLER_28_524 ();
 DECAPx2_ASAP7_75t_R FILLER_28_546 ();
 DECAPx10_ASAP7_75t_R FILLER_28_566 ();
 DECAPx4_ASAP7_75t_R FILLER_28_588 ();
 DECAPx10_ASAP7_75t_R FILLER_28_606 ();
 DECAPx10_ASAP7_75t_R FILLER_28_628 ();
 DECAPx10_ASAP7_75t_R FILLER_28_650 ();
 DECAPx4_ASAP7_75t_R FILLER_28_672 ();
 DECAPx10_ASAP7_75t_R FILLER_28_703 ();
 DECAPx6_ASAP7_75t_R FILLER_28_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_739 ();
 DECAPx6_ASAP7_75t_R FILLER_28_746 ();
 FILLER_ASAP7_75t_R FILLER_28_760 ();
 DECAPx1_ASAP7_75t_R FILLER_28_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_834 ();
 DECAPx10_ASAP7_75t_R FILLER_28_845 ();
 DECAPx10_ASAP7_75t_R FILLER_28_867 ();
 DECAPx6_ASAP7_75t_R FILLER_28_889 ();
 DECAPx1_ASAP7_75t_R FILLER_28_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_907 ();
 DECAPx4_ASAP7_75t_R FILLER_28_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_939 ();
 DECAPx6_ASAP7_75t_R FILLER_28_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_975 ();
 FILLER_ASAP7_75t_R FILLER_28_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_28_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1104 ();
 FILLER_ASAP7_75t_R FILLER_28_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_28_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_28_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_29_68 ();
 DECAPx6_ASAP7_75t_R FILLER_29_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_155 ();
 FILLER_ASAP7_75t_R FILLER_29_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_193 ();
 DECAPx1_ASAP7_75t_R FILLER_29_227 ();
 DECAPx2_ASAP7_75t_R FILLER_29_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_253 ();
 DECAPx4_ASAP7_75t_R FILLER_29_277 ();
 FILLER_ASAP7_75t_R FILLER_29_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_313 ();
 DECAPx10_ASAP7_75t_R FILLER_29_330 ();
 DECAPx1_ASAP7_75t_R FILLER_29_352 ();
 DECAPx4_ASAP7_75t_R FILLER_29_366 ();
 DECAPx4_ASAP7_75t_R FILLER_29_397 ();
 DECAPx1_ASAP7_75t_R FILLER_29_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_423 ();
 DECAPx6_ASAP7_75t_R FILLER_29_430 ();
 DECAPx1_ASAP7_75t_R FILLER_29_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_448 ();
 FILLER_ASAP7_75t_R FILLER_29_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_483 ();
 DECAPx2_ASAP7_75t_R FILLER_29_490 ();
 DECAPx6_ASAP7_75t_R FILLER_29_512 ();
 FILLER_ASAP7_75t_R FILLER_29_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_534 ();
 DECAPx10_ASAP7_75t_R FILLER_29_542 ();
 DECAPx10_ASAP7_75t_R FILLER_29_564 ();
 DECAPx4_ASAP7_75t_R FILLER_29_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_596 ();
 DECAPx10_ASAP7_75t_R FILLER_29_612 ();
 DECAPx10_ASAP7_75t_R FILLER_29_652 ();
 DECAPx4_ASAP7_75t_R FILLER_29_674 ();
 FILLER_ASAP7_75t_R FILLER_29_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_686 ();
 DECAPx10_ASAP7_75t_R FILLER_29_690 ();
 DECAPx10_ASAP7_75t_R FILLER_29_712 ();
 DECAPx6_ASAP7_75t_R FILLER_29_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_748 ();
 FILLER_ASAP7_75t_R FILLER_29_770 ();
 DECAPx4_ASAP7_75t_R FILLER_29_779 ();
 DECAPx4_ASAP7_75t_R FILLER_29_834 ();
 FILLER_ASAP7_75t_R FILLER_29_844 ();
 DECAPx2_ASAP7_75t_R FILLER_29_866 ();
 DECAPx6_ASAP7_75t_R FILLER_29_905 ();
 DECAPx1_ASAP7_75t_R FILLER_29_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_923 ();
 DECAPx2_ASAP7_75t_R FILLER_29_926 ();
 FILLER_ASAP7_75t_R FILLER_29_932 ();
 DECAPx4_ASAP7_75t_R FILLER_29_951 ();
 FILLER_ASAP7_75t_R FILLER_29_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_999 ();
 DECAPx4_ASAP7_75t_R FILLER_29_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1040 ();
 FILLER_ASAP7_75t_R FILLER_29_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1177 ();
 FILLER_ASAP7_75t_R FILLER_29_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_29_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1241 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_30_68 ();
 DECAPx6_ASAP7_75t_R FILLER_30_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_153 ();
 DECAPx2_ASAP7_75t_R FILLER_30_166 ();
 FILLER_ASAP7_75t_R FILLER_30_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_184 ();
 DECAPx1_ASAP7_75t_R FILLER_30_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_201 ();
 DECAPx2_ASAP7_75t_R FILLER_30_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_217 ();
 DECAPx4_ASAP7_75t_R FILLER_30_235 ();
 FILLER_ASAP7_75t_R FILLER_30_245 ();
 DECAPx10_ASAP7_75t_R FILLER_30_259 ();
 DECAPx4_ASAP7_75t_R FILLER_30_281 ();
 DECAPx4_ASAP7_75t_R FILLER_30_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_313 ();
 DECAPx10_ASAP7_75t_R FILLER_30_320 ();
 DECAPx2_ASAP7_75t_R FILLER_30_342 ();
 FILLER_ASAP7_75t_R FILLER_30_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_350 ();
 DECAPx1_ASAP7_75t_R FILLER_30_357 ();
 DECAPx4_ASAP7_75t_R FILLER_30_368 ();
 FILLER_ASAP7_75t_R FILLER_30_378 ();
 DECAPx6_ASAP7_75t_R FILLER_30_390 ();
 DECAPx1_ASAP7_75t_R FILLER_30_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_408 ();
 DECAPx2_ASAP7_75t_R FILLER_30_447 ();
 FILLER_ASAP7_75t_R FILLER_30_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_455 ();
 FILLER_ASAP7_75t_R FILLER_30_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_483 ();
 DECAPx10_ASAP7_75t_R FILLER_30_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_521 ();
 DECAPx1_ASAP7_75t_R FILLER_30_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_535 ();
 DECAPx1_ASAP7_75t_R FILLER_30_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_566 ();
 DECAPx6_ASAP7_75t_R FILLER_30_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_599 ();
 DECAPx6_ASAP7_75t_R FILLER_30_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_624 ();
 FILLER_ASAP7_75t_R FILLER_30_628 ();
 DECAPx1_ASAP7_75t_R FILLER_30_652 ();
 DECAPx10_ASAP7_75t_R FILLER_30_678 ();
 DECAPx10_ASAP7_75t_R FILLER_30_700 ();
 DECAPx10_ASAP7_75t_R FILLER_30_722 ();
 DECAPx10_ASAP7_75t_R FILLER_30_744 ();
 DECAPx10_ASAP7_75t_R FILLER_30_778 ();
 FILLER_ASAP7_75t_R FILLER_30_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_802 ();
 FILLER_ASAP7_75t_R FILLER_30_824 ();
 DECAPx2_ASAP7_75t_R FILLER_30_840 ();
 FILLER_ASAP7_75t_R FILLER_30_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_877 ();
 DECAPx6_ASAP7_75t_R FILLER_30_893 ();
 DECAPx1_ASAP7_75t_R FILLER_30_907 ();
 DECAPx4_ASAP7_75t_R FILLER_30_924 ();
 FILLER_ASAP7_75t_R FILLER_30_934 ();
 FILLER_ASAP7_75t_R FILLER_30_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_955 ();
 FILLER_ASAP7_75t_R FILLER_30_987 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1013 ();
 FILLER_ASAP7_75t_R FILLER_30_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_30_1035 ();
 FILLER_ASAP7_75t_R FILLER_30_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1047 ();
 FILLER_ASAP7_75t_R FILLER_30_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_30_1133 ();
 FILLER_ASAP7_75t_R FILLER_30_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1192 ();
 FILLER_ASAP7_75t_R FILLER_30_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1223 ();
 FILLER_ASAP7_75t_R FILLER_30_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_31_68 ();
 DECAPx10_ASAP7_75t_R FILLER_31_90 ();
 DECAPx4_ASAP7_75t_R FILLER_31_112 ();
 FILLER_ASAP7_75t_R FILLER_31_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_124 ();
 DECAPx2_ASAP7_75t_R FILLER_31_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_149 ();
 DECAPx2_ASAP7_75t_R FILLER_31_159 ();
 DECAPx2_ASAP7_75t_R FILLER_31_174 ();
 FILLER_ASAP7_75t_R FILLER_31_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_196 ();
 FILLER_ASAP7_75t_R FILLER_31_206 ();
 DECAPx1_ASAP7_75t_R FILLER_31_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_225 ();
 DECAPx4_ASAP7_75t_R FILLER_31_234 ();
 FILLER_ASAP7_75t_R FILLER_31_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_246 ();
 DECAPx6_ASAP7_75t_R FILLER_31_265 ();
 DECAPx1_ASAP7_75t_R FILLER_31_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_283 ();
 DECAPx6_ASAP7_75t_R FILLER_31_290 ();
 DECAPx4_ASAP7_75t_R FILLER_31_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_328 ();
 FILLER_ASAP7_75t_R FILLER_31_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_362 ();
 DECAPx2_ASAP7_75t_R FILLER_31_399 ();
 DECAPx2_ASAP7_75t_R FILLER_31_421 ();
 FILLER_ASAP7_75t_R FILLER_31_427 ();
 DECAPx2_ASAP7_75t_R FILLER_31_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_441 ();
 FILLER_ASAP7_75t_R FILLER_31_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_491 ();
 DECAPx2_ASAP7_75t_R FILLER_31_498 ();
 FILLER_ASAP7_75t_R FILLER_31_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_506 ();
 DECAPx10_ASAP7_75t_R FILLER_31_535 ();
 DECAPx1_ASAP7_75t_R FILLER_31_557 ();
 DECAPx4_ASAP7_75t_R FILLER_31_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_591 ();
 FILLER_ASAP7_75t_R FILLER_31_598 ();
 FILLER_ASAP7_75t_R FILLER_31_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_609 ();
 FILLER_ASAP7_75t_R FILLER_31_618 ();
 DECAPx4_ASAP7_75t_R FILLER_31_628 ();
 FILLER_ASAP7_75t_R FILLER_31_638 ();
 DECAPx6_ASAP7_75t_R FILLER_31_646 ();
 FILLER_ASAP7_75t_R FILLER_31_660 ();
 DECAPx6_ASAP7_75t_R FILLER_31_672 ();
 DECAPx2_ASAP7_75t_R FILLER_31_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_692 ();
 DECAPx2_ASAP7_75t_R FILLER_31_708 ();
 FILLER_ASAP7_75t_R FILLER_31_714 ();
 DECAPx4_ASAP7_75t_R FILLER_31_726 ();
 FILLER_ASAP7_75t_R FILLER_31_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_738 ();
 DECAPx6_ASAP7_75t_R FILLER_31_746 ();
 FILLER_ASAP7_75t_R FILLER_31_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_762 ();
 DECAPx10_ASAP7_75t_R FILLER_31_769 ();
 DECAPx10_ASAP7_75t_R FILLER_31_791 ();
 DECAPx2_ASAP7_75t_R FILLER_31_813 ();
 FILLER_ASAP7_75t_R FILLER_31_825 ();
 DECAPx1_ASAP7_75t_R FILLER_31_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_837 ();
 DECAPx2_ASAP7_75t_R FILLER_31_845 ();
 FILLER_ASAP7_75t_R FILLER_31_851 ();
 DECAPx1_ASAP7_75t_R FILLER_31_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_885 ();
 FILLER_ASAP7_75t_R FILLER_31_898 ();
 DECAPx1_ASAP7_75t_R FILLER_31_926 ();
 DECAPx1_ASAP7_75t_R FILLER_31_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_946 ();
 DECAPx6_ASAP7_75t_R FILLER_31_968 ();
 FILLER_ASAP7_75t_R FILLER_31_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_987 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1075 ();
 FILLER_ASAP7_75t_R FILLER_31_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1093 ();
 FILLER_ASAP7_75t_R FILLER_31_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1122 ();
 FILLER_ASAP7_75t_R FILLER_31_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1207 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1225 ();
 FILLER_ASAP7_75t_R FILLER_31_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1248 ();
 DECAPx6_ASAP7_75t_R FILLER_31_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_32_68 ();
 DECAPx10_ASAP7_75t_R FILLER_32_90 ();
 DECAPx1_ASAP7_75t_R FILLER_32_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_141 ();
 DECAPx10_ASAP7_75t_R FILLER_32_154 ();
 DECAPx1_ASAP7_75t_R FILLER_32_176 ();
 DECAPx1_ASAP7_75t_R FILLER_32_200 ();
 FILLER_ASAP7_75t_R FILLER_32_211 ();
 DECAPx1_ASAP7_75t_R FILLER_32_220 ();
 FILLER_ASAP7_75t_R FILLER_32_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_258 ();
 DECAPx10_ASAP7_75t_R FILLER_32_288 ();
 DECAPx10_ASAP7_75t_R FILLER_32_310 ();
 FILLER_ASAP7_75t_R FILLER_32_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_334 ();
 DECAPx10_ASAP7_75t_R FILLER_32_363 ();
 DECAPx6_ASAP7_75t_R FILLER_32_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_416 ();
 DECAPx2_ASAP7_75t_R FILLER_32_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_433 ();
 FILLER_ASAP7_75t_R FILLER_32_441 ();
 DECAPx1_ASAP7_75t_R FILLER_32_458 ();
 FILLER_ASAP7_75t_R FILLER_32_464 ();
 DECAPx4_ASAP7_75t_R FILLER_32_475 ();
 FILLER_ASAP7_75t_R FILLER_32_485 ();
 DECAPx4_ASAP7_75t_R FILLER_32_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_506 ();
 DECAPx4_ASAP7_75t_R FILLER_32_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_553 ();
 DECAPx6_ASAP7_75t_R FILLER_32_563 ();
 DECAPx2_ASAP7_75t_R FILLER_32_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_589 ();
 DECAPx1_ASAP7_75t_R FILLER_32_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_606 ();
 DECAPx10_ASAP7_75t_R FILLER_32_628 ();
 DECAPx2_ASAP7_75t_R FILLER_32_650 ();
 FILLER_ASAP7_75t_R FILLER_32_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_658 ();
 DECAPx4_ASAP7_75t_R FILLER_32_680 ();
 DECAPx10_ASAP7_75t_R FILLER_32_706 ();
 DECAPx10_ASAP7_75t_R FILLER_32_728 ();
 DECAPx4_ASAP7_75t_R FILLER_32_750 ();
 FILLER_ASAP7_75t_R FILLER_32_760 ();
 DECAPx10_ASAP7_75t_R FILLER_32_778 ();
 DECAPx10_ASAP7_75t_R FILLER_32_800 ();
 DECAPx6_ASAP7_75t_R FILLER_32_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_836 ();
 DECAPx2_ASAP7_75t_R FILLER_32_864 ();
 FILLER_ASAP7_75t_R FILLER_32_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_872 ();
 DECAPx4_ASAP7_75t_R FILLER_32_877 ();
 DECAPx10_ASAP7_75t_R FILLER_32_945 ();
 DECAPx10_ASAP7_75t_R FILLER_32_967 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1045 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1067 ();
 FILLER_ASAP7_75t_R FILLER_32_1088 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1167 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_33_68 ();
 DECAPx10_ASAP7_75t_R FILLER_33_90 ();
 DECAPx1_ASAP7_75t_R FILLER_33_112 ();
 FILLER_ASAP7_75t_R FILLER_33_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_131 ();
 DECAPx4_ASAP7_75t_R FILLER_33_139 ();
 FILLER_ASAP7_75t_R FILLER_33_149 ();
 DECAPx4_ASAP7_75t_R FILLER_33_158 ();
 DECAPx1_ASAP7_75t_R FILLER_33_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_178 ();
 FILLER_ASAP7_75t_R FILLER_33_185 ();
 DECAPx6_ASAP7_75t_R FILLER_33_204 ();
 DECAPx2_ASAP7_75t_R FILLER_33_218 ();
 DECAPx2_ASAP7_75t_R FILLER_33_244 ();
 FILLER_ASAP7_75t_R FILLER_33_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_252 ();
 FILLER_ASAP7_75t_R FILLER_33_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_299 ();
 DECAPx10_ASAP7_75t_R FILLER_33_316 ();
 FILLER_ASAP7_75t_R FILLER_33_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_365 ();
 DECAPx10_ASAP7_75t_R FILLER_33_386 ();
 FILLER_ASAP7_75t_R FILLER_33_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_410 ();
 DECAPx6_ASAP7_75t_R FILLER_33_429 ();
 DECAPx2_ASAP7_75t_R FILLER_33_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_449 ();
 DECAPx4_ASAP7_75t_R FILLER_33_456 ();
 DECAPx2_ASAP7_75t_R FILLER_33_475 ();
 FILLER_ASAP7_75t_R FILLER_33_481 ();
 DECAPx10_ASAP7_75t_R FILLER_33_489 ();
 DECAPx2_ASAP7_75t_R FILLER_33_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_517 ();
 DECAPx6_ASAP7_75t_R FILLER_33_534 ();
 DECAPx1_ASAP7_75t_R FILLER_33_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_552 ();
 DECAPx6_ASAP7_75t_R FILLER_33_561 ();
 DECAPx1_ASAP7_75t_R FILLER_33_575 ();
 DECAPx4_ASAP7_75t_R FILLER_33_591 ();
 DECAPx1_ASAP7_75t_R FILLER_33_609 ();
 DECAPx6_ASAP7_75t_R FILLER_33_627 ();
 DECAPx4_ASAP7_75t_R FILLER_33_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_657 ();
 DECAPx4_ASAP7_75t_R FILLER_33_668 ();
 DECAPx6_ASAP7_75t_R FILLER_33_684 ();
 DECAPx2_ASAP7_75t_R FILLER_33_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_704 ();
 DECAPx2_ASAP7_75t_R FILLER_33_711 ();
 DECAPx2_ASAP7_75t_R FILLER_33_729 ();
 DECAPx6_ASAP7_75t_R FILLER_33_741 ();
 FILLER_ASAP7_75t_R FILLER_33_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_757 ();
 DECAPx6_ASAP7_75t_R FILLER_33_764 ();
 DECAPx1_ASAP7_75t_R FILLER_33_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_798 ();
 DECAPx10_ASAP7_75t_R FILLER_33_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_830 ();
 DECAPx10_ASAP7_75t_R FILLER_33_841 ();
 DECAPx2_ASAP7_75t_R FILLER_33_863 ();
 FILLER_ASAP7_75t_R FILLER_33_869 ();
 DECAPx10_ASAP7_75t_R FILLER_33_877 ();
 DECAPx1_ASAP7_75t_R FILLER_33_899 ();
 DECAPx4_ASAP7_75t_R FILLER_33_926 ();
 FILLER_ASAP7_75t_R FILLER_33_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_938 ();
 DECAPx1_ASAP7_75t_R FILLER_33_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_964 ();
 DECAPx1_ASAP7_75t_R FILLER_33_995 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1080 ();
 FILLER_ASAP7_75t_R FILLER_33_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1164 ();
 FILLER_ASAP7_75t_R FILLER_33_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_34_68 ();
 DECAPx10_ASAP7_75t_R FILLER_34_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_112 ();
 DECAPx1_ASAP7_75t_R FILLER_34_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_130 ();
 DECAPx4_ASAP7_75t_R FILLER_34_161 ();
 FILLER_ASAP7_75t_R FILLER_34_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_173 ();
 FILLER_ASAP7_75t_R FILLER_34_192 ();
 DECAPx10_ASAP7_75t_R FILLER_34_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_249 ();
 DECAPx2_ASAP7_75t_R FILLER_34_256 ();
 FILLER_ASAP7_75t_R FILLER_34_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_300 ();
 DECAPx1_ASAP7_75t_R FILLER_34_322 ();
 DECAPx6_ASAP7_75t_R FILLER_34_334 ();
 FILLER_ASAP7_75t_R FILLER_34_348 ();
 DECAPx1_ASAP7_75t_R FILLER_34_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_372 ();
 FILLER_ASAP7_75t_R FILLER_34_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_403 ();
 DECAPx2_ASAP7_75t_R FILLER_34_428 ();
 DECAPx2_ASAP7_75t_R FILLER_34_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_447 ();
 FILLER_ASAP7_75t_R FILLER_34_454 ();
 FILLER_ASAP7_75t_R FILLER_34_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_466 ();
 DECAPx1_ASAP7_75t_R FILLER_34_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_481 ();
 DECAPx2_ASAP7_75t_R FILLER_34_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_529 ();
 DECAPx2_ASAP7_75t_R FILLER_34_536 ();
 FILLER_ASAP7_75t_R FILLER_34_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_544 ();
 DECAPx2_ASAP7_75t_R FILLER_34_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_563 ();
 DECAPx4_ASAP7_75t_R FILLER_34_573 ();
 FILLER_ASAP7_75t_R FILLER_34_583 ();
 FILLER_ASAP7_75t_R FILLER_34_591 ();
 DECAPx6_ASAP7_75t_R FILLER_34_605 ();
 DECAPx1_ASAP7_75t_R FILLER_34_619 ();
 DECAPx10_ASAP7_75t_R FILLER_34_641 ();
 DECAPx2_ASAP7_75t_R FILLER_34_663 ();
 FILLER_ASAP7_75t_R FILLER_34_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_671 ();
 DECAPx10_ASAP7_75t_R FILLER_34_691 ();
 DECAPx10_ASAP7_75t_R FILLER_34_713 ();
 DECAPx10_ASAP7_75t_R FILLER_34_735 ();
 DECAPx10_ASAP7_75t_R FILLER_34_757 ();
 DECAPx10_ASAP7_75t_R FILLER_34_779 ();
 DECAPx1_ASAP7_75t_R FILLER_34_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_805 ();
 FILLER_ASAP7_75t_R FILLER_34_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_831 ();
 DECAPx6_ASAP7_75t_R FILLER_34_839 ();
 FILLER_ASAP7_75t_R FILLER_34_853 ();
 DECAPx2_ASAP7_75t_R FILLER_34_900 ();
 FILLER_ASAP7_75t_R FILLER_34_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_908 ();
 DECAPx10_ASAP7_75t_R FILLER_34_930 ();
 DECAPx1_ASAP7_75t_R FILLER_34_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_971 ();
 DECAPx1_ASAP7_75t_R FILLER_34_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1025 ();
 FILLER_ASAP7_75t_R FILLER_34_1047 ();
 FILLER_ASAP7_75t_R FILLER_34_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1088 ();
 FILLER_ASAP7_75t_R FILLER_34_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1107 ();
 FILLER_ASAP7_75t_R FILLER_34_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1194 ();
 FILLER_ASAP7_75t_R FILLER_34_1209 ();
 FILLER_ASAP7_75t_R FILLER_34_1243 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1268 ();
 FILLER_ASAP7_75t_R FILLER_34_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_35_68 ();
 DECAPx2_ASAP7_75t_R FILLER_35_90 ();
 FILLER_ASAP7_75t_R FILLER_35_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_98 ();
 DECAPx2_ASAP7_75t_R FILLER_35_113 ();
 FILLER_ASAP7_75t_R FILLER_35_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_121 ();
 FILLER_ASAP7_75t_R FILLER_35_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_164 ();
 FILLER_ASAP7_75t_R FILLER_35_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_181 ();
 FILLER_ASAP7_75t_R FILLER_35_189 ();
 DECAPx2_ASAP7_75t_R FILLER_35_200 ();
 FILLER_ASAP7_75t_R FILLER_35_217 ();
 DECAPx2_ASAP7_75t_R FILLER_35_228 ();
 FILLER_ASAP7_75t_R FILLER_35_234 ();
 DECAPx1_ASAP7_75t_R FILLER_35_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_246 ();
 DECAPx2_ASAP7_75t_R FILLER_35_253 ();
 FILLER_ASAP7_75t_R FILLER_35_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_261 ();
 DECAPx1_ASAP7_75t_R FILLER_35_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_311 ();
 DECAPx4_ASAP7_75t_R FILLER_35_321 ();
 DECAPx2_ASAP7_75t_R FILLER_35_340 ();
 DECAPx1_ASAP7_75t_R FILLER_35_352 ();
 FILLER_ASAP7_75t_R FILLER_35_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_365 ();
 FILLER_ASAP7_75t_R FILLER_35_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_382 ();
 DECAPx1_ASAP7_75t_R FILLER_35_403 ();
 DECAPx2_ASAP7_75t_R FILLER_35_425 ();
 FILLER_ASAP7_75t_R FILLER_35_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_463 ();
 FILLER_ASAP7_75t_R FILLER_35_480 ();
 DECAPx1_ASAP7_75t_R FILLER_35_494 ();
 DECAPx2_ASAP7_75t_R FILLER_35_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_514 ();
 DECAPx4_ASAP7_75t_R FILLER_35_533 ();
 FILLER_ASAP7_75t_R FILLER_35_553 ();
 DECAPx1_ASAP7_75t_R FILLER_35_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_592 ();
 DECAPx6_ASAP7_75t_R FILLER_35_606 ();
 FILLER_ASAP7_75t_R FILLER_35_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_622 ();
 DECAPx6_ASAP7_75t_R FILLER_35_632 ();
 DECAPx1_ASAP7_75t_R FILLER_35_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_650 ();
 DECAPx10_ASAP7_75t_R FILLER_35_669 ();
 DECAPx4_ASAP7_75t_R FILLER_35_691 ();
 FILLER_ASAP7_75t_R FILLER_35_701 ();
 DECAPx10_ASAP7_75t_R FILLER_35_709 ();
 DECAPx10_ASAP7_75t_R FILLER_35_731 ();
 DECAPx10_ASAP7_75t_R FILLER_35_753 ();
 FILLER_ASAP7_75t_R FILLER_35_775 ();
 DECAPx10_ASAP7_75t_R FILLER_35_783 ();
 DECAPx6_ASAP7_75t_R FILLER_35_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_819 ();
 DECAPx2_ASAP7_75t_R FILLER_35_827 ();
 DECAPx2_ASAP7_75t_R FILLER_35_854 ();
 FILLER_ASAP7_75t_R FILLER_35_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_862 ();
 DECAPx1_ASAP7_75t_R FILLER_35_885 ();
 DECAPx2_ASAP7_75t_R FILLER_35_896 ();
 FILLER_ASAP7_75t_R FILLER_35_902 ();
 FILLER_ASAP7_75t_R FILLER_35_916 ();
 FILLER_ASAP7_75t_R FILLER_35_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_942 ();
 DECAPx10_ASAP7_75t_R FILLER_35_970 ();
 DECAPx10_ASAP7_75t_R FILLER_35_992 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1089 ();
 FILLER_ASAP7_75t_R FILLER_35_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1107 ();
 FILLER_ASAP7_75t_R FILLER_35_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1184 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1220 ();
 FILLER_ASAP7_75t_R FILLER_35_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1268 ();
 FILLER_ASAP7_75t_R FILLER_35_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_36_68 ();
 DECAPx4_ASAP7_75t_R FILLER_36_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_100 ();
 FILLER_ASAP7_75t_R FILLER_36_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_146 ();
 FILLER_ASAP7_75t_R FILLER_36_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_226 ();
 DECAPx2_ASAP7_75t_R FILLER_36_243 ();
 FILLER_ASAP7_75t_R FILLER_36_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_284 ();
 DECAPx6_ASAP7_75t_R FILLER_36_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_315 ();
 DECAPx2_ASAP7_75t_R FILLER_36_342 ();
 FILLER_ASAP7_75t_R FILLER_36_355 ();
 FILLER_ASAP7_75t_R FILLER_36_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_374 ();
 DECAPx10_ASAP7_75t_R FILLER_36_392 ();
 DECAPx2_ASAP7_75t_R FILLER_36_414 ();
 DECAPx6_ASAP7_75t_R FILLER_36_427 ();
 DECAPx1_ASAP7_75t_R FILLER_36_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_445 ();
 FILLER_ASAP7_75t_R FILLER_36_460 ();
 DECAPx2_ASAP7_75t_R FILLER_36_464 ();
 FILLER_ASAP7_75t_R FILLER_36_470 ();
 DECAPx2_ASAP7_75t_R FILLER_36_492 ();
 DECAPx2_ASAP7_75t_R FILLER_36_522 ();
 DECAPx2_ASAP7_75t_R FILLER_36_538 ();
 FILLER_ASAP7_75t_R FILLER_36_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_561 ();
 DECAPx1_ASAP7_75t_R FILLER_36_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_582 ();
 DECAPx10_ASAP7_75t_R FILLER_36_603 ();
 DECAPx1_ASAP7_75t_R FILLER_36_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_629 ();
 DECAPx2_ASAP7_75t_R FILLER_36_645 ();
 FILLER_ASAP7_75t_R FILLER_36_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_653 ();
 DECAPx10_ASAP7_75t_R FILLER_36_672 ();
 DECAPx2_ASAP7_75t_R FILLER_36_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_716 ();
 DECAPx10_ASAP7_75t_R FILLER_36_740 ();
 DECAPx1_ASAP7_75t_R FILLER_36_762 ();
 DECAPx10_ASAP7_75t_R FILLER_36_788 ();
 DECAPx4_ASAP7_75t_R FILLER_36_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_820 ();
 DECAPx4_ASAP7_75t_R FILLER_36_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_852 ();
 FILLER_ASAP7_75t_R FILLER_36_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_871 ();
 FILLER_ASAP7_75t_R FILLER_36_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_880 ();
 FILLER_ASAP7_75t_R FILLER_36_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_901 ();
 DECAPx6_ASAP7_75t_R FILLER_36_912 ();
 FILLER_ASAP7_75t_R FILLER_36_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_928 ();
 DECAPx10_ASAP7_75t_R FILLER_36_935 ();
 DECAPx6_ASAP7_75t_R FILLER_36_957 ();
 FILLER_ASAP7_75t_R FILLER_36_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1011 ();
 FILLER_ASAP7_75t_R FILLER_36_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1082 ();
 FILLER_ASAP7_75t_R FILLER_36_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_36_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_36_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1159 ();
 FILLER_ASAP7_75t_R FILLER_36_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_36_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1188 ();
 DECAPx4_ASAP7_75t_R FILLER_36_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1269 ();
 FILLER_ASAP7_75t_R FILLER_36_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_37_24 ();
 DECAPx2_ASAP7_75t_R FILLER_37_46 ();
 FILLER_ASAP7_75t_R FILLER_37_52 ();
 DECAPx2_ASAP7_75t_R FILLER_37_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_75 ();
 DECAPx2_ASAP7_75t_R FILLER_37_88 ();
 DECAPx6_ASAP7_75t_R FILLER_37_106 ();
 DECAPx1_ASAP7_75t_R FILLER_37_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_124 ();
 FILLER_ASAP7_75t_R FILLER_37_141 ();
 FILLER_ASAP7_75t_R FILLER_37_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_154 ();
 FILLER_ASAP7_75t_R FILLER_37_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_166 ();
 FILLER_ASAP7_75t_R FILLER_37_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_176 ();
 DECAPx4_ASAP7_75t_R FILLER_37_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_201 ();
 DECAPx4_ASAP7_75t_R FILLER_37_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_219 ();
 DECAPx10_ASAP7_75t_R FILLER_37_226 ();
 DECAPx2_ASAP7_75t_R FILLER_37_248 ();
 DECAPx4_ASAP7_75t_R FILLER_37_263 ();
 FILLER_ASAP7_75t_R FILLER_37_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_275 ();
 DECAPx2_ASAP7_75t_R FILLER_37_285 ();
 DECAPx6_ASAP7_75t_R FILLER_37_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_314 ();
 FILLER_ASAP7_75t_R FILLER_37_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_336 ();
 DECAPx1_ASAP7_75t_R FILLER_37_344 ();
 DECAPx1_ASAP7_75t_R FILLER_37_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_376 ();
 DECAPx10_ASAP7_75t_R FILLER_37_387 ();
 DECAPx1_ASAP7_75t_R FILLER_37_409 ();
 DECAPx2_ASAP7_75t_R FILLER_37_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_431 ();
 FILLER_ASAP7_75t_R FILLER_37_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_440 ();
 DECAPx2_ASAP7_75t_R FILLER_37_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_457 ();
 DECAPx10_ASAP7_75t_R FILLER_37_486 ();
 DECAPx6_ASAP7_75t_R FILLER_37_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_532 ();
 DECAPx4_ASAP7_75t_R FILLER_37_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_549 ();
 DECAPx10_ASAP7_75t_R FILLER_37_560 ();
 DECAPx6_ASAP7_75t_R FILLER_37_582 ();
 FILLER_ASAP7_75t_R FILLER_37_596 ();
 DECAPx6_ASAP7_75t_R FILLER_37_626 ();
 DECAPx2_ASAP7_75t_R FILLER_37_640 ();
 DECAPx1_ASAP7_75t_R FILLER_37_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_676 ();
 DECAPx10_ASAP7_75t_R FILLER_37_683 ();
 DECAPx2_ASAP7_75t_R FILLER_37_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_719 ();
 FILLER_ASAP7_75t_R FILLER_37_730 ();
 DECAPx4_ASAP7_75t_R FILLER_37_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_752 ();
 DECAPx4_ASAP7_75t_R FILLER_37_767 ();
 FILLER_ASAP7_75t_R FILLER_37_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_779 ();
 DECAPx10_ASAP7_75t_R FILLER_37_789 ();
 DECAPx4_ASAP7_75t_R FILLER_37_811 ();
 FILLER_ASAP7_75t_R FILLER_37_821 ();
 DECAPx6_ASAP7_75t_R FILLER_37_837 ();
 FILLER_ASAP7_75t_R FILLER_37_861 ();
 DECAPx2_ASAP7_75t_R FILLER_37_869 ();
 FILLER_ASAP7_75t_R FILLER_37_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_923 ();
 DECAPx2_ASAP7_75t_R FILLER_37_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_932 ();
 DECAPx10_ASAP7_75t_R FILLER_37_939 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1007 ();
 FILLER_ASAP7_75t_R FILLER_37_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1047 ();
 FILLER_ASAP7_75t_R FILLER_37_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1075 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_37_1111 ();
 FILLER_ASAP7_75t_R FILLER_37_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1154 ();
 FILLER_ASAP7_75t_R FILLER_37_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1205 ();
 FILLER_ASAP7_75t_R FILLER_37_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx6_ASAP7_75t_R FILLER_38_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_38 ();
 DECAPx1_ASAP7_75t_R FILLER_38_51 ();
 DECAPx4_ASAP7_75t_R FILLER_38_67 ();
 FILLER_ASAP7_75t_R FILLER_38_92 ();
 DECAPx2_ASAP7_75t_R FILLER_38_97 ();
 DECAPx10_ASAP7_75t_R FILLER_38_115 ();
 DECAPx2_ASAP7_75t_R FILLER_38_137 ();
 FILLER_ASAP7_75t_R FILLER_38_143 ();
 DECAPx2_ASAP7_75t_R FILLER_38_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_158 ();
 DECAPx1_ASAP7_75t_R FILLER_38_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_178 ();
 DECAPx2_ASAP7_75t_R FILLER_38_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_194 ();
 DECAPx2_ASAP7_75t_R FILLER_38_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_207 ();
 DECAPx10_ASAP7_75t_R FILLER_38_220 ();
 FILLER_ASAP7_75t_R FILLER_38_242 ();
 DECAPx10_ASAP7_75t_R FILLER_38_258 ();
 DECAPx6_ASAP7_75t_R FILLER_38_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_318 ();
 FILLER_ASAP7_75t_R FILLER_38_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_358 ();
 DECAPx2_ASAP7_75t_R FILLER_38_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_375 ();
 DECAPx10_ASAP7_75t_R FILLER_38_383 ();
 DECAPx4_ASAP7_75t_R FILLER_38_405 ();
 FILLER_ASAP7_75t_R FILLER_38_415 ();
 DECAPx2_ASAP7_75t_R FILLER_38_423 ();
 FILLER_ASAP7_75t_R FILLER_38_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_431 ();
 DECAPx6_ASAP7_75t_R FILLER_38_448 ();
 DECAPx4_ASAP7_75t_R FILLER_38_464 ();
 DECAPx6_ASAP7_75t_R FILLER_38_480 ();
 DECAPx1_ASAP7_75t_R FILLER_38_494 ();
 DECAPx6_ASAP7_75t_R FILLER_38_508 ();
 DECAPx2_ASAP7_75t_R FILLER_38_522 ();
 DECAPx6_ASAP7_75t_R FILLER_38_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_556 ();
 DECAPx2_ASAP7_75t_R FILLER_38_567 ();
 FILLER_ASAP7_75t_R FILLER_38_573 ();
 DECAPx4_ASAP7_75t_R FILLER_38_581 ();
 FILLER_ASAP7_75t_R FILLER_38_591 ();
 DECAPx2_ASAP7_75t_R FILLER_38_607 ();
 FILLER_ASAP7_75t_R FILLER_38_613 ();
 DECAPx10_ASAP7_75t_R FILLER_38_618 ();
 DECAPx2_ASAP7_75t_R FILLER_38_640 ();
 FILLER_ASAP7_75t_R FILLER_38_646 ();
 DECAPx4_ASAP7_75t_R FILLER_38_662 ();
 FILLER_ASAP7_75t_R FILLER_38_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_674 ();
 DECAPx2_ASAP7_75t_R FILLER_38_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_687 ();
 DECAPx10_ASAP7_75t_R FILLER_38_698 ();
 DECAPx6_ASAP7_75t_R FILLER_38_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_734 ();
 DECAPx10_ASAP7_75t_R FILLER_38_741 ();
 DECAPx4_ASAP7_75t_R FILLER_38_763 ();
 FILLER_ASAP7_75t_R FILLER_38_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_781 ();
 DECAPx6_ASAP7_75t_R FILLER_38_788 ();
 DECAPx2_ASAP7_75t_R FILLER_38_808 ();
 DECAPx4_ASAP7_75t_R FILLER_38_840 ();
 FILLER_ASAP7_75t_R FILLER_38_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_852 ();
 DECAPx10_ASAP7_75t_R FILLER_38_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_889 ();
 DECAPx4_ASAP7_75t_R FILLER_38_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_910 ();
 DECAPx1_ASAP7_75t_R FILLER_38_932 ();
 DECAPx2_ASAP7_75t_R FILLER_38_965 ();
 FILLER_ASAP7_75t_R FILLER_38_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_973 ();
 DECAPx6_ASAP7_75t_R FILLER_38_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1000 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1050 ();
 FILLER_ASAP7_75t_R FILLER_38_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1073 ();
 FILLER_ASAP7_75t_R FILLER_38_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1097 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1171 ();
 FILLER_ASAP7_75t_R FILLER_38_1185 ();
 FILLER_ASAP7_75t_R FILLER_38_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1206 ();
 FILLER_ASAP7_75t_R FILLER_38_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1248 ();
 FILLER_ASAP7_75t_R FILLER_38_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1280 ();
 FILLER_ASAP7_75t_R FILLER_38_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 DECAPx6_ASAP7_75t_R FILLER_39_24 ();
 FILLER_ASAP7_75t_R FILLER_39_38 ();
 DECAPx6_ASAP7_75t_R FILLER_39_52 ();
 FILLER_ASAP7_75t_R FILLER_39_66 ();
 FILLER_ASAP7_75t_R FILLER_39_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_97 ();
 FILLER_ASAP7_75t_R FILLER_39_107 ();
 DECAPx2_ASAP7_75t_R FILLER_39_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_127 ();
 DECAPx10_ASAP7_75t_R FILLER_39_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_162 ();
 DECAPx1_ASAP7_75t_R FILLER_39_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_174 ();
 DECAPx6_ASAP7_75t_R FILLER_39_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_192 ();
 DECAPx1_ASAP7_75t_R FILLER_39_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_221 ();
 DECAPx2_ASAP7_75t_R FILLER_39_246 ();
 FILLER_ASAP7_75t_R FILLER_39_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_279 ();
 DECAPx6_ASAP7_75t_R FILLER_39_288 ();
 DECAPx4_ASAP7_75t_R FILLER_39_309 ();
 FILLER_ASAP7_75t_R FILLER_39_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_321 ();
 DECAPx1_ASAP7_75t_R FILLER_39_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_359 ();
 DECAPx2_ASAP7_75t_R FILLER_39_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_378 ();
 DECAPx4_ASAP7_75t_R FILLER_39_396 ();
 FILLER_ASAP7_75t_R FILLER_39_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_408 ();
 DECAPx1_ASAP7_75t_R FILLER_39_415 ();
 DECAPx2_ASAP7_75t_R FILLER_39_425 ();
 FILLER_ASAP7_75t_R FILLER_39_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_455 ();
 FILLER_ASAP7_75t_R FILLER_39_476 ();
 DECAPx6_ASAP7_75t_R FILLER_39_506 ();
 FILLER_ASAP7_75t_R FILLER_39_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_522 ();
 DECAPx6_ASAP7_75t_R FILLER_39_530 ();
 FILLER_ASAP7_75t_R FILLER_39_544 ();
 FILLER_ASAP7_75t_R FILLER_39_556 ();
 DECAPx1_ASAP7_75t_R FILLER_39_568 ();
 DECAPx6_ASAP7_75t_R FILLER_39_596 ();
 DECAPx10_ASAP7_75t_R FILLER_39_626 ();
 DECAPx6_ASAP7_75t_R FILLER_39_648 ();
 FILLER_ASAP7_75t_R FILLER_39_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_664 ();
 DECAPx6_ASAP7_75t_R FILLER_39_683 ();
 DECAPx1_ASAP7_75t_R FILLER_39_697 ();
 DECAPx10_ASAP7_75t_R FILLER_39_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_733 ();
 DECAPx6_ASAP7_75t_R FILLER_39_750 ();
 FILLER_ASAP7_75t_R FILLER_39_764 ();
 DECAPx10_ASAP7_75t_R FILLER_39_772 ();
 DECAPx1_ASAP7_75t_R FILLER_39_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_798 ();
 DECAPx4_ASAP7_75t_R FILLER_39_805 ();
 DECAPx1_ASAP7_75t_R FILLER_39_832 ();
 DECAPx1_ASAP7_75t_R FILLER_39_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_870 ();
 DECAPx2_ASAP7_75t_R FILLER_39_892 ();
 FILLER_ASAP7_75t_R FILLER_39_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_900 ();
 DECAPx1_ASAP7_75t_R FILLER_39_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_923 ();
 DECAPx2_ASAP7_75t_R FILLER_39_947 ();
 FILLER_ASAP7_75t_R FILLER_39_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_955 ();
 DECAPx2_ASAP7_75t_R FILLER_39_985 ();
 FILLER_ASAP7_75t_R FILLER_39_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_993 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1079 ();
 FILLER_ASAP7_75t_R FILLER_39_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1177 ();
 FILLER_ASAP7_75t_R FILLER_39_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1208 ();
 FILLER_ASAP7_75t_R FILLER_39_1215 ();
 FILLER_ASAP7_75t_R FILLER_39_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1239 ();
 FILLER_ASAP7_75t_R FILLER_39_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_39_1276 ();
 FILLER_ASAP7_75t_R FILLER_39_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx6_ASAP7_75t_R FILLER_40_24 ();
 DECAPx1_ASAP7_75t_R FILLER_40_38 ();
 DECAPx1_ASAP7_75t_R FILLER_40_61 ();
 DECAPx1_ASAP7_75t_R FILLER_40_80 ();
 FILLER_ASAP7_75t_R FILLER_40_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_108 ();
 DECAPx2_ASAP7_75t_R FILLER_40_130 ();
 FILLER_ASAP7_75t_R FILLER_40_136 ();
 DECAPx10_ASAP7_75t_R FILLER_40_150 ();
 DECAPx4_ASAP7_75t_R FILLER_40_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_182 ();
 DECAPx2_ASAP7_75t_R FILLER_40_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_207 ();
 DECAPx2_ASAP7_75t_R FILLER_40_221 ();
 FILLER_ASAP7_75t_R FILLER_40_227 ();
 FILLER_ASAP7_75t_R FILLER_40_250 ();
 DECAPx1_ASAP7_75t_R FILLER_40_296 ();
 FILLER_ASAP7_75t_R FILLER_40_310 ();
 DECAPx10_ASAP7_75t_R FILLER_40_319 ();
 DECAPx4_ASAP7_75t_R FILLER_40_341 ();
 FILLER_ASAP7_75t_R FILLER_40_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_353 ();
 DECAPx2_ASAP7_75t_R FILLER_40_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_366 ();
 FILLER_ASAP7_75t_R FILLER_40_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_377 ();
 DECAPx2_ASAP7_75t_R FILLER_40_399 ();
 DECAPx2_ASAP7_75t_R FILLER_40_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_427 ();
 DECAPx2_ASAP7_75t_R FILLER_40_454 ();
 FILLER_ASAP7_75t_R FILLER_40_460 ();
 DECAPx2_ASAP7_75t_R FILLER_40_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_470 ();
 DECAPx2_ASAP7_75t_R FILLER_40_479 ();
 FILLER_ASAP7_75t_R FILLER_40_485 ();
 DECAPx1_ASAP7_75t_R FILLER_40_493 ();
 DECAPx1_ASAP7_75t_R FILLER_40_507 ();
 FILLER_ASAP7_75t_R FILLER_40_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_523 ();
 FILLER_ASAP7_75t_R FILLER_40_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_544 ();
 FILLER_ASAP7_75t_R FILLER_40_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_554 ();
 DECAPx2_ASAP7_75t_R FILLER_40_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_569 ();
 FILLER_ASAP7_75t_R FILLER_40_576 ();
 DECAPx1_ASAP7_75t_R FILLER_40_585 ();
 DECAPx1_ASAP7_75t_R FILLER_40_597 ();
 DECAPx1_ASAP7_75t_R FILLER_40_609 ();
 DECAPx10_ASAP7_75t_R FILLER_40_623 ();
 DECAPx10_ASAP7_75t_R FILLER_40_645 ();
 DECAPx2_ASAP7_75t_R FILLER_40_691 ();
 FILLER_ASAP7_75t_R FILLER_40_697 ();
 DECAPx4_ASAP7_75t_R FILLER_40_709 ();
 FILLER_ASAP7_75t_R FILLER_40_719 ();
 DECAPx2_ASAP7_75t_R FILLER_40_727 ();
 FILLER_ASAP7_75t_R FILLER_40_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_735 ();
 DECAPx2_ASAP7_75t_R FILLER_40_750 ();
 FILLER_ASAP7_75t_R FILLER_40_756 ();
 DECAPx2_ASAP7_75t_R FILLER_40_774 ();
 FILLER_ASAP7_75t_R FILLER_40_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_782 ();
 DECAPx10_ASAP7_75t_R FILLER_40_789 ();
 DECAPx2_ASAP7_75t_R FILLER_40_811 ();
 FILLER_ASAP7_75t_R FILLER_40_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_819 ();
 DECAPx6_ASAP7_75t_R FILLER_40_826 ();
 DECAPx1_ASAP7_75t_R FILLER_40_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_844 ();
 DECAPx1_ASAP7_75t_R FILLER_40_855 ();
 FILLER_ASAP7_75t_R FILLER_40_875 ();
 DECAPx2_ASAP7_75t_R FILLER_40_892 ();
 DECAPx2_ASAP7_75t_R FILLER_40_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_916 ();
 DECAPx1_ASAP7_75t_R FILLER_40_923 ();
 DECAPx10_ASAP7_75t_R FILLER_40_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1011 ();
 FILLER_ASAP7_75t_R FILLER_40_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1149 ();
 FILLER_ASAP7_75t_R FILLER_40_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1210 ();
 FILLER_ASAP7_75t_R FILLER_40_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1267 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_24 ();
 DECAPx1_ASAP7_75t_R FILLER_41_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_50 ();
 DECAPx4_ASAP7_75t_R FILLER_41_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_95 ();
 DECAPx4_ASAP7_75t_R FILLER_41_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_109 ();
 DECAPx1_ASAP7_75t_R FILLER_41_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_129 ();
 FILLER_ASAP7_75t_R FILLER_41_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_168 ();
 DECAPx2_ASAP7_75t_R FILLER_41_175 ();
 FILLER_ASAP7_75t_R FILLER_41_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_199 ();
 DECAPx6_ASAP7_75t_R FILLER_41_206 ();
 FILLER_ASAP7_75t_R FILLER_41_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_222 ();
 DECAPx4_ASAP7_75t_R FILLER_41_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_240 ();
 FILLER_ASAP7_75t_R FILLER_41_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_258 ();
 DECAPx2_ASAP7_75t_R FILLER_41_273 ();
 FILLER_ASAP7_75t_R FILLER_41_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_307 ();
 DECAPx10_ASAP7_75t_R FILLER_41_318 ();
 DECAPx2_ASAP7_75t_R FILLER_41_340 ();
 DECAPx4_ASAP7_75t_R FILLER_41_355 ();
 FILLER_ASAP7_75t_R FILLER_41_365 ();
 DECAPx4_ASAP7_75t_R FILLER_41_375 ();
 FILLER_ASAP7_75t_R FILLER_41_385 ();
 DECAPx2_ASAP7_75t_R FILLER_41_395 ();
 FILLER_ASAP7_75t_R FILLER_41_401 ();
 DECAPx4_ASAP7_75t_R FILLER_41_421 ();
 FILLER_ASAP7_75t_R FILLER_41_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_433 ();
 DECAPx4_ASAP7_75t_R FILLER_41_440 ();
 DECAPx4_ASAP7_75t_R FILLER_41_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_495 ();
 DECAPx4_ASAP7_75t_R FILLER_41_502 ();
 FILLER_ASAP7_75t_R FILLER_41_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_514 ();
 DECAPx6_ASAP7_75t_R FILLER_41_527 ();
 DECAPx10_ASAP7_75t_R FILLER_41_551 ();
 DECAPx10_ASAP7_75t_R FILLER_41_573 ();
 DECAPx4_ASAP7_75t_R FILLER_41_595 ();
 FILLER_ASAP7_75t_R FILLER_41_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_614 ();
 DECAPx4_ASAP7_75t_R FILLER_41_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_635 ();
 DECAPx10_ASAP7_75t_R FILLER_41_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_667 ();
 DECAPx2_ASAP7_75t_R FILLER_41_674 ();
 FILLER_ASAP7_75t_R FILLER_41_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_682 ();
 DECAPx1_ASAP7_75t_R FILLER_41_693 ();
 FILLER_ASAP7_75t_R FILLER_41_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_723 ();
 DECAPx4_ASAP7_75t_R FILLER_41_730 ();
 FILLER_ASAP7_75t_R FILLER_41_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_742 ();
 FILLER_ASAP7_75t_R FILLER_41_749 ();
 DECAPx6_ASAP7_75t_R FILLER_41_757 ();
 DECAPx1_ASAP7_75t_R FILLER_41_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_775 ();
 DECAPx1_ASAP7_75t_R FILLER_41_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_790 ();
 FILLER_ASAP7_75t_R FILLER_41_803 ();
 DECAPx4_ASAP7_75t_R FILLER_41_811 ();
 DECAPx2_ASAP7_75t_R FILLER_41_833 ();
 DECAPx4_ASAP7_75t_R FILLER_41_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_869 ();
 FILLER_ASAP7_75t_R FILLER_41_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_888 ();
 DECAPx6_ASAP7_75t_R FILLER_41_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_913 ();
 DECAPx1_ASAP7_75t_R FILLER_41_920 ();
 DECAPx1_ASAP7_75t_R FILLER_41_981 ();
 DECAPx1_ASAP7_75t_R FILLER_41_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_995 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1084 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_41_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1237 ();
 FILLER_ASAP7_75t_R FILLER_41_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1285 ();
 FILLER_ASAP7_75t_R FILLER_41_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx6_ASAP7_75t_R FILLER_42_24 ();
 DECAPx1_ASAP7_75t_R FILLER_42_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_70 ();
 FILLER_ASAP7_75t_R FILLER_42_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_98 ();
 FILLER_ASAP7_75t_R FILLER_42_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_139 ();
 FILLER_ASAP7_75t_R FILLER_42_149 ();
 FILLER_ASAP7_75t_R FILLER_42_154 ();
 DECAPx4_ASAP7_75t_R FILLER_42_165 ();
 FILLER_ASAP7_75t_R FILLER_42_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_177 ();
 DECAPx1_ASAP7_75t_R FILLER_42_184 ();
 FILLER_ASAP7_75t_R FILLER_42_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_209 ();
 FILLER_ASAP7_75t_R FILLER_42_213 ();
 FILLER_ASAP7_75t_R FILLER_42_222 ();
 DECAPx1_ASAP7_75t_R FILLER_42_232 ();
 DECAPx1_ASAP7_75t_R FILLER_42_244 ();
 FILLER_ASAP7_75t_R FILLER_42_271 ();
 DECAPx4_ASAP7_75t_R FILLER_42_302 ();
 FILLER_ASAP7_75t_R FILLER_42_312 ();
 FILLER_ASAP7_75t_R FILLER_42_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_330 ();
 DECAPx4_ASAP7_75t_R FILLER_42_337 ();
 DECAPx2_ASAP7_75t_R FILLER_42_382 ();
 FILLER_ASAP7_75t_R FILLER_42_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_390 ();
 DECAPx2_ASAP7_75t_R FILLER_42_399 ();
 FILLER_ASAP7_75t_R FILLER_42_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_407 ();
 DECAPx1_ASAP7_75t_R FILLER_42_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_440 ();
 DECAPx1_ASAP7_75t_R FILLER_42_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_461 ();
 DECAPx2_ASAP7_75t_R FILLER_42_464 ();
 FILLER_ASAP7_75t_R FILLER_42_470 ();
 DECAPx6_ASAP7_75t_R FILLER_42_504 ();
 FILLER_ASAP7_75t_R FILLER_42_518 ();
 DECAPx1_ASAP7_75t_R FILLER_42_530 ();
 DECAPx6_ASAP7_75t_R FILLER_42_548 ();
 DECAPx2_ASAP7_75t_R FILLER_42_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_568 ();
 DECAPx10_ASAP7_75t_R FILLER_42_575 ();
 DECAPx4_ASAP7_75t_R FILLER_42_597 ();
 FILLER_ASAP7_75t_R FILLER_42_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_609 ();
 DECAPx10_ASAP7_75t_R FILLER_42_618 ();
 DECAPx10_ASAP7_75t_R FILLER_42_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_662 ();
 DECAPx2_ASAP7_75t_R FILLER_42_675 ();
 FILLER_ASAP7_75t_R FILLER_42_681 ();
 FILLER_ASAP7_75t_R FILLER_42_695 ();
 DECAPx2_ASAP7_75t_R FILLER_42_705 ();
 DECAPx4_ASAP7_75t_R FILLER_42_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_724 ();
 DECAPx4_ASAP7_75t_R FILLER_42_741 ();
 DECAPx2_ASAP7_75t_R FILLER_42_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_773 ();
 DECAPx2_ASAP7_75t_R FILLER_42_784 ();
 FILLER_ASAP7_75t_R FILLER_42_800 ();
 DECAPx2_ASAP7_75t_R FILLER_42_818 ();
 FILLER_ASAP7_75t_R FILLER_42_824 ();
 DECAPx4_ASAP7_75t_R FILLER_42_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_846 ();
 DECAPx6_ASAP7_75t_R FILLER_42_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_877 ();
 FILLER_ASAP7_75t_R FILLER_42_890 ();
 DECAPx1_ASAP7_75t_R FILLER_42_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_912 ();
 DECAPx6_ASAP7_75t_R FILLER_42_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_975 ();
 DECAPx6_ASAP7_75t_R FILLER_42_992 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1006 ();
 FILLER_ASAP7_75t_R FILLER_42_1016 ();
 FILLER_ASAP7_75t_R FILLER_42_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1038 ();
 FILLER_ASAP7_75t_R FILLER_42_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1161 ();
 FILLER_ASAP7_75t_R FILLER_42_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1200 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1263 ();
 FILLER_ASAP7_75t_R FILLER_42_1269 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1281 ();
 FILLER_ASAP7_75t_R FILLER_42_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx1_ASAP7_75t_R FILLER_43_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_59 ();
 FILLER_ASAP7_75t_R FILLER_43_70 ();
 FILLER_ASAP7_75t_R FILLER_43_78 ();
 FILLER_ASAP7_75t_R FILLER_43_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_90 ();
 DECAPx2_ASAP7_75t_R FILLER_43_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_139 ();
 DECAPx2_ASAP7_75t_R FILLER_43_164 ();
 FILLER_ASAP7_75t_R FILLER_43_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_185 ();
 FILLER_ASAP7_75t_R FILLER_43_217 ();
 DECAPx1_ASAP7_75t_R FILLER_43_227 ();
 FILLER_ASAP7_75t_R FILLER_43_243 ();
 FILLER_ASAP7_75t_R FILLER_43_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_253 ();
 FILLER_ASAP7_75t_R FILLER_43_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_263 ();
 FILLER_ASAP7_75t_R FILLER_43_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_272 ();
 DECAPx2_ASAP7_75t_R FILLER_43_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_316 ();
 FILLER_ASAP7_75t_R FILLER_43_337 ();
 DECAPx2_ASAP7_75t_R FILLER_43_360 ();
 FILLER_ASAP7_75t_R FILLER_43_366 ();
 DECAPx6_ASAP7_75t_R FILLER_43_375 ();
 DECAPx10_ASAP7_75t_R FILLER_43_399 ();
 DECAPx4_ASAP7_75t_R FILLER_43_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_431 ();
 FILLER_ASAP7_75t_R FILLER_43_438 ();
 DECAPx4_ASAP7_75t_R FILLER_43_466 ();
 FILLER_ASAP7_75t_R FILLER_43_476 ();
 DECAPx10_ASAP7_75t_R FILLER_43_498 ();
 DECAPx10_ASAP7_75t_R FILLER_43_520 ();
 DECAPx10_ASAP7_75t_R FILLER_43_542 ();
 DECAPx2_ASAP7_75t_R FILLER_43_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_570 ();
 DECAPx4_ASAP7_75t_R FILLER_43_577 ();
 FILLER_ASAP7_75t_R FILLER_43_587 ();
 DECAPx6_ASAP7_75t_R FILLER_43_595 ();
 FILLER_ASAP7_75t_R FILLER_43_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_611 ();
 DECAPx6_ASAP7_75t_R FILLER_43_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_634 ();
 DECAPx10_ASAP7_75t_R FILLER_43_641 ();
 DECAPx10_ASAP7_75t_R FILLER_43_663 ();
 DECAPx6_ASAP7_75t_R FILLER_43_685 ();
 DECAPx1_ASAP7_75t_R FILLER_43_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_703 ();
 FILLER_ASAP7_75t_R FILLER_43_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_716 ();
 DECAPx10_ASAP7_75t_R FILLER_43_723 ();
 DECAPx4_ASAP7_75t_R FILLER_43_745 ();
 DECAPx6_ASAP7_75t_R FILLER_43_773 ();
 DECAPx2_ASAP7_75t_R FILLER_43_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_793 ();
 DECAPx10_ASAP7_75t_R FILLER_43_804 ();
 DECAPx10_ASAP7_75t_R FILLER_43_826 ();
 DECAPx2_ASAP7_75t_R FILLER_43_848 ();
 DECAPx1_ASAP7_75t_R FILLER_43_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_870 ();
 FILLER_ASAP7_75t_R FILLER_43_900 ();
 DECAPx6_ASAP7_75t_R FILLER_43_908 ();
 FILLER_ASAP7_75t_R FILLER_43_922 ();
 DECAPx2_ASAP7_75t_R FILLER_43_947 ();
 FILLER_ASAP7_75t_R FILLER_43_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_955 ();
 DECAPx1_ASAP7_75t_R FILLER_43_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_985 ();
 DECAPx1_ASAP7_75t_R FILLER_43_992 ();
 DECAPx6_ASAP7_75t_R FILLER_43_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1034 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1046 ();
 FILLER_ASAP7_75t_R FILLER_43_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_43_1087 ();
 FILLER_ASAP7_75t_R FILLER_43_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1162 ();
 FILLER_ASAP7_75t_R FILLER_43_1184 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1200 ();
 FILLER_ASAP7_75t_R FILLER_43_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1239 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx2_ASAP7_75t_R FILLER_44_24 ();
 FILLER_ASAP7_75t_R FILLER_44_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_51 ();
 FILLER_ASAP7_75t_R FILLER_44_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_60 ();
 DECAPx1_ASAP7_75t_R FILLER_44_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_86 ();
 DECAPx6_ASAP7_75t_R FILLER_44_94 ();
 DECAPx10_ASAP7_75t_R FILLER_44_114 ();
 DECAPx10_ASAP7_75t_R FILLER_44_136 ();
 DECAPx6_ASAP7_75t_R FILLER_44_158 ();
 FILLER_ASAP7_75t_R FILLER_44_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_174 ();
 FILLER_ASAP7_75t_R FILLER_44_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_199 ();
 FILLER_ASAP7_75t_R FILLER_44_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_208 ();
 FILLER_ASAP7_75t_R FILLER_44_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_218 ();
 DECAPx1_ASAP7_75t_R FILLER_44_229 ();
 DECAPx4_ASAP7_75t_R FILLER_44_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_258 ();
 DECAPx4_ASAP7_75t_R FILLER_44_266 ();
 DECAPx1_ASAP7_75t_R FILLER_44_282 ();
 DECAPx1_ASAP7_75t_R FILLER_44_292 ();
 DECAPx10_ASAP7_75t_R FILLER_44_302 ();
 DECAPx2_ASAP7_75t_R FILLER_44_324 ();
 FILLER_ASAP7_75t_R FILLER_44_330 ();
 FILLER_ASAP7_75t_R FILLER_44_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_344 ();
 DECAPx10_ASAP7_75t_R FILLER_44_383 ();
 DECAPx4_ASAP7_75t_R FILLER_44_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_415 ();
 DECAPx6_ASAP7_75t_R FILLER_44_422 ();
 DECAPx2_ASAP7_75t_R FILLER_44_456 ();
 DECAPx4_ASAP7_75t_R FILLER_44_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_474 ();
 FILLER_ASAP7_75t_R FILLER_44_489 ();
 DECAPx10_ASAP7_75t_R FILLER_44_501 ();
 DECAPx10_ASAP7_75t_R FILLER_44_523 ();
 DECAPx10_ASAP7_75t_R FILLER_44_545 ();
 DECAPx10_ASAP7_75t_R FILLER_44_567 ();
 FILLER_ASAP7_75t_R FILLER_44_589 ();
 DECAPx10_ASAP7_75t_R FILLER_44_599 ();
 DECAPx6_ASAP7_75t_R FILLER_44_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_635 ();
 DECAPx1_ASAP7_75t_R FILLER_44_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_648 ();
 DECAPx10_ASAP7_75t_R FILLER_44_655 ();
 DECAPx10_ASAP7_75t_R FILLER_44_677 ();
 DECAPx4_ASAP7_75t_R FILLER_44_699 ();
 FILLER_ASAP7_75t_R FILLER_44_709 ();
 DECAPx6_ASAP7_75t_R FILLER_44_723 ();
 FILLER_ASAP7_75t_R FILLER_44_747 ();
 DECAPx10_ASAP7_75t_R FILLER_44_785 ();
 DECAPx2_ASAP7_75t_R FILLER_44_807 ();
 DECAPx10_ASAP7_75t_R FILLER_44_819 ();
 DECAPx4_ASAP7_75t_R FILLER_44_841 ();
 FILLER_ASAP7_75t_R FILLER_44_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_861 ();
 DECAPx4_ASAP7_75t_R FILLER_44_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_882 ();
 FILLER_ASAP7_75t_R FILLER_44_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_888 ();
 DECAPx6_ASAP7_75t_R FILLER_44_911 ();
 FILLER_ASAP7_75t_R FILLER_44_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_935 ();
 DECAPx10_ASAP7_75t_R FILLER_44_939 ();
 DECAPx10_ASAP7_75t_R FILLER_44_961 ();
 DECAPx4_ASAP7_75t_R FILLER_44_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_993 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1064 ();
 FILLER_ASAP7_75t_R FILLER_44_1086 ();
 FILLER_ASAP7_75t_R FILLER_44_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1149 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1166 ();
 FILLER_ASAP7_75t_R FILLER_44_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1199 ();
 FILLER_ASAP7_75t_R FILLER_44_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_45_2 ();
 FILLER_ASAP7_75t_R FILLER_45_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_18 ();
 FILLER_ASAP7_75t_R FILLER_45_31 ();
 DECAPx10_ASAP7_75t_R FILLER_45_51 ();
 DECAPx4_ASAP7_75t_R FILLER_45_73 ();
 FILLER_ASAP7_75t_R FILLER_45_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_85 ();
 DECAPx1_ASAP7_75t_R FILLER_45_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_97 ();
 DECAPx2_ASAP7_75t_R FILLER_45_122 ();
 DECAPx2_ASAP7_75t_R FILLER_45_150 ();
 DECAPx6_ASAP7_75t_R FILLER_45_167 ();
 DECAPx4_ASAP7_75t_R FILLER_45_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_220 ();
 FILLER_ASAP7_75t_R FILLER_45_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_230 ();
 DECAPx6_ASAP7_75t_R FILLER_45_238 ();
 DECAPx2_ASAP7_75t_R FILLER_45_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_258 ();
 DECAPx10_ASAP7_75t_R FILLER_45_266 ();
 DECAPx4_ASAP7_75t_R FILLER_45_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_314 ();
 DECAPx1_ASAP7_75t_R FILLER_45_353 ();
 DECAPx4_ASAP7_75t_R FILLER_45_367 ();
 FILLER_ASAP7_75t_R FILLER_45_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_379 ();
 DECAPx4_ASAP7_75t_R FILLER_45_401 ();
 FILLER_ASAP7_75t_R FILLER_45_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_423 ();
 DECAPx2_ASAP7_75t_R FILLER_45_442 ();
 FILLER_ASAP7_75t_R FILLER_45_448 ();
 DECAPx4_ASAP7_75t_R FILLER_45_462 ();
 FILLER_ASAP7_75t_R FILLER_45_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_474 ();
 FILLER_ASAP7_75t_R FILLER_45_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_483 ();
 FILLER_ASAP7_75t_R FILLER_45_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_492 ();
 DECAPx6_ASAP7_75t_R FILLER_45_499 ();
 FILLER_ASAP7_75t_R FILLER_45_513 ();
 DECAPx4_ASAP7_75t_R FILLER_45_529 ();
 FILLER_ASAP7_75t_R FILLER_45_539 ();
 FILLER_ASAP7_75t_R FILLER_45_548 ();
 DECAPx1_ASAP7_75t_R FILLER_45_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_560 ();
 DECAPx2_ASAP7_75t_R FILLER_45_567 ();
 FILLER_ASAP7_75t_R FILLER_45_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_575 ();
 DECAPx1_ASAP7_75t_R FILLER_45_588 ();
 DECAPx6_ASAP7_75t_R FILLER_45_602 ();
 FILLER_ASAP7_75t_R FILLER_45_616 ();
 DECAPx2_ASAP7_75t_R FILLER_45_630 ();
 FILLER_ASAP7_75t_R FILLER_45_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_644 ();
 DECAPx10_ASAP7_75t_R FILLER_45_657 ();
 DECAPx6_ASAP7_75t_R FILLER_45_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_743 ();
 FILLER_ASAP7_75t_R FILLER_45_750 ();
 FILLER_ASAP7_75t_R FILLER_45_760 ();
 FILLER_ASAP7_75t_R FILLER_45_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_778 ();
 DECAPx10_ASAP7_75t_R FILLER_45_785 ();
 DECAPx6_ASAP7_75t_R FILLER_45_807 ();
 DECAPx1_ASAP7_75t_R FILLER_45_821 ();
 FILLER_ASAP7_75t_R FILLER_45_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_840 ();
 DECAPx1_ASAP7_75t_R FILLER_45_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_859 ();
 DECAPx4_ASAP7_75t_R FILLER_45_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_882 ();
 DECAPx10_ASAP7_75t_R FILLER_45_895 ();
 DECAPx2_ASAP7_75t_R FILLER_45_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_923 ();
 DECAPx6_ASAP7_75t_R FILLER_45_926 ();
 FILLER_ASAP7_75t_R FILLER_45_940 ();
 DECAPx2_ASAP7_75t_R FILLER_45_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_964 ();
 DECAPx6_ASAP7_75t_R FILLER_45_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_988 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1016 ();
 FILLER_ASAP7_75t_R FILLER_45_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1025 ();
 FILLER_ASAP7_75t_R FILLER_45_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1044 ();
 FILLER_ASAP7_75t_R FILLER_45_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1052 ();
 DECAPx4_ASAP7_75t_R FILLER_45_1069 ();
 FILLER_ASAP7_75t_R FILLER_45_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1190 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1225 ();
 FILLER_ASAP7_75t_R FILLER_45_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1249 ();
 FILLER_ASAP7_75t_R FILLER_45_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_45_1280 ();
 FILLER_ASAP7_75t_R FILLER_45_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_46_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_16 ();
 DECAPx4_ASAP7_75t_R FILLER_46_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_55 ();
 DECAPx1_ASAP7_75t_R FILLER_46_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_66 ();
 DECAPx2_ASAP7_75t_R FILLER_46_73 ();
 FILLER_ASAP7_75t_R FILLER_46_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_145 ();
 DECAPx10_ASAP7_75t_R FILLER_46_153 ();
 DECAPx2_ASAP7_75t_R FILLER_46_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_181 ();
 DECAPx1_ASAP7_75t_R FILLER_46_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_209 ();
 DECAPx1_ASAP7_75t_R FILLER_46_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_242 ();
 DECAPx6_ASAP7_75t_R FILLER_46_249 ();
 DECAPx2_ASAP7_75t_R FILLER_46_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_269 ();
 FILLER_ASAP7_75t_R FILLER_46_289 ();
 DECAPx4_ASAP7_75t_R FILLER_46_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_311 ();
 DECAPx1_ASAP7_75t_R FILLER_46_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_326 ();
 DECAPx2_ASAP7_75t_R FILLER_46_334 ();
 DECAPx10_ASAP7_75t_R FILLER_46_347 ();
 DECAPx4_ASAP7_75t_R FILLER_46_369 ();
 DECAPx2_ASAP7_75t_R FILLER_46_396 ();
 FILLER_ASAP7_75t_R FILLER_46_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_404 ();
 DECAPx6_ASAP7_75t_R FILLER_46_411 ();
 FILLER_ASAP7_75t_R FILLER_46_425 ();
 DECAPx2_ASAP7_75t_R FILLER_46_440 ();
 DECAPx2_ASAP7_75t_R FILLER_46_464 ();
 FILLER_ASAP7_75t_R FILLER_46_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_472 ();
 DECAPx10_ASAP7_75t_R FILLER_46_482 ();
 FILLER_ASAP7_75t_R FILLER_46_520 ();
 DECAPx10_ASAP7_75t_R FILLER_46_538 ();
 DECAPx10_ASAP7_75t_R FILLER_46_560 ();
 DECAPx10_ASAP7_75t_R FILLER_46_582 ();
 DECAPx10_ASAP7_75t_R FILLER_46_604 ();
 DECAPx4_ASAP7_75t_R FILLER_46_626 ();
 FILLER_ASAP7_75t_R FILLER_46_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_638 ();
 DECAPx2_ASAP7_75t_R FILLER_46_660 ();
 FILLER_ASAP7_75t_R FILLER_46_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_668 ();
 DECAPx2_ASAP7_75t_R FILLER_46_679 ();
 FILLER_ASAP7_75t_R FILLER_46_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_687 ();
 DECAPx1_ASAP7_75t_R FILLER_46_694 ();
 DECAPx10_ASAP7_75t_R FILLER_46_711 ();
 DECAPx6_ASAP7_75t_R FILLER_46_733 ();
 DECAPx2_ASAP7_75t_R FILLER_46_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_753 ();
 DECAPx10_ASAP7_75t_R FILLER_46_764 ();
 DECAPx6_ASAP7_75t_R FILLER_46_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_800 ();
 DECAPx10_ASAP7_75t_R FILLER_46_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_847 ();
 DECAPx6_ASAP7_75t_R FILLER_46_858 ();
 DECAPx6_ASAP7_75t_R FILLER_46_875 ();
 DECAPx1_ASAP7_75t_R FILLER_46_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_917 ();
 DECAPx6_ASAP7_75t_R FILLER_46_930 ();
 DECAPx1_ASAP7_75t_R FILLER_46_953 ();
 DECAPx6_ASAP7_75t_R FILLER_46_963 ();
 DECAPx2_ASAP7_75t_R FILLER_46_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_983 ();
 DECAPx6_ASAP7_75t_R FILLER_46_992 ();
 FILLER_ASAP7_75t_R FILLER_46_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1039 ();
 FILLER_ASAP7_75t_R FILLER_46_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1070 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1092 ();
 FILLER_ASAP7_75t_R FILLER_46_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1160 ();
 FILLER_ASAP7_75t_R FILLER_46_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1168 ();
 FILLER_ASAP7_75t_R FILLER_46_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1177 ();
 FILLER_ASAP7_75t_R FILLER_46_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1203 ();
 FILLER_ASAP7_75t_R FILLER_46_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx6_ASAP7_75t_R FILLER_47_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_38 ();
 DECAPx1_ASAP7_75t_R FILLER_47_45 ();
 DECAPx2_ASAP7_75t_R FILLER_47_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_81 ();
 DECAPx1_ASAP7_75t_R FILLER_47_85 ();
 FILLER_ASAP7_75t_R FILLER_47_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_98 ();
 DECAPx1_ASAP7_75t_R FILLER_47_111 ();
 DECAPx1_ASAP7_75t_R FILLER_47_122 ();
 FILLER_ASAP7_75t_R FILLER_47_141 ();
 DECAPx4_ASAP7_75t_R FILLER_47_167 ();
 DECAPx2_ASAP7_75t_R FILLER_47_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_194 ();
 DECAPx4_ASAP7_75t_R FILLER_47_201 ();
 FILLER_ASAP7_75t_R FILLER_47_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_213 ();
 DECAPx4_ASAP7_75t_R FILLER_47_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_244 ();
 DECAPx6_ASAP7_75t_R FILLER_47_254 ();
 DECAPx1_ASAP7_75t_R FILLER_47_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_272 ();
 FILLER_ASAP7_75t_R FILLER_47_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_290 ();
 DECAPx6_ASAP7_75t_R FILLER_47_301 ();
 DECAPx1_ASAP7_75t_R FILLER_47_315 ();
 DECAPx1_ASAP7_75t_R FILLER_47_334 ();
 DECAPx10_ASAP7_75t_R FILLER_47_348 ();
 FILLER_ASAP7_75t_R FILLER_47_370 ();
 FILLER_ASAP7_75t_R FILLER_47_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_381 ();
 DECAPx6_ASAP7_75t_R FILLER_47_392 ();
 FILLER_ASAP7_75t_R FILLER_47_406 ();
 DECAPx1_ASAP7_75t_R FILLER_47_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_418 ();
 FILLER_ASAP7_75t_R FILLER_47_429 ();
 DECAPx10_ASAP7_75t_R FILLER_47_439 ();
 FILLER_ASAP7_75t_R FILLER_47_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_463 ();
 DECAPx10_ASAP7_75t_R FILLER_47_486 ();
 DECAPx10_ASAP7_75t_R FILLER_47_508 ();
 DECAPx10_ASAP7_75t_R FILLER_47_530 ();
 DECAPx10_ASAP7_75t_R FILLER_47_552 ();
 DECAPx10_ASAP7_75t_R FILLER_47_574 ();
 DECAPx10_ASAP7_75t_R FILLER_47_596 ();
 DECAPx10_ASAP7_75t_R FILLER_47_618 ();
 DECAPx10_ASAP7_75t_R FILLER_47_640 ();
 DECAPx10_ASAP7_75t_R FILLER_47_662 ();
 DECAPx10_ASAP7_75t_R FILLER_47_684 ();
 DECAPx10_ASAP7_75t_R FILLER_47_706 ();
 DECAPx6_ASAP7_75t_R FILLER_47_728 ();
 DECAPx2_ASAP7_75t_R FILLER_47_742 ();
 DECAPx6_ASAP7_75t_R FILLER_47_758 ();
 FILLER_ASAP7_75t_R FILLER_47_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_774 ();
 DECAPx10_ASAP7_75t_R FILLER_47_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_807 ();
 FILLER_ASAP7_75t_R FILLER_47_814 ();
 DECAPx4_ASAP7_75t_R FILLER_47_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_852 ();
 DECAPx10_ASAP7_75t_R FILLER_47_886 ();
 DECAPx2_ASAP7_75t_R FILLER_47_908 ();
 FILLER_ASAP7_75t_R FILLER_47_914 ();
 FILLER_ASAP7_75t_R FILLER_47_922 ();
 DECAPx2_ASAP7_75t_R FILLER_47_970 ();
 FILLER_ASAP7_75t_R FILLER_47_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_978 ();
 DECAPx4_ASAP7_75t_R FILLER_47_994 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_47_1038 ();
 FILLER_ASAP7_75t_R FILLER_47_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1060 ();
 FILLER_ASAP7_75t_R FILLER_47_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1074 ();
 FILLER_ASAP7_75t_R FILLER_47_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1121 ();
 FILLER_ASAP7_75t_R FILLER_47_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1136 ();
 FILLER_ASAP7_75t_R FILLER_47_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_47_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_48_2 ();
 DECAPx1_ASAP7_75t_R FILLER_48_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_28 ();
 DECAPx2_ASAP7_75t_R FILLER_48_35 ();
 FILLER_ASAP7_75t_R FILLER_48_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_50 ();
 FILLER_ASAP7_75t_R FILLER_48_57 ();
 DECAPx2_ASAP7_75t_R FILLER_48_71 ();
 DECAPx1_ASAP7_75t_R FILLER_48_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_124 ();
 DECAPx1_ASAP7_75t_R FILLER_48_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_150 ();
 DECAPx6_ASAP7_75t_R FILLER_48_163 ();
 DECAPx1_ASAP7_75t_R FILLER_48_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_181 ();
 DECAPx2_ASAP7_75t_R FILLER_48_188 ();
 FILLER_ASAP7_75t_R FILLER_48_194 ();
 DECAPx1_ASAP7_75t_R FILLER_48_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_215 ();
 FILLER_ASAP7_75t_R FILLER_48_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_230 ();
 FILLER_ASAP7_75t_R FILLER_48_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_243 ();
 DECAPx6_ASAP7_75t_R FILLER_48_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_273 ();
 DECAPx2_ASAP7_75t_R FILLER_48_280 ();
 FILLER_ASAP7_75t_R FILLER_48_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_296 ();
 DECAPx6_ASAP7_75t_R FILLER_48_319 ();
 DECAPx1_ASAP7_75t_R FILLER_48_333 ();
 DECAPx4_ASAP7_75t_R FILLER_48_344 ();
 DECAPx2_ASAP7_75t_R FILLER_48_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_377 ();
 DECAPx2_ASAP7_75t_R FILLER_48_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_405 ();
 DECAPx2_ASAP7_75t_R FILLER_48_428 ();
 DECAPx1_ASAP7_75t_R FILLER_48_440 ();
 DECAPx10_ASAP7_75t_R FILLER_48_464 ();
 DECAPx2_ASAP7_75t_R FILLER_48_486 ();
 FILLER_ASAP7_75t_R FILLER_48_492 ();
 DECAPx2_ASAP7_75t_R FILLER_48_506 ();
 FILLER_ASAP7_75t_R FILLER_48_512 ();
 FILLER_ASAP7_75t_R FILLER_48_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_526 ();
 DECAPx10_ASAP7_75t_R FILLER_48_535 ();
 DECAPx6_ASAP7_75t_R FILLER_48_557 ();
 DECAPx2_ASAP7_75t_R FILLER_48_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_577 ();
 DECAPx4_ASAP7_75t_R FILLER_48_594 ();
 DECAPx10_ASAP7_75t_R FILLER_48_621 ();
 DECAPx10_ASAP7_75t_R FILLER_48_643 ();
 DECAPx10_ASAP7_75t_R FILLER_48_665 ();
 DECAPx10_ASAP7_75t_R FILLER_48_687 ();
 DECAPx10_ASAP7_75t_R FILLER_48_709 ();
 DECAPx2_ASAP7_75t_R FILLER_48_731 ();
 FILLER_ASAP7_75t_R FILLER_48_737 ();
 DECAPx2_ASAP7_75t_R FILLER_48_745 ();
 DECAPx10_ASAP7_75t_R FILLER_48_765 ();
 DECAPx6_ASAP7_75t_R FILLER_48_787 ();
 DECAPx1_ASAP7_75t_R FILLER_48_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_805 ();
 DECAPx2_ASAP7_75t_R FILLER_48_824 ();
 FILLER_ASAP7_75t_R FILLER_48_830 ();
 DECAPx6_ASAP7_75t_R FILLER_48_842 ();
 FILLER_ASAP7_75t_R FILLER_48_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_858 ();
 DECAPx10_ASAP7_75t_R FILLER_48_871 ();
 DECAPx2_ASAP7_75t_R FILLER_48_893 ();
 DECAPx4_ASAP7_75t_R FILLER_48_905 ();
 DECAPx2_ASAP7_75t_R FILLER_48_925 ();
 FILLER_ASAP7_75t_R FILLER_48_961 ();
 FILLER_ASAP7_75t_R FILLER_48_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_971 ();
 DECAPx10_ASAP7_75t_R FILLER_48_982 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1026 ();
 FILLER_ASAP7_75t_R FILLER_48_1036 ();
 FILLER_ASAP7_75t_R FILLER_48_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1046 ();
 FILLER_ASAP7_75t_R FILLER_48_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1097 ();
 FILLER_ASAP7_75t_R FILLER_48_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1243 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_49_2 ();
 DECAPx2_ASAP7_75t_R FILLER_49_16 ();
 FILLER_ASAP7_75t_R FILLER_49_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_41 ();
 DECAPx4_ASAP7_75t_R FILLER_49_68 ();
 FILLER_ASAP7_75t_R FILLER_49_78 ();
 DECAPx2_ASAP7_75t_R FILLER_49_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_101 ();
 DECAPx1_ASAP7_75t_R FILLER_49_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_113 ();
 DECAPx6_ASAP7_75t_R FILLER_49_121 ();
 DECAPx2_ASAP7_75t_R FILLER_49_135 ();
 DECAPx1_ASAP7_75t_R FILLER_49_153 ();
 FILLER_ASAP7_75t_R FILLER_49_166 ();
 FILLER_ASAP7_75t_R FILLER_49_172 ();
 DECAPx2_ASAP7_75t_R FILLER_49_186 ();
 DECAPx2_ASAP7_75t_R FILLER_49_202 ();
 FILLER_ASAP7_75t_R FILLER_49_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_210 ();
 DECAPx4_ASAP7_75t_R FILLER_49_217 ();
 FILLER_ASAP7_75t_R FILLER_49_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_229 ();
 DECAPx2_ASAP7_75t_R FILLER_49_237 ();
 DECAPx2_ASAP7_75t_R FILLER_49_262 ();
 DECAPx10_ASAP7_75t_R FILLER_49_278 ();
 DECAPx4_ASAP7_75t_R FILLER_49_300 ();
 FILLER_ASAP7_75t_R FILLER_49_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_312 ();
 DECAPx4_ASAP7_75t_R FILLER_49_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_385 ();
 FILLER_ASAP7_75t_R FILLER_49_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_415 ();
 FILLER_ASAP7_75t_R FILLER_49_426 ();
 DECAPx1_ASAP7_75t_R FILLER_49_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_448 ();
 DECAPx4_ASAP7_75t_R FILLER_49_461 ();
 FILLER_ASAP7_75t_R FILLER_49_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_473 ();
 DECAPx6_ASAP7_75t_R FILLER_49_505 ();
 DECAPx1_ASAP7_75t_R FILLER_49_519 ();
 DECAPx4_ASAP7_75t_R FILLER_49_537 ();
 FILLER_ASAP7_75t_R FILLER_49_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_549 ();
 DECAPx1_ASAP7_75t_R FILLER_49_557 ();
 DECAPx6_ASAP7_75t_R FILLER_49_587 ();
 DECAPx1_ASAP7_75t_R FILLER_49_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_605 ();
 DECAPx4_ASAP7_75t_R FILLER_49_616 ();
 FILLER_ASAP7_75t_R FILLER_49_626 ();
 DECAPx4_ASAP7_75t_R FILLER_49_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_654 ();
 DECAPx2_ASAP7_75t_R FILLER_49_667 ();
 FILLER_ASAP7_75t_R FILLER_49_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_675 ();
 DECAPx2_ASAP7_75t_R FILLER_49_686 ();
 DECAPx10_ASAP7_75t_R FILLER_49_716 ();
 FILLER_ASAP7_75t_R FILLER_49_738 ();
 DECAPx2_ASAP7_75t_R FILLER_49_750 ();
 FILLER_ASAP7_75t_R FILLER_49_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_758 ();
 DECAPx10_ASAP7_75t_R FILLER_49_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_793 ();
 DECAPx10_ASAP7_75t_R FILLER_49_805 ();
 DECAPx4_ASAP7_75t_R FILLER_49_827 ();
 FILLER_ASAP7_75t_R FILLER_49_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_839 ();
 DECAPx10_ASAP7_75t_R FILLER_49_846 ();
 DECAPx6_ASAP7_75t_R FILLER_49_868 ();
 DECAPx1_ASAP7_75t_R FILLER_49_882 ();
 DECAPx1_ASAP7_75t_R FILLER_49_898 ();
 DECAPx6_ASAP7_75t_R FILLER_49_908 ();
 FILLER_ASAP7_75t_R FILLER_49_922 ();
 DECAPx1_ASAP7_75t_R FILLER_49_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_930 ();
 FILLER_ASAP7_75t_R FILLER_49_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_977 ();
 DECAPx4_ASAP7_75t_R FILLER_49_985 ();
 FILLER_ASAP7_75t_R FILLER_49_995 ();
 FILLER_ASAP7_75t_R FILLER_49_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_49_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1056 ();
 FILLER_ASAP7_75t_R FILLER_49_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_49_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_49_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1143 ();
 FILLER_ASAP7_75t_R FILLER_49_1153 ();
 FILLER_ASAP7_75t_R FILLER_49_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_50_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_40 ();
 FILLER_ASAP7_75t_R FILLER_50_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_49 ();
 FILLER_ASAP7_75t_R FILLER_50_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_58 ();
 DECAPx4_ASAP7_75t_R FILLER_50_66 ();
 FILLER_ASAP7_75t_R FILLER_50_76 ();
 DECAPx2_ASAP7_75t_R FILLER_50_93 ();
 DECAPx1_ASAP7_75t_R FILLER_50_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_109 ();
 DECAPx4_ASAP7_75t_R FILLER_50_122 ();
 FILLER_ASAP7_75t_R FILLER_50_132 ();
 DECAPx4_ASAP7_75t_R FILLER_50_155 ();
 FILLER_ASAP7_75t_R FILLER_50_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_192 ();
 FILLER_ASAP7_75t_R FILLER_50_199 ();
 DECAPx2_ASAP7_75t_R FILLER_50_207 ();
 FILLER_ASAP7_75t_R FILLER_50_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_222 ();
 FILLER_ASAP7_75t_R FILLER_50_229 ();
 FILLER_ASAP7_75t_R FILLER_50_237 ();
 FILLER_ASAP7_75t_R FILLER_50_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_250 ();
 DECAPx6_ASAP7_75t_R FILLER_50_260 ();
 DECAPx2_ASAP7_75t_R FILLER_50_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_294 ();
 DECAPx4_ASAP7_75t_R FILLER_50_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_313 ();
 DECAPx6_ASAP7_75t_R FILLER_50_329 ();
 FILLER_ASAP7_75t_R FILLER_50_343 ();
 FILLER_ASAP7_75t_R FILLER_50_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_355 ();
 DECAPx1_ASAP7_75t_R FILLER_50_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_375 ();
 DECAPx6_ASAP7_75t_R FILLER_50_416 ();
 DECAPx2_ASAP7_75t_R FILLER_50_430 ();
 FILLER_ASAP7_75t_R FILLER_50_442 ();
 DECAPx1_ASAP7_75t_R FILLER_50_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_461 ();
 DECAPx2_ASAP7_75t_R FILLER_50_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_470 ();
 DECAPx10_ASAP7_75t_R FILLER_50_488 ();
 DECAPx10_ASAP7_75t_R FILLER_50_510 ();
 DECAPx2_ASAP7_75t_R FILLER_50_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_538 ();
 DECAPx2_ASAP7_75t_R FILLER_50_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_576 ();
 DECAPx10_ASAP7_75t_R FILLER_50_591 ();
 DECAPx1_ASAP7_75t_R FILLER_50_613 ();
 DECAPx2_ASAP7_75t_R FILLER_50_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_630 ();
 DECAPx2_ASAP7_75t_R FILLER_50_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_643 ();
 DECAPx10_ASAP7_75t_R FILLER_50_654 ();
 DECAPx2_ASAP7_75t_R FILLER_50_676 ();
 FILLER_ASAP7_75t_R FILLER_50_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_684 ();
 DECAPx6_ASAP7_75t_R FILLER_50_705 ();
 FILLER_ASAP7_75t_R FILLER_50_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_721 ();
 DECAPx10_ASAP7_75t_R FILLER_50_732 ();
 DECAPx2_ASAP7_75t_R FILLER_50_754 ();
 FILLER_ASAP7_75t_R FILLER_50_760 ();
 DECAPx10_ASAP7_75t_R FILLER_50_768 ();
 DECAPx10_ASAP7_75t_R FILLER_50_790 ();
 DECAPx10_ASAP7_75t_R FILLER_50_812 ();
 DECAPx2_ASAP7_75t_R FILLER_50_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_840 ();
 DECAPx4_ASAP7_75t_R FILLER_50_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_881 ();
 DECAPx10_ASAP7_75t_R FILLER_50_890 ();
 DECAPx2_ASAP7_75t_R FILLER_50_912 ();
 FILLER_ASAP7_75t_R FILLER_50_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_920 ();
 DECAPx2_ASAP7_75t_R FILLER_50_933 ();
 FILLER_ASAP7_75t_R FILLER_50_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_941 ();
 DECAPx1_ASAP7_75t_R FILLER_50_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_991 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1079 ();
 FILLER_ASAP7_75t_R FILLER_50_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1191 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1241 ();
 FILLER_ASAP7_75t_R FILLER_50_1263 ();
 DECAPx4_ASAP7_75t_R FILLER_50_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_51_2 ();
 DECAPx2_ASAP7_75t_R FILLER_51_24 ();
 FILLER_ASAP7_75t_R FILLER_51_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_67 ();
 DECAPx6_ASAP7_75t_R FILLER_51_76 ();
 FILLER_ASAP7_75t_R FILLER_51_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_98 ();
 DECAPx2_ASAP7_75t_R FILLER_51_106 ();
 DECAPx1_ASAP7_75t_R FILLER_51_115 ();
 DECAPx10_ASAP7_75t_R FILLER_51_126 ();
 DECAPx6_ASAP7_75t_R FILLER_51_148 ();
 DECAPx2_ASAP7_75t_R FILLER_51_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_182 ();
 FILLER_ASAP7_75t_R FILLER_51_201 ();
 DECAPx2_ASAP7_75t_R FILLER_51_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_222 ();
 DECAPx4_ASAP7_75t_R FILLER_51_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_240 ();
 DECAPx4_ASAP7_75t_R FILLER_51_247 ();
 FILLER_ASAP7_75t_R FILLER_51_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_259 ();
 FILLER_ASAP7_75t_R FILLER_51_303 ();
 DECAPx6_ASAP7_75t_R FILLER_51_311 ();
 FILLER_ASAP7_75t_R FILLER_51_325 ();
 DECAPx4_ASAP7_75t_R FILLER_51_342 ();
 FILLER_ASAP7_75t_R FILLER_51_352 ();
 DECAPx4_ASAP7_75t_R FILLER_51_403 ();
 FILLER_ASAP7_75t_R FILLER_51_413 ();
 FILLER_ASAP7_75t_R FILLER_51_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_423 ();
 DECAPx6_ASAP7_75t_R FILLER_51_430 ();
 DECAPx1_ASAP7_75t_R FILLER_51_444 ();
 DECAPx2_ASAP7_75t_R FILLER_51_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_466 ();
 DECAPx6_ASAP7_75t_R FILLER_51_473 ();
 DECAPx1_ASAP7_75t_R FILLER_51_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_491 ();
 DECAPx4_ASAP7_75t_R FILLER_51_510 ();
 FILLER_ASAP7_75t_R FILLER_51_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_538 ();
 DECAPx6_ASAP7_75t_R FILLER_51_553 ();
 FILLER_ASAP7_75t_R FILLER_51_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_569 ();
 DECAPx10_ASAP7_75t_R FILLER_51_576 ();
 DECAPx10_ASAP7_75t_R FILLER_51_598 ();
 DECAPx10_ASAP7_75t_R FILLER_51_620 ();
 DECAPx4_ASAP7_75t_R FILLER_51_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_652 ();
 DECAPx1_ASAP7_75t_R FILLER_51_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_663 ();
 DECAPx10_ASAP7_75t_R FILLER_51_674 ();
 DECAPx10_ASAP7_75t_R FILLER_51_696 ();
 DECAPx1_ASAP7_75t_R FILLER_51_718 ();
 DECAPx10_ASAP7_75t_R FILLER_51_736 ();
 DECAPx6_ASAP7_75t_R FILLER_51_758 ();
 DECAPx1_ASAP7_75t_R FILLER_51_772 ();
 DECAPx6_ASAP7_75t_R FILLER_51_786 ();
 DECAPx2_ASAP7_75t_R FILLER_51_800 ();
 DECAPx1_ASAP7_75t_R FILLER_51_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_819 ();
 DECAPx6_ASAP7_75t_R FILLER_51_826 ();
 DECAPx1_ASAP7_75t_R FILLER_51_840 ();
 DECAPx6_ASAP7_75t_R FILLER_51_850 ();
 DECAPx10_ASAP7_75t_R FILLER_51_871 ();
 DECAPx4_ASAP7_75t_R FILLER_51_893 ();
 FILLER_ASAP7_75t_R FILLER_51_903 ();
 DECAPx4_ASAP7_75t_R FILLER_51_911 ();
 FILLER_ASAP7_75t_R FILLER_51_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_923 ();
 DECAPx1_ASAP7_75t_R FILLER_51_926 ();
 DECAPx10_ASAP7_75t_R FILLER_51_951 ();
 DECAPx1_ASAP7_75t_R FILLER_51_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_996 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1050 ();
 FILLER_ASAP7_75t_R FILLER_51_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1107 ();
 FILLER_ASAP7_75t_R FILLER_51_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_51_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1200 ();
 FILLER_ASAP7_75t_R FILLER_51_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1229 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_51_1277 ();
 FILLER_ASAP7_75t_R FILLER_51_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_52_2 ();
 DECAPx1_ASAP7_75t_R FILLER_52_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_20 ();
 DECAPx1_ASAP7_75t_R FILLER_52_36 ();
 DECAPx2_ASAP7_75t_R FILLER_52_50 ();
 FILLER_ASAP7_75t_R FILLER_52_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_58 ();
 DECAPx2_ASAP7_75t_R FILLER_52_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_88 ();
 DECAPx4_ASAP7_75t_R FILLER_52_95 ();
 FILLER_ASAP7_75t_R FILLER_52_108 ();
 DECAPx1_ASAP7_75t_R FILLER_52_154 ();
 DECAPx6_ASAP7_75t_R FILLER_52_164 ();
 FILLER_ASAP7_75t_R FILLER_52_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_180 ();
 DECAPx2_ASAP7_75t_R FILLER_52_193 ();
 FILLER_ASAP7_75t_R FILLER_52_199 ();
 FILLER_ASAP7_75t_R FILLER_52_207 ();
 DECAPx6_ASAP7_75t_R FILLER_52_223 ();
 FILLER_ASAP7_75t_R FILLER_52_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_239 ();
 DECAPx4_ASAP7_75t_R FILLER_52_256 ();
 DECAPx2_ASAP7_75t_R FILLER_52_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_279 ();
 FILLER_ASAP7_75t_R FILLER_52_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_288 ();
 FILLER_ASAP7_75t_R FILLER_52_297 ();
 DECAPx10_ASAP7_75t_R FILLER_52_307 ();
 DECAPx4_ASAP7_75t_R FILLER_52_329 ();
 FILLER_ASAP7_75t_R FILLER_52_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_358 ();
 DECAPx2_ASAP7_75t_R FILLER_52_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_375 ();
 DECAPx2_ASAP7_75t_R FILLER_52_392 ();
 FILLER_ASAP7_75t_R FILLER_52_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_400 ();
 DECAPx1_ASAP7_75t_R FILLER_52_411 ();
 DECAPx4_ASAP7_75t_R FILLER_52_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_439 ();
 FILLER_ASAP7_75t_R FILLER_52_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_461 ();
 DECAPx10_ASAP7_75t_R FILLER_52_464 ();
 DECAPx4_ASAP7_75t_R FILLER_52_486 ();
 FILLER_ASAP7_75t_R FILLER_52_496 ();
 FILLER_ASAP7_75t_R FILLER_52_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_535 ();
 FILLER_ASAP7_75t_R FILLER_52_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_544 ();
 DECAPx4_ASAP7_75t_R FILLER_52_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_585 ();
 FILLER_ASAP7_75t_R FILLER_52_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_598 ();
 FILLER_ASAP7_75t_R FILLER_52_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_611 ();
 DECAPx2_ASAP7_75t_R FILLER_52_620 ();
 DECAPx2_ASAP7_75t_R FILLER_52_641 ();
 FILLER_ASAP7_75t_R FILLER_52_647 ();
 DECAPx10_ASAP7_75t_R FILLER_52_655 ();
 DECAPx2_ASAP7_75t_R FILLER_52_677 ();
 FILLER_ASAP7_75t_R FILLER_52_683 ();
 DECAPx10_ASAP7_75t_R FILLER_52_695 ();
 DECAPx10_ASAP7_75t_R FILLER_52_717 ();
 DECAPx1_ASAP7_75t_R FILLER_52_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_743 ();
 DECAPx1_ASAP7_75t_R FILLER_52_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_756 ();
 DECAPx10_ASAP7_75t_R FILLER_52_767 ();
 DECAPx6_ASAP7_75t_R FILLER_52_789 ();
 DECAPx4_ASAP7_75t_R FILLER_52_812 ();
 FILLER_ASAP7_75t_R FILLER_52_822 ();
 DECAPx2_ASAP7_75t_R FILLER_52_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_842 ();
 DECAPx4_ASAP7_75t_R FILLER_52_851 ();
 DECAPx6_ASAP7_75t_R FILLER_52_882 ();
 DECAPx2_ASAP7_75t_R FILLER_52_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_902 ();
 DECAPx6_ASAP7_75t_R FILLER_52_909 ();
 FILLER_ASAP7_75t_R FILLER_52_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_925 ();
 DECAPx6_ASAP7_75t_R FILLER_52_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_946 ();
 DECAPx4_ASAP7_75t_R FILLER_52_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_960 ();
 DECAPx10_ASAP7_75t_R FILLER_52_981 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1003 ();
 FILLER_ASAP7_75t_R FILLER_52_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1068 ();
 FILLER_ASAP7_75t_R FILLER_52_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1200 ();
 FILLER_ASAP7_75t_R FILLER_52_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_53_2 ();
 FILLER_ASAP7_75t_R FILLER_53_16 ();
 DECAPx2_ASAP7_75t_R FILLER_53_47 ();
 FILLER_ASAP7_75t_R FILLER_53_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_55 ();
 DECAPx2_ASAP7_75t_R FILLER_53_79 ();
 FILLER_ASAP7_75t_R FILLER_53_85 ();
 DECAPx1_ASAP7_75t_R FILLER_53_93 ();
 FILLER_ASAP7_75t_R FILLER_53_112 ();
 DECAPx1_ASAP7_75t_R FILLER_53_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_133 ();
 FILLER_ASAP7_75t_R FILLER_53_137 ();
 DECAPx2_ASAP7_75t_R FILLER_53_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_154 ();
 FILLER_ASAP7_75t_R FILLER_53_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_177 ();
 DECAPx6_ASAP7_75t_R FILLER_53_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_204 ();
 FILLER_ASAP7_75t_R FILLER_53_213 ();
 DECAPx4_ASAP7_75t_R FILLER_53_222 ();
 FILLER_ASAP7_75t_R FILLER_53_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_234 ();
 DECAPx2_ASAP7_75t_R FILLER_53_252 ();
 FILLER_ASAP7_75t_R FILLER_53_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_267 ();
 FILLER_ASAP7_75t_R FILLER_53_271 ();
 FILLER_ASAP7_75t_R FILLER_53_276 ();
 DECAPx2_ASAP7_75t_R FILLER_53_295 ();
 FILLER_ASAP7_75t_R FILLER_53_301 ();
 DECAPx2_ASAP7_75t_R FILLER_53_309 ();
 FILLER_ASAP7_75t_R FILLER_53_315 ();
 DECAPx4_ASAP7_75t_R FILLER_53_333 ();
 FILLER_ASAP7_75t_R FILLER_53_343 ();
 DECAPx2_ASAP7_75t_R FILLER_53_366 ();
 FILLER_ASAP7_75t_R FILLER_53_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_382 ();
 DECAPx1_ASAP7_75t_R FILLER_53_393 ();
 DECAPx6_ASAP7_75t_R FILLER_53_404 ();
 DECAPx1_ASAP7_75t_R FILLER_53_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_422 ();
 DECAPx10_ASAP7_75t_R FILLER_53_435 ();
 DECAPx2_ASAP7_75t_R FILLER_53_457 ();
 FILLER_ASAP7_75t_R FILLER_53_463 ();
 DECAPx2_ASAP7_75t_R FILLER_53_471 ();
 FILLER_ASAP7_75t_R FILLER_53_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_479 ();
 DECAPx1_ASAP7_75t_R FILLER_53_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_496 ();
 DECAPx2_ASAP7_75t_R FILLER_53_515 ();
 DECAPx2_ASAP7_75t_R FILLER_53_527 ();
 FILLER_ASAP7_75t_R FILLER_53_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_535 ();
 DECAPx2_ASAP7_75t_R FILLER_53_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_558 ();
 DECAPx1_ASAP7_75t_R FILLER_53_567 ();
 DECAPx2_ASAP7_75t_R FILLER_53_577 ();
 DECAPx2_ASAP7_75t_R FILLER_53_589 ();
 FILLER_ASAP7_75t_R FILLER_53_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_632 ();
 DECAPx10_ASAP7_75t_R FILLER_53_640 ();
 DECAPx10_ASAP7_75t_R FILLER_53_662 ();
 DECAPx10_ASAP7_75t_R FILLER_53_684 ();
 DECAPx2_ASAP7_75t_R FILLER_53_706 ();
 FILLER_ASAP7_75t_R FILLER_53_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_714 ();
 FILLER_ASAP7_75t_R FILLER_53_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_730 ();
 DECAPx6_ASAP7_75t_R FILLER_53_741 ();
 DECAPx2_ASAP7_75t_R FILLER_53_755 ();
 DECAPx10_ASAP7_75t_R FILLER_53_767 ();
 DECAPx10_ASAP7_75t_R FILLER_53_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_811 ();
 DECAPx10_ASAP7_75t_R FILLER_53_832 ();
 DECAPx10_ASAP7_75t_R FILLER_53_854 ();
 DECAPx10_ASAP7_75t_R FILLER_53_876 ();
 FILLER_ASAP7_75t_R FILLER_53_898 ();
 FILLER_ASAP7_75t_R FILLER_53_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_912 ();
 DECAPx1_ASAP7_75t_R FILLER_53_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_926 ();
 DECAPx2_ASAP7_75t_R FILLER_53_934 ();
 FILLER_ASAP7_75t_R FILLER_53_940 ();
 DECAPx4_ASAP7_75t_R FILLER_53_960 ();
 DECAPx10_ASAP7_75t_R FILLER_53_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1017 ();
 FILLER_ASAP7_75t_R FILLER_53_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1227 ();
 FILLER_ASAP7_75t_R FILLER_53_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1241 ();
 FILLER_ASAP7_75t_R FILLER_53_1251 ();
 FILLER_ASAP7_75t_R FILLER_53_1263 ();
 DECAPx4_ASAP7_75t_R FILLER_54_2 ();
 FILLER_ASAP7_75t_R FILLER_54_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_14 ();
 FILLER_ASAP7_75t_R FILLER_54_28 ();
 FILLER_ASAP7_75t_R FILLER_54_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_46 ();
 DECAPx2_ASAP7_75t_R FILLER_54_59 ();
 DECAPx6_ASAP7_75t_R FILLER_54_77 ();
 DECAPx2_ASAP7_75t_R FILLER_54_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_107 ();
 FILLER_ASAP7_75t_R FILLER_54_124 ();
 DECAPx2_ASAP7_75t_R FILLER_54_144 ();
 FILLER_ASAP7_75t_R FILLER_54_150 ();
 FILLER_ASAP7_75t_R FILLER_54_172 ();
 DECAPx2_ASAP7_75t_R FILLER_54_185 ();
 FILLER_ASAP7_75t_R FILLER_54_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_193 ();
 DECAPx1_ASAP7_75t_R FILLER_54_208 ();
 FILLER_ASAP7_75t_R FILLER_54_218 ();
 FILLER_ASAP7_75t_R FILLER_54_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_238 ();
 FILLER_ASAP7_75t_R FILLER_54_246 ();
 FILLER_ASAP7_75t_R FILLER_54_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_256 ();
 FILLER_ASAP7_75t_R FILLER_54_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_267 ();
 FILLER_ASAP7_75t_R FILLER_54_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_276 ();
 DECAPx2_ASAP7_75t_R FILLER_54_289 ();
 FILLER_ASAP7_75t_R FILLER_54_295 ();
 DECAPx2_ASAP7_75t_R FILLER_54_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_315 ();
 DECAPx6_ASAP7_75t_R FILLER_54_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_342 ();
 DECAPx1_ASAP7_75t_R FILLER_54_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_376 ();
 DECAPx4_ASAP7_75t_R FILLER_54_419 ();
 FILLER_ASAP7_75t_R FILLER_54_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_437 ();
 DECAPx1_ASAP7_75t_R FILLER_54_452 ();
 FILLER_ASAP7_75t_R FILLER_54_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_461 ();
 DECAPx6_ASAP7_75t_R FILLER_54_464 ();
 DECAPx2_ASAP7_75t_R FILLER_54_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_484 ();
 DECAPx6_ASAP7_75t_R FILLER_54_497 ();
 DECAPx2_ASAP7_75t_R FILLER_54_511 ();
 FILLER_ASAP7_75t_R FILLER_54_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_533 ();
 DECAPx6_ASAP7_75t_R FILLER_54_541 ();
 DECAPx2_ASAP7_75t_R FILLER_54_565 ();
 FILLER_ASAP7_75t_R FILLER_54_571 ();
 DECAPx10_ASAP7_75t_R FILLER_54_583 ();
 DECAPx10_ASAP7_75t_R FILLER_54_605 ();
 DECAPx10_ASAP7_75t_R FILLER_54_627 ();
 DECAPx6_ASAP7_75t_R FILLER_54_649 ();
 FILLER_ASAP7_75t_R FILLER_54_663 ();
 DECAPx6_ASAP7_75t_R FILLER_54_680 ();
 FILLER_ASAP7_75t_R FILLER_54_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_696 ();
 DECAPx4_ASAP7_75t_R FILLER_54_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_717 ();
 DECAPx10_ASAP7_75t_R FILLER_54_730 ();
 DECAPx2_ASAP7_75t_R FILLER_54_752 ();
 FILLER_ASAP7_75t_R FILLER_54_758 ();
 FILLER_ASAP7_75t_R FILLER_54_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_768 ();
 DECAPx1_ASAP7_75t_R FILLER_54_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_794 ();
 DECAPx6_ASAP7_75t_R FILLER_54_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_819 ();
 DECAPx10_ASAP7_75t_R FILLER_54_826 ();
 DECAPx6_ASAP7_75t_R FILLER_54_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_862 ();
 DECAPx1_ASAP7_75t_R FILLER_54_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_877 ();
 DECAPx1_ASAP7_75t_R FILLER_54_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_885 ();
 DECAPx6_ASAP7_75t_R FILLER_54_898 ();
 FILLER_ASAP7_75t_R FILLER_54_912 ();
 DECAPx2_ASAP7_75t_R FILLER_54_922 ();
 FILLER_ASAP7_75t_R FILLER_54_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_930 ();
 DECAPx6_ASAP7_75t_R FILLER_54_939 ();
 DECAPx1_ASAP7_75t_R FILLER_54_953 ();
 DECAPx10_ASAP7_75t_R FILLER_54_965 ();
 DECAPx4_ASAP7_75t_R FILLER_54_987 ();
 FILLER_ASAP7_75t_R FILLER_54_997 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_54_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1158 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1181 ();
 FILLER_ASAP7_75t_R FILLER_54_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1247 ();
 FILLER_ASAP7_75t_R FILLER_54_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_55_2 ();
 FILLER_ASAP7_75t_R FILLER_55_8 ();
 FILLER_ASAP7_75t_R FILLER_55_23 ();
 FILLER_ASAP7_75t_R FILLER_55_33 ();
 FILLER_ASAP7_75t_R FILLER_55_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_43 ();
 DECAPx10_ASAP7_75t_R FILLER_55_56 ();
 DECAPx1_ASAP7_75t_R FILLER_55_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_98 ();
 FILLER_ASAP7_75t_R FILLER_55_119 ();
 DECAPx1_ASAP7_75t_R FILLER_55_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_148 ();
 FILLER_ASAP7_75t_R FILLER_55_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_193 ();
 DECAPx4_ASAP7_75t_R FILLER_55_201 ();
 FILLER_ASAP7_75t_R FILLER_55_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_213 ();
 FILLER_ASAP7_75t_R FILLER_55_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_277 ();
 DECAPx1_ASAP7_75t_R FILLER_55_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_288 ();
 DECAPx1_ASAP7_75t_R FILLER_55_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_301 ();
 DECAPx10_ASAP7_75t_R FILLER_55_312 ();
 DECAPx6_ASAP7_75t_R FILLER_55_334 ();
 FILLER_ASAP7_75t_R FILLER_55_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_350 ();
 DECAPx4_ASAP7_75t_R FILLER_55_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_378 ();
 DECAPx4_ASAP7_75t_R FILLER_55_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_406 ();
 DECAPx6_ASAP7_75t_R FILLER_55_415 ();
 DECAPx1_ASAP7_75t_R FILLER_55_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_433 ();
 DECAPx4_ASAP7_75t_R FILLER_55_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_453 ();
 DECAPx4_ASAP7_75t_R FILLER_55_475 ();
 FILLER_ASAP7_75t_R FILLER_55_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_487 ();
 DECAPx6_ASAP7_75t_R FILLER_55_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_508 ();
 DECAPx1_ASAP7_75t_R FILLER_55_531 ();
 DECAPx10_ASAP7_75t_R FILLER_55_556 ();
 DECAPx6_ASAP7_75t_R FILLER_55_578 ();
 DECAPx2_ASAP7_75t_R FILLER_55_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_598 ();
 DECAPx6_ASAP7_75t_R FILLER_55_605 ();
 DECAPx2_ASAP7_75t_R FILLER_55_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_625 ();
 DECAPx6_ASAP7_75t_R FILLER_55_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_646 ();
 DECAPx6_ASAP7_75t_R FILLER_55_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_688 ();
 DECAPx6_ASAP7_75t_R FILLER_55_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_713 ();
 DECAPx6_ASAP7_75t_R FILLER_55_728 ();
 FILLER_ASAP7_75t_R FILLER_55_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_744 ();
 DECAPx1_ASAP7_75t_R FILLER_55_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_771 ();
 DECAPx2_ASAP7_75t_R FILLER_55_784 ();
 DECAPx10_ASAP7_75t_R FILLER_55_796 ();
 DECAPx2_ASAP7_75t_R FILLER_55_818 ();
 DECAPx10_ASAP7_75t_R FILLER_55_832 ();
 FILLER_ASAP7_75t_R FILLER_55_854 ();
 DECAPx10_ASAP7_75t_R FILLER_55_862 ();
 DECAPx10_ASAP7_75t_R FILLER_55_884 ();
 DECAPx6_ASAP7_75t_R FILLER_55_906 ();
 DECAPx1_ASAP7_75t_R FILLER_55_920 ();
 DECAPx1_ASAP7_75t_R FILLER_55_926 ();
 DECAPx10_ASAP7_75t_R FILLER_55_940 ();
 DECAPx2_ASAP7_75t_R FILLER_55_962 ();
 FILLER_ASAP7_75t_R FILLER_55_968 ();
 DECAPx10_ASAP7_75t_R FILLER_55_978 ();
 FILLER_ASAP7_75t_R FILLER_55_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_55_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1140 ();
 FILLER_ASAP7_75t_R FILLER_55_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1155 ();
 FILLER_ASAP7_75t_R FILLER_55_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_56_2 ();
 FILLER_ASAP7_75t_R FILLER_56_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_14 ();
 DECAPx1_ASAP7_75t_R FILLER_56_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_26 ();
 FILLER_ASAP7_75t_R FILLER_56_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_43 ();
 DECAPx4_ASAP7_75t_R FILLER_56_56 ();
 FILLER_ASAP7_75t_R FILLER_56_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_68 ();
 DECAPx6_ASAP7_75t_R FILLER_56_72 ();
 DECAPx1_ASAP7_75t_R FILLER_56_86 ();
 FILLER_ASAP7_75t_R FILLER_56_116 ();
 DECAPx6_ASAP7_75t_R FILLER_56_134 ();
 DECAPx4_ASAP7_75t_R FILLER_56_160 ();
 FILLER_ASAP7_75t_R FILLER_56_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_172 ();
 DECAPx1_ASAP7_75t_R FILLER_56_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_189 ();
 DECAPx1_ASAP7_75t_R FILLER_56_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_213 ();
 DECAPx2_ASAP7_75t_R FILLER_56_220 ();
 FILLER_ASAP7_75t_R FILLER_56_226 ();
 DECAPx2_ASAP7_75t_R FILLER_56_234 ();
 DECAPx1_ASAP7_75t_R FILLER_56_258 ();
 DECAPx2_ASAP7_75t_R FILLER_56_269 ();
 FILLER_ASAP7_75t_R FILLER_56_301 ();
 DECAPx6_ASAP7_75t_R FILLER_56_313 ();
 DECAPx1_ASAP7_75t_R FILLER_56_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_331 ();
 DECAPx6_ASAP7_75t_R FILLER_56_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_356 ();
 DECAPx10_ASAP7_75t_R FILLER_56_367 ();
 FILLER_ASAP7_75t_R FILLER_56_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_391 ();
 DECAPx4_ASAP7_75t_R FILLER_56_398 ();
 DECAPx6_ASAP7_75t_R FILLER_56_414 ();
 DECAPx1_ASAP7_75t_R FILLER_56_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_432 ();
 DECAPx4_ASAP7_75t_R FILLER_56_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_449 ();
 DECAPx1_ASAP7_75t_R FILLER_56_464 ();
 DECAPx10_ASAP7_75t_R FILLER_56_496 ();
 DECAPx2_ASAP7_75t_R FILLER_56_518 ();
 FILLER_ASAP7_75t_R FILLER_56_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_526 ();
 DECAPx10_ASAP7_75t_R FILLER_56_533 ();
 DECAPx6_ASAP7_75t_R FILLER_56_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_569 ();
 DECAPx10_ASAP7_75t_R FILLER_56_576 ();
 DECAPx2_ASAP7_75t_R FILLER_56_598 ();
 DECAPx2_ASAP7_75t_R FILLER_56_634 ();
 FILLER_ASAP7_75t_R FILLER_56_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_648 ();
 DECAPx1_ASAP7_75t_R FILLER_56_655 ();
 DECAPx4_ASAP7_75t_R FILLER_56_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_685 ();
 DECAPx4_ASAP7_75t_R FILLER_56_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_699 ();
 DECAPx10_ASAP7_75t_R FILLER_56_710 ();
 DECAPx6_ASAP7_75t_R FILLER_56_732 ();
 FILLER_ASAP7_75t_R FILLER_56_746 ();
 DECAPx1_ASAP7_75t_R FILLER_56_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_758 ();
 FILLER_ASAP7_75t_R FILLER_56_783 ();
 DECAPx10_ASAP7_75t_R FILLER_56_791 ();
 DECAPx1_ASAP7_75t_R FILLER_56_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_817 ();
 DECAPx4_ASAP7_75t_R FILLER_56_834 ();
 FILLER_ASAP7_75t_R FILLER_56_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_854 ();
 DECAPx10_ASAP7_75t_R FILLER_56_871 ();
 DECAPx2_ASAP7_75t_R FILLER_56_893 ();
 FILLER_ASAP7_75t_R FILLER_56_899 ();
 DECAPx1_ASAP7_75t_R FILLER_56_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_918 ();
 DECAPx10_ASAP7_75t_R FILLER_56_935 ();
 DECAPx10_ASAP7_75t_R FILLER_56_957 ();
 DECAPx1_ASAP7_75t_R FILLER_56_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_983 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1028 ();
 FILLER_ASAP7_75t_R FILLER_56_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1052 ();
 FILLER_ASAP7_75t_R FILLER_56_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1091 ();
 FILLER_ASAP7_75t_R FILLER_56_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1128 ();
 FILLER_ASAP7_75t_R FILLER_56_1149 ();
 FILLER_ASAP7_75t_R FILLER_56_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_56_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1276 ();
 FILLER_ASAP7_75t_R FILLER_56_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_57_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_8 ();
 DECAPx4_ASAP7_75t_R FILLER_57_16 ();
 FILLER_ASAP7_75t_R FILLER_57_26 ();
 DECAPx2_ASAP7_75t_R FILLER_57_35 ();
 FILLER_ASAP7_75t_R FILLER_57_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_43 ();
 FILLER_ASAP7_75t_R FILLER_57_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_52 ();
 DECAPx4_ASAP7_75t_R FILLER_57_77 ();
 FILLER_ASAP7_75t_R FILLER_57_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_89 ();
 DECAPx4_ASAP7_75t_R FILLER_57_111 ();
 FILLER_ASAP7_75t_R FILLER_57_121 ();
 FILLER_ASAP7_75t_R FILLER_57_129 ();
 DECAPx10_ASAP7_75t_R FILLER_57_138 ();
 DECAPx2_ASAP7_75t_R FILLER_57_160 ();
 FILLER_ASAP7_75t_R FILLER_57_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_168 ();
 DECAPx4_ASAP7_75t_R FILLER_57_180 ();
 FILLER_ASAP7_75t_R FILLER_57_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_192 ();
 DECAPx2_ASAP7_75t_R FILLER_57_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_207 ();
 DECAPx1_ASAP7_75t_R FILLER_57_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_220 ();
 DECAPx1_ASAP7_75t_R FILLER_57_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_231 ();
 DECAPx1_ASAP7_75t_R FILLER_57_238 ();
 DECAPx1_ASAP7_75t_R FILLER_57_258 ();
 DECAPx2_ASAP7_75t_R FILLER_57_271 ();
 FILLER_ASAP7_75t_R FILLER_57_277 ();
 DECAPx1_ASAP7_75t_R FILLER_57_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_358 ();
 DECAPx2_ASAP7_75t_R FILLER_57_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_372 ();
 DECAPx4_ASAP7_75t_R FILLER_57_383 ();
 DECAPx2_ASAP7_75t_R FILLER_57_415 ();
 FILLER_ASAP7_75t_R FILLER_57_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_423 ();
 FILLER_ASAP7_75t_R FILLER_57_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_441 ();
 DECAPx6_ASAP7_75t_R FILLER_57_454 ();
 FILLER_ASAP7_75t_R FILLER_57_474 ();
 DECAPx6_ASAP7_75t_R FILLER_57_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_510 ();
 DECAPx2_ASAP7_75t_R FILLER_57_521 ();
 DECAPx6_ASAP7_75t_R FILLER_57_538 ();
 DECAPx1_ASAP7_75t_R FILLER_57_552 ();
 DECAPx2_ASAP7_75t_R FILLER_57_566 ();
 DECAPx6_ASAP7_75t_R FILLER_57_578 ();
 DECAPx10_ASAP7_75t_R FILLER_57_606 ();
 DECAPx6_ASAP7_75t_R FILLER_57_628 ();
 FILLER_ASAP7_75t_R FILLER_57_642 ();
 DECAPx1_ASAP7_75t_R FILLER_57_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_667 ();
 DECAPx6_ASAP7_75t_R FILLER_57_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_702 ();
 DECAPx6_ASAP7_75t_R FILLER_57_713 ();
 DECAPx10_ASAP7_75t_R FILLER_57_759 ();
 DECAPx10_ASAP7_75t_R FILLER_57_781 ();
 DECAPx10_ASAP7_75t_R FILLER_57_803 ();
 DECAPx10_ASAP7_75t_R FILLER_57_825 ();
 DECAPx2_ASAP7_75t_R FILLER_57_847 ();
 FILLER_ASAP7_75t_R FILLER_57_853 ();
 DECAPx2_ASAP7_75t_R FILLER_57_895 ();
 FILLER_ASAP7_75t_R FILLER_57_901 ();
 DECAPx6_ASAP7_75t_R FILLER_57_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_923 ();
 DECAPx10_ASAP7_75t_R FILLER_57_926 ();
 DECAPx10_ASAP7_75t_R FILLER_57_948 ();
 DECAPx10_ASAP7_75t_R FILLER_57_970 ();
 DECAPx10_ASAP7_75t_R FILLER_57_992 ();
 FILLER_ASAP7_75t_R FILLER_57_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1106 ();
 FILLER_ASAP7_75t_R FILLER_57_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1210 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_58_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_22 ();
 FILLER_ASAP7_75t_R FILLER_58_80 ();
 DECAPx1_ASAP7_75t_R FILLER_58_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_116 ();
 DECAPx1_ASAP7_75t_R FILLER_58_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_128 ();
 FILLER_ASAP7_75t_R FILLER_58_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_146 ();
 FILLER_ASAP7_75t_R FILLER_58_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_180 ();
 DECAPx4_ASAP7_75t_R FILLER_58_188 ();
 DECAPx4_ASAP7_75t_R FILLER_58_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_211 ();
 DECAPx4_ASAP7_75t_R FILLER_58_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_260 ();
 DECAPx2_ASAP7_75t_R FILLER_58_267 ();
 DECAPx10_ASAP7_75t_R FILLER_58_291 ();
 FILLER_ASAP7_75t_R FILLER_58_313 ();
 DECAPx2_ASAP7_75t_R FILLER_58_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_332 ();
 DECAPx4_ASAP7_75t_R FILLER_58_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_357 ();
 DECAPx10_ASAP7_75t_R FILLER_58_379 ();
 DECAPx6_ASAP7_75t_R FILLER_58_401 ();
 DECAPx2_ASAP7_75t_R FILLER_58_415 ();
 DECAPx6_ASAP7_75t_R FILLER_58_439 ();
 FILLER_ASAP7_75t_R FILLER_58_453 ();
 DECAPx6_ASAP7_75t_R FILLER_58_464 ();
 FILLER_ASAP7_75t_R FILLER_58_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_480 ();
 FILLER_ASAP7_75t_R FILLER_58_528 ();
 DECAPx4_ASAP7_75t_R FILLER_58_542 ();
 FILLER_ASAP7_75t_R FILLER_58_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_554 ();
 DECAPx10_ASAP7_75t_R FILLER_58_616 ();
 DECAPx2_ASAP7_75t_R FILLER_58_638 ();
 FILLER_ASAP7_75t_R FILLER_58_644 ();
 DECAPx10_ASAP7_75t_R FILLER_58_654 ();
 DECAPx10_ASAP7_75t_R FILLER_58_676 ();
 DECAPx10_ASAP7_75t_R FILLER_58_698 ();
 DECAPx2_ASAP7_75t_R FILLER_58_720 ();
 FILLER_ASAP7_75t_R FILLER_58_726 ();
 DECAPx4_ASAP7_75t_R FILLER_58_736 ();
 FILLER_ASAP7_75t_R FILLER_58_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_748 ();
 FILLER_ASAP7_75t_R FILLER_58_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_757 ();
 DECAPx6_ASAP7_75t_R FILLER_58_764 ();
 DECAPx1_ASAP7_75t_R FILLER_58_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_782 ();
 DECAPx4_ASAP7_75t_R FILLER_58_793 ();
 FILLER_ASAP7_75t_R FILLER_58_803 ();
 DECAPx10_ASAP7_75t_R FILLER_58_811 ();
 DECAPx10_ASAP7_75t_R FILLER_58_833 ();
 DECAPx2_ASAP7_75t_R FILLER_58_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_861 ();
 DECAPx6_ASAP7_75t_R FILLER_58_869 ();
 DECAPx2_ASAP7_75t_R FILLER_58_883 ();
 DECAPx6_ASAP7_75t_R FILLER_58_895 ();
 DECAPx2_ASAP7_75t_R FILLER_58_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_915 ();
 DECAPx4_ASAP7_75t_R FILLER_58_922 ();
 DECAPx10_ASAP7_75t_R FILLER_58_944 ();
 DECAPx10_ASAP7_75t_R FILLER_58_966 ();
 FILLER_ASAP7_75t_R FILLER_58_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_990 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1001 ();
 FILLER_ASAP7_75t_R FILLER_58_1007 ();
 FILLER_ASAP7_75t_R FILLER_58_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1052 ();
 FILLER_ASAP7_75t_R FILLER_58_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_58_1076 ();
 FILLER_ASAP7_75t_R FILLER_58_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_58_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1182 ();
 FILLER_ASAP7_75t_R FILLER_58_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_59_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_23 ();
 DECAPx2_ASAP7_75t_R FILLER_59_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_63 ();
 DECAPx6_ASAP7_75t_R FILLER_59_67 ();
 DECAPx10_ASAP7_75t_R FILLER_59_87 ();
 DECAPx2_ASAP7_75t_R FILLER_59_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_115 ();
 FILLER_ASAP7_75t_R FILLER_59_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_127 ();
 DECAPx2_ASAP7_75t_R FILLER_59_135 ();
 FILLER_ASAP7_75t_R FILLER_59_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_152 ();
 DECAPx2_ASAP7_75t_R FILLER_59_162 ();
 FILLER_ASAP7_75t_R FILLER_59_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_170 ();
 FILLER_ASAP7_75t_R FILLER_59_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_197 ();
 FILLER_ASAP7_75t_R FILLER_59_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_213 ();
 DECAPx10_ASAP7_75t_R FILLER_59_225 ();
 DECAPx10_ASAP7_75t_R FILLER_59_247 ();
 DECAPx1_ASAP7_75t_R FILLER_59_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_273 ();
 DECAPx10_ASAP7_75t_R FILLER_59_284 ();
 DECAPx1_ASAP7_75t_R FILLER_59_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_310 ();
 DECAPx6_ASAP7_75t_R FILLER_59_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_339 ();
 DECAPx10_ASAP7_75t_R FILLER_59_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_372 ();
 DECAPx6_ASAP7_75t_R FILLER_59_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_424 ();
 DECAPx10_ASAP7_75t_R FILLER_59_442 ();
 DECAPx6_ASAP7_75t_R FILLER_59_464 ();
 FILLER_ASAP7_75t_R FILLER_59_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_525 ();
 DECAPx1_ASAP7_75t_R FILLER_59_538 ();
 DECAPx6_ASAP7_75t_R FILLER_59_549 ();
 FILLER_ASAP7_75t_R FILLER_59_563 ();
 DECAPx6_ASAP7_75t_R FILLER_59_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_609 ();
 DECAPx10_ASAP7_75t_R FILLER_59_616 ();
 DECAPx6_ASAP7_75t_R FILLER_59_638 ();
 FILLER_ASAP7_75t_R FILLER_59_652 ();
 DECAPx4_ASAP7_75t_R FILLER_59_660 ();
 FILLER_ASAP7_75t_R FILLER_59_670 ();
 DECAPx10_ASAP7_75t_R FILLER_59_678 ();
 DECAPx6_ASAP7_75t_R FILLER_59_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_714 ();
 DECAPx10_ASAP7_75t_R FILLER_59_721 ();
 FILLER_ASAP7_75t_R FILLER_59_743 ();
 FILLER_ASAP7_75t_R FILLER_59_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_758 ();
 DECAPx4_ASAP7_75t_R FILLER_59_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_779 ();
 DECAPx4_ASAP7_75t_R FILLER_59_786 ();
 FILLER_ASAP7_75t_R FILLER_59_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_798 ();
 DECAPx10_ASAP7_75t_R FILLER_59_809 ();
 DECAPx10_ASAP7_75t_R FILLER_59_831 ();
 DECAPx2_ASAP7_75t_R FILLER_59_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_859 ();
 DECAPx10_ASAP7_75t_R FILLER_59_877 ();
 DECAPx2_ASAP7_75t_R FILLER_59_899 ();
 FILLER_ASAP7_75t_R FILLER_59_905 ();
 DECAPx4_ASAP7_75t_R FILLER_59_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_923 ();
 DECAPx1_ASAP7_75t_R FILLER_59_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_930 ();
 DECAPx2_ASAP7_75t_R FILLER_59_943 ();
 FILLER_ASAP7_75t_R FILLER_59_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_951 ();
 DECAPx10_ASAP7_75t_R FILLER_59_962 ();
 DECAPx2_ASAP7_75t_R FILLER_59_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_990 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1023 ();
 FILLER_ASAP7_75t_R FILLER_59_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1069 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1091 ();
 FILLER_ASAP7_75t_R FILLER_59_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1139 ();
 FILLER_ASAP7_75t_R FILLER_59_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1203 ();
 FILLER_ASAP7_75t_R FILLER_59_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_59_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_60_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_34 ();
 FILLER_ASAP7_75t_R FILLER_60_50 ();
 DECAPx1_ASAP7_75t_R FILLER_60_58 ();
 DECAPx4_ASAP7_75t_R FILLER_60_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_75 ();
 DECAPx1_ASAP7_75t_R FILLER_60_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_95 ();
 DECAPx1_ASAP7_75t_R FILLER_60_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_134 ();
 DECAPx2_ASAP7_75t_R FILLER_60_147 ();
 DECAPx6_ASAP7_75t_R FILLER_60_168 ();
 DECAPx2_ASAP7_75t_R FILLER_60_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_188 ();
 DECAPx2_ASAP7_75t_R FILLER_60_217 ();
 FILLER_ASAP7_75t_R FILLER_60_223 ();
 DECAPx6_ASAP7_75t_R FILLER_60_231 ();
 DECAPx2_ASAP7_75t_R FILLER_60_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_251 ();
 FILLER_ASAP7_75t_R FILLER_60_269 ();
 DECAPx6_ASAP7_75t_R FILLER_60_294 ();
 FILLER_ASAP7_75t_R FILLER_60_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_310 ();
 DECAPx2_ASAP7_75t_R FILLER_60_319 ();
 FILLER_ASAP7_75t_R FILLER_60_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_349 ();
 DECAPx2_ASAP7_75t_R FILLER_60_399 ();
 DECAPx10_ASAP7_75t_R FILLER_60_411 ();
 FILLER_ASAP7_75t_R FILLER_60_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_435 ();
 DECAPx4_ASAP7_75t_R FILLER_60_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_452 ();
 FILLER_ASAP7_75t_R FILLER_60_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_466 ();
 DECAPx2_ASAP7_75t_R FILLER_60_473 ();
 FILLER_ASAP7_75t_R FILLER_60_479 ();
 DECAPx6_ASAP7_75t_R FILLER_60_505 ();
 FILLER_ASAP7_75t_R FILLER_60_519 ();
 DECAPx2_ASAP7_75t_R FILLER_60_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_537 ();
 DECAPx10_ASAP7_75t_R FILLER_60_546 ();
 DECAPx4_ASAP7_75t_R FILLER_60_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_578 ();
 DECAPx10_ASAP7_75t_R FILLER_60_587 ();
 DECAPx6_ASAP7_75t_R FILLER_60_609 ();
 DECAPx1_ASAP7_75t_R FILLER_60_623 ();
 DECAPx6_ASAP7_75t_R FILLER_60_637 ();
 DECAPx1_ASAP7_75t_R FILLER_60_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_655 ();
 DECAPx1_ASAP7_75t_R FILLER_60_662 ();
 DECAPx10_ASAP7_75t_R FILLER_60_676 ();
 FILLER_ASAP7_75t_R FILLER_60_698 ();
 DECAPx2_ASAP7_75t_R FILLER_60_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_715 ();
 DECAPx10_ASAP7_75t_R FILLER_60_722 ();
 DECAPx2_ASAP7_75t_R FILLER_60_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_750 ();
 DECAPx2_ASAP7_75t_R FILLER_60_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_763 ();
 DECAPx6_ASAP7_75t_R FILLER_60_774 ();
 FILLER_ASAP7_75t_R FILLER_60_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_790 ();
 DECAPx4_ASAP7_75t_R FILLER_60_800 ();
 FILLER_ASAP7_75t_R FILLER_60_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_825 ();
 DECAPx10_ASAP7_75t_R FILLER_60_836 ();
 DECAPx10_ASAP7_75t_R FILLER_60_858 ();
 DECAPx4_ASAP7_75t_R FILLER_60_880 ();
 FILLER_ASAP7_75t_R FILLER_60_890 ();
 DECAPx10_ASAP7_75t_R FILLER_60_902 ();
 DECAPx2_ASAP7_75t_R FILLER_60_924 ();
 FILLER_ASAP7_75t_R FILLER_60_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_932 ();
 FILLER_ASAP7_75t_R FILLER_60_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_942 ();
 DECAPx10_ASAP7_75t_R FILLER_60_957 ();
 DECAPx10_ASAP7_75t_R FILLER_60_979 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1033 ();
 FILLER_ASAP7_75t_R FILLER_60_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1060 ();
 FILLER_ASAP7_75t_R FILLER_60_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1092 ();
 FILLER_ASAP7_75t_R FILLER_60_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1114 ();
 FILLER_ASAP7_75t_R FILLER_60_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1137 ();
 FILLER_ASAP7_75t_R FILLER_60_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1203 ();
 FILLER_ASAP7_75t_R FILLER_60_1209 ();
 FILLER_ASAP7_75t_R FILLER_60_1225 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_61_2 ();
 FILLER_ASAP7_75t_R FILLER_61_8 ();
 DECAPx6_ASAP7_75t_R FILLER_61_30 ();
 DECAPx2_ASAP7_75t_R FILLER_61_44 ();
 DECAPx1_ASAP7_75t_R FILLER_61_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_100 ();
 FILLER_ASAP7_75t_R FILLER_61_109 ();
 FILLER_ASAP7_75t_R FILLER_61_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_127 ();
 DECAPx4_ASAP7_75t_R FILLER_61_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_145 ();
 FILLER_ASAP7_75t_R FILLER_61_154 ();
 FILLER_ASAP7_75t_R FILLER_61_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_161 ();
 DECAPx10_ASAP7_75t_R FILLER_61_194 ();
 DECAPx2_ASAP7_75t_R FILLER_61_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_232 ();
 FILLER_ASAP7_75t_R FILLER_61_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_251 ();
 FILLER_ASAP7_75t_R FILLER_61_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_267 ();
 FILLER_ASAP7_75t_R FILLER_61_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_285 ();
 DECAPx10_ASAP7_75t_R FILLER_61_302 ();
 DECAPx6_ASAP7_75t_R FILLER_61_324 ();
 DECAPx1_ASAP7_75t_R FILLER_61_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_349 ();
 FILLER_ASAP7_75t_R FILLER_61_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_359 ();
 DECAPx2_ASAP7_75t_R FILLER_61_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_376 ();
 DECAPx10_ASAP7_75t_R FILLER_61_394 ();
 DECAPx6_ASAP7_75t_R FILLER_61_416 ();
 DECAPx2_ASAP7_75t_R FILLER_61_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_436 ();
 DECAPx6_ASAP7_75t_R FILLER_61_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_459 ();
 FILLER_ASAP7_75t_R FILLER_61_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_483 ();
 DECAPx1_ASAP7_75t_R FILLER_61_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_494 ();
 DECAPx10_ASAP7_75t_R FILLER_61_503 ();
 DECAPx10_ASAP7_75t_R FILLER_61_525 ();
 DECAPx4_ASAP7_75t_R FILLER_61_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_557 ();
 DECAPx6_ASAP7_75t_R FILLER_61_568 ();
 DECAPx1_ASAP7_75t_R FILLER_61_582 ();
 DECAPx4_ASAP7_75t_R FILLER_61_596 ();
 DECAPx2_ASAP7_75t_R FILLER_61_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_622 ();
 DECAPx10_ASAP7_75t_R FILLER_61_629 ();
 DECAPx10_ASAP7_75t_R FILLER_61_651 ();
 DECAPx10_ASAP7_75t_R FILLER_61_673 ();
 DECAPx10_ASAP7_75t_R FILLER_61_695 ();
 DECAPx10_ASAP7_75t_R FILLER_61_717 ();
 DECAPx2_ASAP7_75t_R FILLER_61_739 ();
 FILLER_ASAP7_75t_R FILLER_61_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_747 ();
 DECAPx10_ASAP7_75t_R FILLER_61_756 ();
 DECAPx10_ASAP7_75t_R FILLER_61_778 ();
 DECAPx10_ASAP7_75t_R FILLER_61_800 ();
 DECAPx2_ASAP7_75t_R FILLER_61_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_828 ();
 DECAPx2_ASAP7_75t_R FILLER_61_836 ();
 FILLER_ASAP7_75t_R FILLER_61_849 ();
 DECAPx4_ASAP7_75t_R FILLER_61_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_867 ();
 DECAPx10_ASAP7_75t_R FILLER_61_891 ();
 DECAPx1_ASAP7_75t_R FILLER_61_920 ();
 DECAPx2_ASAP7_75t_R FILLER_61_926 ();
 FILLER_ASAP7_75t_R FILLER_61_932 ();
 DECAPx10_ASAP7_75t_R FILLER_61_940 ();
 DECAPx6_ASAP7_75t_R FILLER_61_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_976 ();
 DECAPx10_ASAP7_75t_R FILLER_61_983 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1027 ();
 FILLER_ASAP7_75t_R FILLER_61_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1045 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1183 ();
 FILLER_ASAP7_75t_R FILLER_61_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1209 ();
 FILLER_ASAP7_75t_R FILLER_61_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_62_2 ();
 FILLER_ASAP7_75t_R FILLER_62_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_30 ();
 FILLER_ASAP7_75t_R FILLER_62_37 ();
 DECAPx10_ASAP7_75t_R FILLER_62_54 ();
 DECAPx6_ASAP7_75t_R FILLER_62_76 ();
 FILLER_ASAP7_75t_R FILLER_62_96 ();
 DECAPx2_ASAP7_75t_R FILLER_62_104 ();
 FILLER_ASAP7_75t_R FILLER_62_110 ();
 FILLER_ASAP7_75t_R FILLER_62_133 ();
 DECAPx10_ASAP7_75t_R FILLER_62_142 ();
 DECAPx2_ASAP7_75t_R FILLER_62_164 ();
 FILLER_ASAP7_75t_R FILLER_62_170 ();
 DECAPx10_ASAP7_75t_R FILLER_62_184 ();
 DECAPx2_ASAP7_75t_R FILLER_62_212 ();
 FILLER_ASAP7_75t_R FILLER_62_218 ();
 DECAPx6_ASAP7_75t_R FILLER_62_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_258 ();
 DECAPx10_ASAP7_75t_R FILLER_62_284 ();
 FILLER_ASAP7_75t_R FILLER_62_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_308 ();
 DECAPx10_ASAP7_75t_R FILLER_62_330 ();
 DECAPx10_ASAP7_75t_R FILLER_62_352 ();
 DECAPx10_ASAP7_75t_R FILLER_62_374 ();
 FILLER_ASAP7_75t_R FILLER_62_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_398 ();
 DECAPx4_ASAP7_75t_R FILLER_62_411 ();
 FILLER_ASAP7_75t_R FILLER_62_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_423 ();
 DECAPx2_ASAP7_75t_R FILLER_62_431 ();
 FILLER_ASAP7_75t_R FILLER_62_437 ();
 DECAPx6_ASAP7_75t_R FILLER_62_445 ();
 FILLER_ASAP7_75t_R FILLER_62_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_461 ();
 DECAPx10_ASAP7_75t_R FILLER_62_464 ();
 DECAPx10_ASAP7_75t_R FILLER_62_486 ();
 DECAPx2_ASAP7_75t_R FILLER_62_508 ();
 FILLER_ASAP7_75t_R FILLER_62_514 ();
 DECAPx6_ASAP7_75t_R FILLER_62_537 ();
 DECAPx2_ASAP7_75t_R FILLER_62_551 ();
 DECAPx10_ASAP7_75t_R FILLER_62_567 ();
 FILLER_ASAP7_75t_R FILLER_62_589 ();
 FILLER_ASAP7_75t_R FILLER_62_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_603 ();
 DECAPx10_ASAP7_75t_R FILLER_62_616 ();
 DECAPx2_ASAP7_75t_R FILLER_62_638 ();
 DECAPx10_ASAP7_75t_R FILLER_62_651 ();
 DECAPx10_ASAP7_75t_R FILLER_62_673 ();
 DECAPx2_ASAP7_75t_R FILLER_62_695 ();
 FILLER_ASAP7_75t_R FILLER_62_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_703 ();
 DECAPx2_ASAP7_75t_R FILLER_62_726 ();
 DECAPx10_ASAP7_75t_R FILLER_62_738 ();
 DECAPx10_ASAP7_75t_R FILLER_62_760 ();
 DECAPx10_ASAP7_75t_R FILLER_62_782 ();
 DECAPx10_ASAP7_75t_R FILLER_62_804 ();
 DECAPx10_ASAP7_75t_R FILLER_62_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_848 ();
 DECAPx1_ASAP7_75t_R FILLER_62_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_863 ();
 DECAPx10_ASAP7_75t_R FILLER_62_872 ();
 DECAPx6_ASAP7_75t_R FILLER_62_894 ();
 DECAPx2_ASAP7_75t_R FILLER_62_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_914 ();
 DECAPx10_ASAP7_75t_R FILLER_62_939 ();
 DECAPx4_ASAP7_75t_R FILLER_62_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_971 ();
 DECAPx10_ASAP7_75t_R FILLER_62_978 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_62_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1044 ();
 FILLER_ASAP7_75t_R FILLER_62_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1143 ();
 FILLER_ASAP7_75t_R FILLER_62_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1182 ();
 FILLER_ASAP7_75t_R FILLER_62_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1205 ();
 FILLER_ASAP7_75t_R FILLER_62_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1245 ();
 DECAPx6_ASAP7_75t_R FILLER_63_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_16 ();
 FILLER_ASAP7_75t_R FILLER_63_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_26 ();
 FILLER_ASAP7_75t_R FILLER_63_40 ();
 FILLER_ASAP7_75t_R FILLER_63_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_69 ();
 DECAPx6_ASAP7_75t_R FILLER_63_82 ();
 DECAPx1_ASAP7_75t_R FILLER_63_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_100 ();
 FILLER_ASAP7_75t_R FILLER_63_110 ();
 FILLER_ASAP7_75t_R FILLER_63_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_136 ();
 DECAPx2_ASAP7_75t_R FILLER_63_157 ();
 DECAPx6_ASAP7_75t_R FILLER_63_166 ();
 DECAPx2_ASAP7_75t_R FILLER_63_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_186 ();
 FILLER_ASAP7_75t_R FILLER_63_206 ();
 FILLER_ASAP7_75t_R FILLER_63_221 ();
 DECAPx1_ASAP7_75t_R FILLER_63_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_258 ();
 DECAPx10_ASAP7_75t_R FILLER_63_265 ();
 DECAPx10_ASAP7_75t_R FILLER_63_287 ();
 FILLER_ASAP7_75t_R FILLER_63_309 ();
 DECAPx6_ASAP7_75t_R FILLER_63_317 ();
 DECAPx2_ASAP7_75t_R FILLER_63_352 ();
 DECAPx10_ASAP7_75t_R FILLER_63_368 ();
 DECAPx4_ASAP7_75t_R FILLER_63_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_410 ();
 DECAPx2_ASAP7_75t_R FILLER_63_417 ();
 DECAPx6_ASAP7_75t_R FILLER_63_429 ();
 FILLER_ASAP7_75t_R FILLER_63_443 ();
 DECAPx10_ASAP7_75t_R FILLER_63_461 ();
 DECAPx10_ASAP7_75t_R FILLER_63_483 ();
 DECAPx4_ASAP7_75t_R FILLER_63_505 ();
 FILLER_ASAP7_75t_R FILLER_63_515 ();
 FILLER_ASAP7_75t_R FILLER_63_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_522 ();
 FILLER_ASAP7_75t_R FILLER_63_535 ();
 FILLER_ASAP7_75t_R FILLER_63_554 ();
 DECAPx10_ASAP7_75t_R FILLER_63_572 ();
 DECAPx10_ASAP7_75t_R FILLER_63_594 ();
 DECAPx10_ASAP7_75t_R FILLER_63_616 ();
 DECAPx2_ASAP7_75t_R FILLER_63_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_644 ();
 DECAPx10_ASAP7_75t_R FILLER_63_655 ();
 DECAPx2_ASAP7_75t_R FILLER_63_677 ();
 FILLER_ASAP7_75t_R FILLER_63_683 ();
 DECAPx10_ASAP7_75t_R FILLER_63_695 ();
 DECAPx6_ASAP7_75t_R FILLER_63_717 ();
 FILLER_ASAP7_75t_R FILLER_63_731 ();
 DECAPx4_ASAP7_75t_R FILLER_63_739 ();
 FILLER_ASAP7_75t_R FILLER_63_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_759 ();
 DECAPx6_ASAP7_75t_R FILLER_63_774 ();
 FILLER_ASAP7_75t_R FILLER_63_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_790 ();
 DECAPx10_ASAP7_75t_R FILLER_63_797 ();
 DECAPx10_ASAP7_75t_R FILLER_63_819 ();
 DECAPx10_ASAP7_75t_R FILLER_63_841 ();
 DECAPx10_ASAP7_75t_R FILLER_63_863 ();
 DECAPx10_ASAP7_75t_R FILLER_63_885 ();
 DECAPx6_ASAP7_75t_R FILLER_63_907 ();
 FILLER_ASAP7_75t_R FILLER_63_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_923 ();
 DECAPx6_ASAP7_75t_R FILLER_63_926 ();
 DECAPx10_ASAP7_75t_R FILLER_63_960 ();
 DECAPx10_ASAP7_75t_R FILLER_63_982 ();
 FILLER_ASAP7_75t_R FILLER_63_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1006 ();
 FILLER_ASAP7_75t_R FILLER_63_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1027 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1174 ();
 FILLER_ASAP7_75t_R FILLER_63_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1269 ();
 FILLER_ASAP7_75t_R FILLER_63_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_64_2 ();
 FILLER_ASAP7_75t_R FILLER_64_24 ();
 DECAPx4_ASAP7_75t_R FILLER_64_38 ();
 FILLER_ASAP7_75t_R FILLER_64_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_50 ();
 FILLER_ASAP7_75t_R FILLER_64_77 ();
 DECAPx1_ASAP7_75t_R FILLER_64_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_159 ();
 DECAPx4_ASAP7_75t_R FILLER_64_172 ();
 FILLER_ASAP7_75t_R FILLER_64_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_184 ();
 FILLER_ASAP7_75t_R FILLER_64_188 ();
 DECAPx2_ASAP7_75t_R FILLER_64_253 ();
 DECAPx10_ASAP7_75t_R FILLER_64_275 ();
 DECAPx6_ASAP7_75t_R FILLER_64_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_368 ();
 DECAPx4_ASAP7_75t_R FILLER_64_397 ();
 FILLER_ASAP7_75t_R FILLER_64_407 ();
 DECAPx2_ASAP7_75t_R FILLER_64_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_421 ();
 DECAPx10_ASAP7_75t_R FILLER_64_440 ();
 DECAPx2_ASAP7_75t_R FILLER_64_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_470 ();
 DECAPx4_ASAP7_75t_R FILLER_64_487 ();
 FILLER_ASAP7_75t_R FILLER_64_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_499 ();
 DECAPx6_ASAP7_75t_R FILLER_64_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_522 ();
 DECAPx2_ASAP7_75t_R FILLER_64_544 ();
 FILLER_ASAP7_75t_R FILLER_64_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_562 ();
 DECAPx10_ASAP7_75t_R FILLER_64_569 ();
 FILLER_ASAP7_75t_R FILLER_64_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_593 ();
 FILLER_ASAP7_75t_R FILLER_64_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_614 ();
 DECAPx2_ASAP7_75t_R FILLER_64_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_627 ();
 DECAPx2_ASAP7_75t_R FILLER_64_638 ();
 FILLER_ASAP7_75t_R FILLER_64_644 ();
 DECAPx6_ASAP7_75t_R FILLER_64_673 ();
 DECAPx1_ASAP7_75t_R FILLER_64_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_691 ();
 DECAPx10_ASAP7_75t_R FILLER_64_702 ();
 DECAPx10_ASAP7_75t_R FILLER_64_724 ();
 DECAPx6_ASAP7_75t_R FILLER_64_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_760 ();
 DECAPx4_ASAP7_75t_R FILLER_64_773 ();
 FILLER_ASAP7_75t_R FILLER_64_783 ();
 DECAPx2_ASAP7_75t_R FILLER_64_795 ();
 DECAPx10_ASAP7_75t_R FILLER_64_811 ();
 DECAPx4_ASAP7_75t_R FILLER_64_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_843 ();
 DECAPx10_ASAP7_75t_R FILLER_64_854 ();
 FILLER_ASAP7_75t_R FILLER_64_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_878 ();
 DECAPx2_ASAP7_75t_R FILLER_64_885 ();
 FILLER_ASAP7_75t_R FILLER_64_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_893 ();
 DECAPx10_ASAP7_75t_R FILLER_64_900 ();
 DECAPx4_ASAP7_75t_R FILLER_64_922 ();
 DECAPx4_ASAP7_75t_R FILLER_64_938 ();
 DECAPx4_ASAP7_75t_R FILLER_64_962 ();
 FILLER_ASAP7_75t_R FILLER_64_972 ();
 DECAPx1_ASAP7_75t_R FILLER_64_990 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1048 ();
 FILLER_ASAP7_75t_R FILLER_64_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1079 ();
 FILLER_ASAP7_75t_R FILLER_64_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1119 ();
 FILLER_ASAP7_75t_R FILLER_64_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1143 ();
 FILLER_ASAP7_75t_R FILLER_64_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1191 ();
 FILLER_ASAP7_75t_R FILLER_64_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1229 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1281 ();
 FILLER_ASAP7_75t_R FILLER_64_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_65_2 ();
 FILLER_ASAP7_75t_R FILLER_65_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_10 ();
 FILLER_ASAP7_75t_R FILLER_65_19 ();
 DECAPx1_ASAP7_75t_R FILLER_65_39 ();
 DECAPx6_ASAP7_75t_R FILLER_65_73 ();
 DECAPx1_ASAP7_75t_R FILLER_65_87 ();
 FILLER_ASAP7_75t_R FILLER_65_103 ();
 FILLER_ASAP7_75t_R FILLER_65_114 ();
 DECAPx1_ASAP7_75t_R FILLER_65_122 ();
 DECAPx2_ASAP7_75t_R FILLER_65_134 ();
 DECAPx2_ASAP7_75t_R FILLER_65_153 ();
 FILLER_ASAP7_75t_R FILLER_65_159 ();
 DECAPx2_ASAP7_75t_R FILLER_65_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_176 ();
 DECAPx2_ASAP7_75t_R FILLER_65_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_187 ();
 FILLER_ASAP7_75t_R FILLER_65_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_214 ();
 FILLER_ASAP7_75t_R FILLER_65_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_225 ();
 FILLER_ASAP7_75t_R FILLER_65_251 ();
 DECAPx1_ASAP7_75t_R FILLER_65_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_281 ();
 DECAPx1_ASAP7_75t_R FILLER_65_288 ();
 DECAPx6_ASAP7_75t_R FILLER_65_312 ();
 DECAPx1_ASAP7_75t_R FILLER_65_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_340 ();
 DECAPx1_ASAP7_75t_R FILLER_65_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_367 ();
 DECAPx6_ASAP7_75t_R FILLER_65_399 ();
 DECAPx2_ASAP7_75t_R FILLER_65_413 ();
 DECAPx4_ASAP7_75t_R FILLER_65_427 ();
 DECAPx1_ASAP7_75t_R FILLER_65_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_447 ();
 DECAPx4_ASAP7_75t_R FILLER_65_461 ();
 FILLER_ASAP7_75t_R FILLER_65_471 ();
 FILLER_ASAP7_75t_R FILLER_65_479 ();
 DECAPx1_ASAP7_75t_R FILLER_65_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_493 ();
 DECAPx10_ASAP7_75t_R FILLER_65_504 ();
 DECAPx6_ASAP7_75t_R FILLER_65_526 ();
 DECAPx2_ASAP7_75t_R FILLER_65_540 ();
 DECAPx4_ASAP7_75t_R FILLER_65_555 ();
 DECAPx4_ASAP7_75t_R FILLER_65_571 ();
 FILLER_ASAP7_75t_R FILLER_65_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_583 ();
 DECAPx10_ASAP7_75t_R FILLER_65_590 ();
 DECAPx1_ASAP7_75t_R FILLER_65_612 ();
 DECAPx1_ASAP7_75t_R FILLER_65_622 ();
 DECAPx6_ASAP7_75t_R FILLER_65_632 ();
 FILLER_ASAP7_75t_R FILLER_65_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_662 ();
 DECAPx10_ASAP7_75t_R FILLER_65_669 ();
 DECAPx4_ASAP7_75t_R FILLER_65_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_701 ();
 DECAPx10_ASAP7_75t_R FILLER_65_708 ();
 DECAPx10_ASAP7_75t_R FILLER_65_730 ();
 DECAPx10_ASAP7_75t_R FILLER_65_752 ();
 DECAPx6_ASAP7_75t_R FILLER_65_774 ();
 DECAPx10_ASAP7_75t_R FILLER_65_794 ();
 DECAPx10_ASAP7_75t_R FILLER_65_816 ();
 DECAPx10_ASAP7_75t_R FILLER_65_838 ();
 DECAPx2_ASAP7_75t_R FILLER_65_860 ();
 DECAPx10_ASAP7_75t_R FILLER_65_874 ();
 FILLER_ASAP7_75t_R FILLER_65_896 ();
 DECAPx6_ASAP7_75t_R FILLER_65_906 ();
 DECAPx1_ASAP7_75t_R FILLER_65_920 ();
 DECAPx2_ASAP7_75t_R FILLER_65_926 ();
 DECAPx10_ASAP7_75t_R FILLER_65_938 ();
 DECAPx6_ASAP7_75t_R FILLER_65_960 ();
 DECAPx1_ASAP7_75t_R FILLER_65_974 ();
 DECAPx10_ASAP7_75t_R FILLER_65_990 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1051 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1073 ();
 FILLER_ASAP7_75t_R FILLER_65_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1120 ();
 FILLER_ASAP7_75t_R FILLER_65_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1172 ();
 FILLER_ASAP7_75t_R FILLER_65_1207 ();
 FILLER_ASAP7_75t_R FILLER_65_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1245 ();
 FILLER_ASAP7_75t_R FILLER_65_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1255 ();
 FILLER_ASAP7_75t_R FILLER_65_1266 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_66_2 ();
 FILLER_ASAP7_75t_R FILLER_66_8 ();
 FILLER_ASAP7_75t_R FILLER_66_41 ();
 DECAPx10_ASAP7_75t_R FILLER_66_58 ();
 DECAPx6_ASAP7_75t_R FILLER_66_80 ();
 FILLER_ASAP7_75t_R FILLER_66_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_125 ();
 DECAPx4_ASAP7_75t_R FILLER_66_150 ();
 DECAPx2_ASAP7_75t_R FILLER_66_166 ();
 DECAPx2_ASAP7_75t_R FILLER_66_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_189 ();
 DECAPx10_ASAP7_75t_R FILLER_66_197 ();
 DECAPx1_ASAP7_75t_R FILLER_66_219 ();
 FILLER_ASAP7_75t_R FILLER_66_229 ();
 FILLER_ASAP7_75t_R FILLER_66_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_249 ();
 DECAPx4_ASAP7_75t_R FILLER_66_272 ();
 FILLER_ASAP7_75t_R FILLER_66_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_284 ();
 DECAPx4_ASAP7_75t_R FILLER_66_293 ();
 FILLER_ASAP7_75t_R FILLER_66_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_305 ();
 DECAPx1_ASAP7_75t_R FILLER_66_337 ();
 DECAPx1_ASAP7_75t_R FILLER_66_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_375 ();
 DECAPx10_ASAP7_75t_R FILLER_66_386 ();
 DECAPx4_ASAP7_75t_R FILLER_66_408 ();
 DECAPx4_ASAP7_75t_R FILLER_66_424 ();
 DECAPx2_ASAP7_75t_R FILLER_66_443 ();
 FILLER_ASAP7_75t_R FILLER_66_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_451 ();
 DECAPx2_ASAP7_75t_R FILLER_66_464 ();
 DECAPx2_ASAP7_75t_R FILLER_66_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_488 ();
 DECAPx10_ASAP7_75t_R FILLER_66_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_517 ();
 DECAPx1_ASAP7_75t_R FILLER_66_524 ();
 DECAPx10_ASAP7_75t_R FILLER_66_535 ();
 DECAPx6_ASAP7_75t_R FILLER_66_557 ();
 DECAPx1_ASAP7_75t_R FILLER_66_571 ();
 DECAPx10_ASAP7_75t_R FILLER_66_585 ();
 DECAPx4_ASAP7_75t_R FILLER_66_607 ();
 FILLER_ASAP7_75t_R FILLER_66_617 ();
 DECAPx10_ASAP7_75t_R FILLER_66_629 ();
 FILLER_ASAP7_75t_R FILLER_66_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_653 ();
 DECAPx4_ASAP7_75t_R FILLER_66_660 ();
 FILLER_ASAP7_75t_R FILLER_66_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_672 ();
 DECAPx10_ASAP7_75t_R FILLER_66_680 ();
 DECAPx10_ASAP7_75t_R FILLER_66_702 ();
 DECAPx6_ASAP7_75t_R FILLER_66_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_738 ();
 DECAPx6_ASAP7_75t_R FILLER_66_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_762 ();
 DECAPx10_ASAP7_75t_R FILLER_66_769 ();
 DECAPx6_ASAP7_75t_R FILLER_66_791 ();
 DECAPx1_ASAP7_75t_R FILLER_66_805 ();
 DECAPx6_ASAP7_75t_R FILLER_66_815 ();
 FILLER_ASAP7_75t_R FILLER_66_829 ();
 DECAPx6_ASAP7_75t_R FILLER_66_837 ();
 FILLER_ASAP7_75t_R FILLER_66_851 ();
 DECAPx10_ASAP7_75t_R FILLER_66_859 ();
 DECAPx10_ASAP7_75t_R FILLER_66_881 ();
 DECAPx10_ASAP7_75t_R FILLER_66_903 ();
 DECAPx4_ASAP7_75t_R FILLER_66_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_935 ();
 DECAPx10_ASAP7_75t_R FILLER_66_946 ();
 DECAPx10_ASAP7_75t_R FILLER_66_968 ();
 DECAPx10_ASAP7_75t_R FILLER_66_990 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1083 ();
 FILLER_ASAP7_75t_R FILLER_66_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1160 ();
 FILLER_ASAP7_75t_R FILLER_66_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1168 ();
 FILLER_ASAP7_75t_R FILLER_66_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1219 ();
 FILLER_ASAP7_75t_R FILLER_66_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_67_2 ();
 FILLER_ASAP7_75t_R FILLER_67_24 ();
 FILLER_ASAP7_75t_R FILLER_67_34 ();
 DECAPx2_ASAP7_75t_R FILLER_67_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_48 ();
 DECAPx10_ASAP7_75t_R FILLER_67_52 ();
 DECAPx2_ASAP7_75t_R FILLER_67_74 ();
 DECAPx1_ASAP7_75t_R FILLER_67_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_104 ();
 DECAPx2_ASAP7_75t_R FILLER_67_108 ();
 DECAPx10_ASAP7_75t_R FILLER_67_122 ();
 DECAPx10_ASAP7_75t_R FILLER_67_144 ();
 DECAPx6_ASAP7_75t_R FILLER_67_166 ();
 FILLER_ASAP7_75t_R FILLER_67_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_182 ();
 DECAPx1_ASAP7_75t_R FILLER_67_190 ();
 DECAPx1_ASAP7_75t_R FILLER_67_202 ();
 DECAPx1_ASAP7_75t_R FILLER_67_212 ();
 FILLER_ASAP7_75t_R FILLER_67_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_224 ();
 DECAPx4_ASAP7_75t_R FILLER_67_270 ();
 FILLER_ASAP7_75t_R FILLER_67_280 ();
 DECAPx1_ASAP7_75t_R FILLER_67_288 ();
 DECAPx10_ASAP7_75t_R FILLER_67_376 ();
 DECAPx2_ASAP7_75t_R FILLER_67_398 ();
 FILLER_ASAP7_75t_R FILLER_67_404 ();
 DECAPx1_ASAP7_75t_R FILLER_67_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_422 ();
 DECAPx10_ASAP7_75t_R FILLER_67_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_460 ();
 DECAPx1_ASAP7_75t_R FILLER_67_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_471 ();
 DECAPx10_ASAP7_75t_R FILLER_67_478 ();
 FILLER_ASAP7_75t_R FILLER_67_525 ();
 FILLER_ASAP7_75t_R FILLER_67_548 ();
 DECAPx4_ASAP7_75t_R FILLER_67_568 ();
 FILLER_ASAP7_75t_R FILLER_67_578 ();
 DECAPx10_ASAP7_75t_R FILLER_67_586 ();
 DECAPx10_ASAP7_75t_R FILLER_67_608 ();
 DECAPx10_ASAP7_75t_R FILLER_67_630 ();
 DECAPx10_ASAP7_75t_R FILLER_67_652 ();
 DECAPx6_ASAP7_75t_R FILLER_67_674 ();
 DECAPx1_ASAP7_75t_R FILLER_67_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_692 ();
 DECAPx4_ASAP7_75t_R FILLER_67_699 ();
 FILLER_ASAP7_75t_R FILLER_67_709 ();
 DECAPx10_ASAP7_75t_R FILLER_67_717 ();
 FILLER_ASAP7_75t_R FILLER_67_739 ();
 DECAPx10_ASAP7_75t_R FILLER_67_747 ();
 DECAPx10_ASAP7_75t_R FILLER_67_769 ();
 DECAPx10_ASAP7_75t_R FILLER_67_791 ();
 DECAPx10_ASAP7_75t_R FILLER_67_813 ();
 DECAPx10_ASAP7_75t_R FILLER_67_835 ();
 DECAPx10_ASAP7_75t_R FILLER_67_857 ();
 DECAPx10_ASAP7_75t_R FILLER_67_879 ();
 DECAPx2_ASAP7_75t_R FILLER_67_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_907 ();
 DECAPx2_ASAP7_75t_R FILLER_67_916 ();
 FILLER_ASAP7_75t_R FILLER_67_922 ();
 DECAPx10_ASAP7_75t_R FILLER_67_926 ();
 DECAPx10_ASAP7_75t_R FILLER_67_948 ();
 DECAPx10_ASAP7_75t_R FILLER_67_970 ();
 DECAPx10_ASAP7_75t_R FILLER_67_992 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1044 ();
 FILLER_ASAP7_75t_R FILLER_67_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1096 ();
 FILLER_ASAP7_75t_R FILLER_67_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1111 ();
 FILLER_ASAP7_75t_R FILLER_67_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1136 ();
 FILLER_ASAP7_75t_R FILLER_67_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1152 ();
 FILLER_ASAP7_75t_R FILLER_67_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1241 ();
 FILLER_ASAP7_75t_R FILLER_67_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_68_2 ();
 FILLER_ASAP7_75t_R FILLER_68_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_26 ();
 DECAPx1_ASAP7_75t_R FILLER_68_30 ();
 DECAPx2_ASAP7_75t_R FILLER_68_46 ();
 FILLER_ASAP7_75t_R FILLER_68_52 ();
 DECAPx2_ASAP7_75t_R FILLER_68_63 ();
 FILLER_ASAP7_75t_R FILLER_68_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_84 ();
 DECAPx6_ASAP7_75t_R FILLER_68_93 ();
 FILLER_ASAP7_75t_R FILLER_68_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_109 ();
 FILLER_ASAP7_75t_R FILLER_68_128 ();
 DECAPx6_ASAP7_75t_R FILLER_68_136 ();
 FILLER_ASAP7_75t_R FILLER_68_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_152 ();
 DECAPx10_ASAP7_75t_R FILLER_68_183 ();
 FILLER_ASAP7_75t_R FILLER_68_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_207 ();
 DECAPx2_ASAP7_75t_R FILLER_68_214 ();
 DECAPx1_ASAP7_75t_R FILLER_68_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_254 ();
 DECAPx4_ASAP7_75t_R FILLER_68_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_271 ();
 DECAPx2_ASAP7_75t_R FILLER_68_278 ();
 DECAPx1_ASAP7_75t_R FILLER_68_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_296 ();
 DECAPx4_ASAP7_75t_R FILLER_68_326 ();
 DECAPx10_ASAP7_75t_R FILLER_68_367 ();
 DECAPx10_ASAP7_75t_R FILLER_68_389 ();
 DECAPx10_ASAP7_75t_R FILLER_68_411 ();
 DECAPx10_ASAP7_75t_R FILLER_68_433 ();
 DECAPx2_ASAP7_75t_R FILLER_68_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_461 ();
 DECAPx4_ASAP7_75t_R FILLER_68_464 ();
 FILLER_ASAP7_75t_R FILLER_68_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_518 ();
 DECAPx2_ASAP7_75t_R FILLER_68_525 ();
 DECAPx2_ASAP7_75t_R FILLER_68_541 ();
 FILLER_ASAP7_75t_R FILLER_68_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_555 ();
 DECAPx2_ASAP7_75t_R FILLER_68_571 ();
 FILLER_ASAP7_75t_R FILLER_68_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_579 ();
 DECAPx2_ASAP7_75t_R FILLER_68_586 ();
 DECAPx10_ASAP7_75t_R FILLER_68_599 ();
 DECAPx1_ASAP7_75t_R FILLER_68_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_625 ();
 DECAPx2_ASAP7_75t_R FILLER_68_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_648 ();
 DECAPx10_ASAP7_75t_R FILLER_68_659 ();
 DECAPx10_ASAP7_75t_R FILLER_68_681 ();
 DECAPx6_ASAP7_75t_R FILLER_68_703 ();
 DECAPx10_ASAP7_75t_R FILLER_68_723 ();
 DECAPx10_ASAP7_75t_R FILLER_68_745 ();
 DECAPx6_ASAP7_75t_R FILLER_68_767 ();
 DECAPx2_ASAP7_75t_R FILLER_68_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_787 ();
 DECAPx10_ASAP7_75t_R FILLER_68_794 ();
 DECAPx10_ASAP7_75t_R FILLER_68_816 ();
 DECAPx6_ASAP7_75t_R FILLER_68_838 ();
 DECAPx2_ASAP7_75t_R FILLER_68_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_858 ();
 DECAPx10_ASAP7_75t_R FILLER_68_875 ();
 DECAPx10_ASAP7_75t_R FILLER_68_897 ();
 DECAPx10_ASAP7_75t_R FILLER_68_919 ();
 FILLER_ASAP7_75t_R FILLER_68_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_943 ();
 DECAPx4_ASAP7_75t_R FILLER_68_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_957 ();
 DECAPx4_ASAP7_75t_R FILLER_68_970 ();
 FILLER_ASAP7_75t_R FILLER_68_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_982 ();
 DECAPx10_ASAP7_75t_R FILLER_68_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1055 ();
 FILLER_ASAP7_75t_R FILLER_68_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1138 ();
 FILLER_ASAP7_75t_R FILLER_68_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1182 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1220 ();
 FILLER_ASAP7_75t_R FILLER_68_1226 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_69_2 ();
 FILLER_ASAP7_75t_R FILLER_69_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_37 ();
 DECAPx1_ASAP7_75t_R FILLER_69_41 ();
 FILLER_ASAP7_75t_R FILLER_69_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_77 ();
 DECAPx1_ASAP7_75t_R FILLER_69_84 ();
 DECAPx2_ASAP7_75t_R FILLER_69_95 ();
 FILLER_ASAP7_75t_R FILLER_69_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_111 ();
 FILLER_ASAP7_75t_R FILLER_69_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_144 ();
 DECAPx10_ASAP7_75t_R FILLER_69_165 ();
 FILLER_ASAP7_75t_R FILLER_69_187 ();
 DECAPx2_ASAP7_75t_R FILLER_69_195 ();
 DECAPx6_ASAP7_75t_R FILLER_69_248 ();
 FILLER_ASAP7_75t_R FILLER_69_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_272 ();
 DECAPx4_ASAP7_75t_R FILLER_69_287 ();
 DECAPx2_ASAP7_75t_R FILLER_69_327 ();
 DECAPx6_ASAP7_75t_R FILLER_69_350 ();
 FILLER_ASAP7_75t_R FILLER_69_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_374 ();
 DECAPx10_ASAP7_75t_R FILLER_69_385 ();
 DECAPx10_ASAP7_75t_R FILLER_69_417 ();
 DECAPx4_ASAP7_75t_R FILLER_69_439 ();
 DECAPx10_ASAP7_75t_R FILLER_69_455 ();
 DECAPx1_ASAP7_75t_R FILLER_69_477 ();
 DECAPx6_ASAP7_75t_R FILLER_69_495 ();
 DECAPx2_ASAP7_75t_R FILLER_69_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_522 ();
 DECAPx10_ASAP7_75t_R FILLER_69_531 ();
 DECAPx10_ASAP7_75t_R FILLER_69_553 ();
 DECAPx10_ASAP7_75t_R FILLER_69_575 ();
 DECAPx1_ASAP7_75t_R FILLER_69_597 ();
 DECAPx6_ASAP7_75t_R FILLER_69_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_647 ();
 DECAPx10_ASAP7_75t_R FILLER_69_655 ();
 DECAPx10_ASAP7_75t_R FILLER_69_677 ();
 DECAPx10_ASAP7_75t_R FILLER_69_699 ();
 DECAPx10_ASAP7_75t_R FILLER_69_721 ();
 DECAPx6_ASAP7_75t_R FILLER_69_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_757 ();
 DECAPx10_ASAP7_75t_R FILLER_69_764 ();
 DECAPx1_ASAP7_75t_R FILLER_69_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_790 ();
 DECAPx2_ASAP7_75t_R FILLER_69_797 ();
 FILLER_ASAP7_75t_R FILLER_69_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_805 ();
 DECAPx6_ASAP7_75t_R FILLER_69_812 ();
 DECAPx1_ASAP7_75t_R FILLER_69_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_830 ();
 DECAPx10_ASAP7_75t_R FILLER_69_838 ();
 DECAPx2_ASAP7_75t_R FILLER_69_860 ();
 FILLER_ASAP7_75t_R FILLER_69_866 ();
 DECAPx10_ASAP7_75t_R FILLER_69_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_896 ();
 DECAPx6_ASAP7_75t_R FILLER_69_904 ();
 DECAPx2_ASAP7_75t_R FILLER_69_918 ();
 FILLER_ASAP7_75t_R FILLER_69_926 ();
 DECAPx2_ASAP7_75t_R FILLER_69_934 ();
 FILLER_ASAP7_75t_R FILLER_69_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_942 ();
 FILLER_ASAP7_75t_R FILLER_69_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_963 ();
 DECAPx1_ASAP7_75t_R FILLER_69_978 ();
 DECAPx10_ASAP7_75t_R FILLER_69_990 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1012 ();
 FILLER_ASAP7_75t_R FILLER_69_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1078 ();
 FILLER_ASAP7_75t_R FILLER_69_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1130 ();
 FILLER_ASAP7_75t_R FILLER_69_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1215 ();
 FILLER_ASAP7_75t_R FILLER_69_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1224 ();
 FILLER_ASAP7_75t_R FILLER_69_1251 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1281 ();
 FILLER_ASAP7_75t_R FILLER_69_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_70_2 ();
 FILLER_ASAP7_75t_R FILLER_70_22 ();
 DECAPx1_ASAP7_75t_R FILLER_70_48 ();
 FILLER_ASAP7_75t_R FILLER_70_58 ();
 FILLER_ASAP7_75t_R FILLER_70_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_76 ();
 FILLER_ASAP7_75t_R FILLER_70_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_140 ();
 DECAPx2_ASAP7_75t_R FILLER_70_150 ();
 FILLER_ASAP7_75t_R FILLER_70_156 ();
 FILLER_ASAP7_75t_R FILLER_70_179 ();
 FILLER_ASAP7_75t_R FILLER_70_188 ();
 FILLER_ASAP7_75t_R FILLER_70_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_209 ();
 FILLER_ASAP7_75t_R FILLER_70_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_224 ();
 DECAPx10_ASAP7_75t_R FILLER_70_234 ();
 FILLER_ASAP7_75t_R FILLER_70_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_258 ();
 DECAPx10_ASAP7_75t_R FILLER_70_284 ();
 FILLER_ASAP7_75t_R FILLER_70_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_350 ();
 FILLER_ASAP7_75t_R FILLER_70_358 ();
 DECAPx4_ASAP7_75t_R FILLER_70_391 ();
 DECAPx10_ASAP7_75t_R FILLER_70_413 ();
 DECAPx2_ASAP7_75t_R FILLER_70_435 ();
 FILLER_ASAP7_75t_R FILLER_70_441 ();
 DECAPx2_ASAP7_75t_R FILLER_70_453 ();
 FILLER_ASAP7_75t_R FILLER_70_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_461 ();
 DECAPx10_ASAP7_75t_R FILLER_70_464 ();
 FILLER_ASAP7_75t_R FILLER_70_486 ();
 DECAPx2_ASAP7_75t_R FILLER_70_494 ();
 FILLER_ASAP7_75t_R FILLER_70_500 ();
 DECAPx6_ASAP7_75t_R FILLER_70_533 ();
 FILLER_ASAP7_75t_R FILLER_70_547 ();
 DECAPx10_ASAP7_75t_R FILLER_70_558 ();
 DECAPx10_ASAP7_75t_R FILLER_70_580 ();
 DECAPx10_ASAP7_75t_R FILLER_70_602 ();
 DECAPx10_ASAP7_75t_R FILLER_70_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_646 ();
 DECAPx10_ASAP7_75t_R FILLER_70_684 ();
 DECAPx2_ASAP7_75t_R FILLER_70_706 ();
 DECAPx4_ASAP7_75t_R FILLER_70_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_732 ();
 DECAPx10_ASAP7_75t_R FILLER_70_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_765 ();
 DECAPx2_ASAP7_75t_R FILLER_70_772 ();
 FILLER_ASAP7_75t_R FILLER_70_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_780 ();
 DECAPx6_ASAP7_75t_R FILLER_70_788 ();
 DECAPx2_ASAP7_75t_R FILLER_70_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_808 ();
 DECAPx10_ASAP7_75t_R FILLER_70_827 ();
 DECAPx10_ASAP7_75t_R FILLER_70_849 ();
 FILLER_ASAP7_75t_R FILLER_70_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_873 ();
 DECAPx6_ASAP7_75t_R FILLER_70_880 ();
 DECAPx1_ASAP7_75t_R FILLER_70_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_898 ();
 DECAPx6_ASAP7_75t_R FILLER_70_911 ();
 DECAPx2_ASAP7_75t_R FILLER_70_925 ();
 DECAPx2_ASAP7_75t_R FILLER_70_937 ();
 FILLER_ASAP7_75t_R FILLER_70_943 ();
 DECAPx4_ASAP7_75t_R FILLER_70_965 ();
 FILLER_ASAP7_75t_R FILLER_70_975 ();
 DECAPx10_ASAP7_75t_R FILLER_70_988 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1032 ();
 FILLER_ASAP7_75t_R FILLER_70_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1070 ();
 FILLER_ASAP7_75t_R FILLER_70_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_70_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1163 ();
 FILLER_ASAP7_75t_R FILLER_70_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1252 ();
 FILLER_ASAP7_75t_R FILLER_70_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1265 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1276 ();
 FILLER_ASAP7_75t_R FILLER_70_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_71_2 ();
 FILLER_ASAP7_75t_R FILLER_71_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_26 ();
 DECAPx2_ASAP7_75t_R FILLER_71_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_57 ();
 DECAPx4_ASAP7_75t_R FILLER_71_62 ();
 FILLER_ASAP7_75t_R FILLER_71_72 ();
 DECAPx2_ASAP7_75t_R FILLER_71_82 ();
 FILLER_ASAP7_75t_R FILLER_71_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_90 ();
 DECAPx6_ASAP7_75t_R FILLER_71_101 ();
 DECAPx1_ASAP7_75t_R FILLER_71_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_172 ();
 DECAPx2_ASAP7_75t_R FILLER_71_187 ();
 DECAPx6_ASAP7_75t_R FILLER_71_207 ();
 FILLER_ASAP7_75t_R FILLER_71_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_223 ();
 DECAPx1_ASAP7_75t_R FILLER_71_230 ();
 FILLER_ASAP7_75t_R FILLER_71_250 ();
 DECAPx1_ASAP7_75t_R FILLER_71_267 ();
 DECAPx6_ASAP7_75t_R FILLER_71_277 ();
 DECAPx2_ASAP7_75t_R FILLER_71_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_297 ();
 DECAPx4_ASAP7_75t_R FILLER_71_322 ();
 FILLER_ASAP7_75t_R FILLER_71_349 ();
 DECAPx10_ASAP7_75t_R FILLER_71_372 ();
 DECAPx6_ASAP7_75t_R FILLER_71_394 ();
 DECAPx2_ASAP7_75t_R FILLER_71_424 ();
 FILLER_ASAP7_75t_R FILLER_71_430 ();
 DECAPx6_ASAP7_75t_R FILLER_71_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_471 ();
 FILLER_ASAP7_75t_R FILLER_71_482 ();
 FILLER_ASAP7_75t_R FILLER_71_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_502 ();
 DECAPx2_ASAP7_75t_R FILLER_71_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_536 ();
 DECAPx1_ASAP7_75t_R FILLER_71_558 ();
 DECAPx4_ASAP7_75t_R FILLER_71_568 ();
 DECAPx10_ASAP7_75t_R FILLER_71_605 ();
 FILLER_ASAP7_75t_R FILLER_71_627 ();
 DECAPx6_ASAP7_75t_R FILLER_71_635 ();
 DECAPx2_ASAP7_75t_R FILLER_71_649 ();
 DECAPx10_ASAP7_75t_R FILLER_71_680 ();
 DECAPx10_ASAP7_75t_R FILLER_71_702 ();
 DECAPx10_ASAP7_75t_R FILLER_71_724 ();
 DECAPx10_ASAP7_75t_R FILLER_71_746 ();
 DECAPx2_ASAP7_75t_R FILLER_71_768 ();
 FILLER_ASAP7_75t_R FILLER_71_774 ();
 DECAPx10_ASAP7_75t_R FILLER_71_782 ();
 DECAPx10_ASAP7_75t_R FILLER_71_804 ();
 DECAPx10_ASAP7_75t_R FILLER_71_826 ();
 DECAPx10_ASAP7_75t_R FILLER_71_848 ();
 FILLER_ASAP7_75t_R FILLER_71_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_872 ();
 DECAPx10_ASAP7_75t_R FILLER_71_883 ();
 DECAPx6_ASAP7_75t_R FILLER_71_905 ();
 DECAPx1_ASAP7_75t_R FILLER_71_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_923 ();
 DECAPx6_ASAP7_75t_R FILLER_71_926 ();
 DECAPx1_ASAP7_75t_R FILLER_71_954 ();
 DECAPx10_ASAP7_75t_R FILLER_71_961 ();
 DECAPx6_ASAP7_75t_R FILLER_71_983 ();
 DECAPx2_ASAP7_75t_R FILLER_71_997 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1022 ();
 FILLER_ASAP7_75t_R FILLER_71_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1041 ();
 FILLER_ASAP7_75t_R FILLER_71_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1050 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1069 ();
 FILLER_ASAP7_75t_R FILLER_71_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1089 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1123 ();
 FILLER_ASAP7_75t_R FILLER_71_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1177 ();
 FILLER_ASAP7_75t_R FILLER_71_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1185 ();
 FILLER_ASAP7_75t_R FILLER_71_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1268 ();
 FILLER_ASAP7_75t_R FILLER_71_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_72_2 ();
 FILLER_ASAP7_75t_R FILLER_72_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_14 ();
 DECAPx6_ASAP7_75t_R FILLER_72_29 ();
 DECAPx10_ASAP7_75t_R FILLER_72_50 ();
 DECAPx6_ASAP7_75t_R FILLER_72_72 ();
 DECAPx2_ASAP7_75t_R FILLER_72_86 ();
 FILLER_ASAP7_75t_R FILLER_72_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_106 ();
 DECAPx4_ASAP7_75t_R FILLER_72_119 ();
 FILLER_ASAP7_75t_R FILLER_72_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_131 ();
 DECAPx1_ASAP7_75t_R FILLER_72_147 ();
 FILLER_ASAP7_75t_R FILLER_72_165 ();
 DECAPx10_ASAP7_75t_R FILLER_72_176 ();
 DECAPx10_ASAP7_75t_R FILLER_72_198 ();
 DECAPx1_ASAP7_75t_R FILLER_72_220 ();
 FILLER_ASAP7_75t_R FILLER_72_244 ();
 DECAPx2_ASAP7_75t_R FILLER_72_254 ();
 FILLER_ASAP7_75t_R FILLER_72_260 ();
 DECAPx6_ASAP7_75t_R FILLER_72_272 ();
 DECAPx2_ASAP7_75t_R FILLER_72_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_292 ();
 DECAPx6_ASAP7_75t_R FILLER_72_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_313 ();
 DECAPx10_ASAP7_75t_R FILLER_72_324 ();
 DECAPx2_ASAP7_75t_R FILLER_72_346 ();
 DECAPx10_ASAP7_75t_R FILLER_72_362 ();
 DECAPx6_ASAP7_75t_R FILLER_72_384 ();
 FILLER_ASAP7_75t_R FILLER_72_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_400 ();
 FILLER_ASAP7_75t_R FILLER_72_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_411 ();
 FILLER_ASAP7_75t_R FILLER_72_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_424 ();
 DECAPx4_ASAP7_75t_R FILLER_72_431 ();
 FILLER_ASAP7_75t_R FILLER_72_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_443 ();
 DECAPx4_ASAP7_75t_R FILLER_72_450 ();
 FILLER_ASAP7_75t_R FILLER_72_460 ();
 DECAPx10_ASAP7_75t_R FILLER_72_464 ();
 DECAPx6_ASAP7_75t_R FILLER_72_486 ();
 FILLER_ASAP7_75t_R FILLER_72_500 ();
 DECAPx1_ASAP7_75t_R FILLER_72_512 ();
 DECAPx6_ASAP7_75t_R FILLER_72_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_536 ();
 DECAPx4_ASAP7_75t_R FILLER_72_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_557 ();
 FILLER_ASAP7_75t_R FILLER_72_568 ();
 FILLER_ASAP7_75t_R FILLER_72_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_581 ();
 DECAPx10_ASAP7_75t_R FILLER_72_605 ();
 DECAPx1_ASAP7_75t_R FILLER_72_627 ();
 DECAPx10_ASAP7_75t_R FILLER_72_637 ();
 DECAPx6_ASAP7_75t_R FILLER_72_659 ();
 DECAPx1_ASAP7_75t_R FILLER_72_673 ();
 DECAPx10_ASAP7_75t_R FILLER_72_683 ();
 DECAPx1_ASAP7_75t_R FILLER_72_705 ();
 DECAPx10_ASAP7_75t_R FILLER_72_725 ();
 DECAPx4_ASAP7_75t_R FILLER_72_747 ();
 FILLER_ASAP7_75t_R FILLER_72_757 ();
 DECAPx10_ASAP7_75t_R FILLER_72_769 ();
 DECAPx10_ASAP7_75t_R FILLER_72_791 ();
 DECAPx2_ASAP7_75t_R FILLER_72_813 ();
 DECAPx6_ASAP7_75t_R FILLER_72_835 ();
 DECAPx1_ASAP7_75t_R FILLER_72_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_853 ();
 DECAPx10_ASAP7_75t_R FILLER_72_860 ();
 DECAPx10_ASAP7_75t_R FILLER_72_882 ();
 DECAPx10_ASAP7_75t_R FILLER_72_904 ();
 DECAPx2_ASAP7_75t_R FILLER_72_926 ();
 FILLER_ASAP7_75t_R FILLER_72_932 ();
 DECAPx6_ASAP7_75t_R FILLER_72_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_958 ();
 DECAPx10_ASAP7_75t_R FILLER_72_965 ();
 DECAPx10_ASAP7_75t_R FILLER_72_987 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1160 ();
 FILLER_ASAP7_75t_R FILLER_72_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1195 ();
 FILLER_ASAP7_75t_R FILLER_72_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1235 ();
 FILLER_ASAP7_75t_R FILLER_72_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_73_2 ();
 DECAPx6_ASAP7_75t_R FILLER_73_24 ();
 DECAPx6_ASAP7_75t_R FILLER_73_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_59 ();
 DECAPx2_ASAP7_75t_R FILLER_73_66 ();
 FILLER_ASAP7_75t_R FILLER_73_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_74 ();
 DECAPx2_ASAP7_75t_R FILLER_73_83 ();
 FILLER_ASAP7_75t_R FILLER_73_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_133 ();
 DECAPx10_ASAP7_75t_R FILLER_73_168 ();
 FILLER_ASAP7_75t_R FILLER_73_190 ();
 FILLER_ASAP7_75t_R FILLER_73_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_250 ();
 FILLER_ASAP7_75t_R FILLER_73_259 ();
 DECAPx2_ASAP7_75t_R FILLER_73_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_277 ();
 DECAPx4_ASAP7_75t_R FILLER_73_286 ();
 FILLER_ASAP7_75t_R FILLER_73_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_298 ();
 DECAPx6_ASAP7_75t_R FILLER_73_327 ();
 FILLER_ASAP7_75t_R FILLER_73_341 ();
 DECAPx1_ASAP7_75t_R FILLER_73_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_368 ();
 DECAPx1_ASAP7_75t_R FILLER_73_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_380 ();
 DECAPx6_ASAP7_75t_R FILLER_73_391 ();
 DECAPx4_ASAP7_75t_R FILLER_73_411 ();
 FILLER_ASAP7_75t_R FILLER_73_421 ();
 DECAPx6_ASAP7_75t_R FILLER_73_431 ();
 DECAPx1_ASAP7_75t_R FILLER_73_445 ();
 DECAPx10_ASAP7_75t_R FILLER_73_455 ();
 DECAPx4_ASAP7_75t_R FILLER_73_477 ();
 DECAPx6_ASAP7_75t_R FILLER_73_505 ();
 DECAPx2_ASAP7_75t_R FILLER_73_519 ();
 DECAPx2_ASAP7_75t_R FILLER_73_531 ();
 DECAPx10_ASAP7_75t_R FILLER_73_544 ();
 DECAPx10_ASAP7_75t_R FILLER_73_566 ();
 DECAPx4_ASAP7_75t_R FILLER_73_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_598 ();
 DECAPx10_ASAP7_75t_R FILLER_73_613 ();
 DECAPx4_ASAP7_75t_R FILLER_73_635 ();
 FILLER_ASAP7_75t_R FILLER_73_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_657 ();
 DECAPx1_ASAP7_75t_R FILLER_73_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_680 ();
 DECAPx10_ASAP7_75t_R FILLER_73_687 ();
 DECAPx10_ASAP7_75t_R FILLER_73_709 ();
 DECAPx6_ASAP7_75t_R FILLER_73_731 ();
 DECAPx10_ASAP7_75t_R FILLER_73_755 ();
 DECAPx2_ASAP7_75t_R FILLER_73_777 ();
 DECAPx10_ASAP7_75t_R FILLER_73_797 ();
 DECAPx10_ASAP7_75t_R FILLER_73_819 ();
 DECAPx4_ASAP7_75t_R FILLER_73_841 ();
 FILLER_ASAP7_75t_R FILLER_73_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_853 ();
 DECAPx6_ASAP7_75t_R FILLER_73_864 ();
 DECAPx2_ASAP7_75t_R FILLER_73_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_905 ();
 DECAPx4_ASAP7_75t_R FILLER_73_912 ();
 FILLER_ASAP7_75t_R FILLER_73_922 ();
 DECAPx4_ASAP7_75t_R FILLER_73_936 ();
 DECAPx1_ASAP7_75t_R FILLER_73_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_956 ();
 DECAPx6_ASAP7_75t_R FILLER_73_973 ();
 DECAPx2_ASAP7_75t_R FILLER_73_996 ();
 FILLER_ASAP7_75t_R FILLER_73_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1047 ();
 FILLER_ASAP7_75t_R FILLER_73_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1111 ();
 FILLER_ASAP7_75t_R FILLER_73_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1130 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1179 ();
 FILLER_ASAP7_75t_R FILLER_73_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1187 ();
 FILLER_ASAP7_75t_R FILLER_73_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1235 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_74_2 ();
 DECAPx10_ASAP7_75t_R FILLER_74_24 ();
 DECAPx6_ASAP7_75t_R FILLER_74_56 ();
 DECAPx1_ASAP7_75t_R FILLER_74_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_74 ();
 DECAPx2_ASAP7_75t_R FILLER_74_85 ();
 FILLER_ASAP7_75t_R FILLER_74_101 ();
 DECAPx6_ASAP7_75t_R FILLER_74_117 ();
 FILLER_ASAP7_75t_R FILLER_74_131 ();
 DECAPx10_ASAP7_75t_R FILLER_74_145 ();
 DECAPx4_ASAP7_75t_R FILLER_74_167 ();
 FILLER_ASAP7_75t_R FILLER_74_177 ();
 FILLER_ASAP7_75t_R FILLER_74_185 ();
 DECAPx2_ASAP7_75t_R FILLER_74_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_201 ();
 DECAPx2_ASAP7_75t_R FILLER_74_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_214 ();
 FILLER_ASAP7_75t_R FILLER_74_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_271 ();
 DECAPx10_ASAP7_75t_R FILLER_74_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_314 ();
 FILLER_ASAP7_75t_R FILLER_74_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_327 ();
 DECAPx6_ASAP7_75t_R FILLER_74_356 ();
 DECAPx4_ASAP7_75t_R FILLER_74_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_401 ();
 DECAPx2_ASAP7_75t_R FILLER_74_418 ();
 FILLER_ASAP7_75t_R FILLER_74_424 ();
 DECAPx6_ASAP7_75t_R FILLER_74_436 ();
 DECAPx1_ASAP7_75t_R FILLER_74_450 ();
 DECAPx10_ASAP7_75t_R FILLER_74_464 ();
 DECAPx6_ASAP7_75t_R FILLER_74_486 ();
 FILLER_ASAP7_75t_R FILLER_74_500 ();
 DECAPx10_ASAP7_75t_R FILLER_74_536 ();
 DECAPx10_ASAP7_75t_R FILLER_74_558 ();
 DECAPx2_ASAP7_75t_R FILLER_74_580 ();
 FILLER_ASAP7_75t_R FILLER_74_586 ();
 FILLER_ASAP7_75t_R FILLER_74_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_600 ();
 DECAPx1_ASAP7_75t_R FILLER_74_609 ();
 FILLER_ASAP7_75t_R FILLER_74_626 ();
 DECAPx10_ASAP7_75t_R FILLER_74_634 ();
 DECAPx6_ASAP7_75t_R FILLER_74_656 ();
 DECAPx2_ASAP7_75t_R FILLER_74_670 ();
 DECAPx10_ASAP7_75t_R FILLER_74_686 ();
 DECAPx10_ASAP7_75t_R FILLER_74_708 ();
 DECAPx10_ASAP7_75t_R FILLER_74_730 ();
 DECAPx10_ASAP7_75t_R FILLER_74_752 ();
 DECAPx6_ASAP7_75t_R FILLER_74_774 ();
 DECAPx1_ASAP7_75t_R FILLER_74_788 ();
 DECAPx10_ASAP7_75t_R FILLER_74_799 ();
 DECAPx10_ASAP7_75t_R FILLER_74_821 ();
 DECAPx10_ASAP7_75t_R FILLER_74_843 ();
 DECAPx10_ASAP7_75t_R FILLER_74_865 ();
 DECAPx10_ASAP7_75t_R FILLER_74_887 ();
 DECAPx10_ASAP7_75t_R FILLER_74_909 ();
 DECAPx2_ASAP7_75t_R FILLER_74_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_943 ();
 DECAPx10_ASAP7_75t_R FILLER_74_964 ();
 FILLER_ASAP7_75t_R FILLER_74_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_988 ();
 DECAPx10_ASAP7_75t_R FILLER_74_995 ();
 DECAPx10_ASAP7_75t_R FILLER_74_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1057 ();
 FILLER_ASAP7_75t_R FILLER_74_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1074 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1177 ();
 FILLER_ASAP7_75t_R FILLER_74_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1199 ();
 FILLER_ASAP7_75t_R FILLER_74_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_74_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1236 ();
 FILLER_ASAP7_75t_R FILLER_74_1252 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_75_2 ();
 DECAPx1_ASAP7_75t_R FILLER_75_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_20 ();
 DECAPx4_ASAP7_75t_R FILLER_75_48 ();
 DECAPx1_ASAP7_75t_R FILLER_75_64 ();
 DECAPx2_ASAP7_75t_R FILLER_75_98 ();
 FILLER_ASAP7_75t_R FILLER_75_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_106 ();
 DECAPx10_ASAP7_75t_R FILLER_75_115 ();
 DECAPx10_ASAP7_75t_R FILLER_75_137 ();
 FILLER_ASAP7_75t_R FILLER_75_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_161 ();
 FILLER_ASAP7_75t_R FILLER_75_185 ();
 DECAPx2_ASAP7_75t_R FILLER_75_194 ();
 FILLER_ASAP7_75t_R FILLER_75_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_211 ();
 DECAPx1_ASAP7_75t_R FILLER_75_219 ();
 DECAPx6_ASAP7_75t_R FILLER_75_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_243 ();
 DECAPx10_ASAP7_75t_R FILLER_75_250 ();
 DECAPx10_ASAP7_75t_R FILLER_75_272 ();
 DECAPx1_ASAP7_75t_R FILLER_75_294 ();
 DECAPx2_ASAP7_75t_R FILLER_75_319 ();
 DECAPx6_ASAP7_75t_R FILLER_75_352 ();
 FILLER_ASAP7_75t_R FILLER_75_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_368 ();
 DECAPx2_ASAP7_75t_R FILLER_75_376 ();
 FILLER_ASAP7_75t_R FILLER_75_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_384 ();
 DECAPx1_ASAP7_75t_R FILLER_75_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_410 ();
 DECAPx2_ASAP7_75t_R FILLER_75_449 ();
 FILLER_ASAP7_75t_R FILLER_75_455 ();
 DECAPx6_ASAP7_75t_R FILLER_75_471 ();
 DECAPx2_ASAP7_75t_R FILLER_75_485 ();
 DECAPx1_ASAP7_75t_R FILLER_75_512 ();
 FILLER_ASAP7_75t_R FILLER_75_536 ();
 DECAPx10_ASAP7_75t_R FILLER_75_559 ();
 FILLER_ASAP7_75t_R FILLER_75_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_583 ();
 DECAPx10_ASAP7_75t_R FILLER_75_611 ();
 DECAPx10_ASAP7_75t_R FILLER_75_633 ();
 DECAPx10_ASAP7_75t_R FILLER_75_655 ();
 DECAPx1_ASAP7_75t_R FILLER_75_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_681 ();
 DECAPx10_ASAP7_75t_R FILLER_75_688 ();
 DECAPx2_ASAP7_75t_R FILLER_75_710 ();
 FILLER_ASAP7_75t_R FILLER_75_716 ();
 DECAPx10_ASAP7_75t_R FILLER_75_724 ();
 DECAPx10_ASAP7_75t_R FILLER_75_746 ();
 DECAPx10_ASAP7_75t_R FILLER_75_768 ();
 DECAPx10_ASAP7_75t_R FILLER_75_790 ();
 DECAPx10_ASAP7_75t_R FILLER_75_812 ();
 DECAPx10_ASAP7_75t_R FILLER_75_834 ();
 DECAPx10_ASAP7_75t_R FILLER_75_856 ();
 DECAPx10_ASAP7_75t_R FILLER_75_878 ();
 DECAPx10_ASAP7_75t_R FILLER_75_900 ();
 FILLER_ASAP7_75t_R FILLER_75_922 ();
 DECAPx1_ASAP7_75t_R FILLER_75_926 ();
 DECAPx10_ASAP7_75t_R FILLER_75_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_968 ();
 DECAPx10_ASAP7_75t_R FILLER_75_998 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1070 ();
 FILLER_ASAP7_75t_R FILLER_75_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1116 ();
 FILLER_ASAP7_75t_R FILLER_75_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1214 ();
 FILLER_ASAP7_75t_R FILLER_75_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_76_2 ();
 DECAPx2_ASAP7_75t_R FILLER_76_24 ();
 FILLER_ASAP7_75t_R FILLER_76_30 ();
 DECAPx1_ASAP7_75t_R FILLER_76_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_44 ();
 DECAPx6_ASAP7_75t_R FILLER_76_51 ();
 DECAPx2_ASAP7_75t_R FILLER_76_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_77 ();
 DECAPx2_ASAP7_75t_R FILLER_76_101 ();
 DECAPx2_ASAP7_75t_R FILLER_76_115 ();
 DECAPx1_ASAP7_75t_R FILLER_76_129 ();
 DECAPx1_ASAP7_75t_R FILLER_76_140 ();
 DECAPx10_ASAP7_75t_R FILLER_76_162 ();
 FILLER_ASAP7_75t_R FILLER_76_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_201 ();
 DECAPx6_ASAP7_75t_R FILLER_76_218 ();
 DECAPx2_ASAP7_75t_R FILLER_76_232 ();
 DECAPx2_ASAP7_75t_R FILLER_76_265 ();
 DECAPx1_ASAP7_75t_R FILLER_76_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_291 ();
 DECAPx2_ASAP7_75t_R FILLER_76_302 ();
 FILLER_ASAP7_75t_R FILLER_76_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_310 ();
 DECAPx1_ASAP7_75t_R FILLER_76_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_343 ();
 DECAPx1_ASAP7_75t_R FILLER_76_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_390 ();
 FILLER_ASAP7_75t_R FILLER_76_398 ();
 DECAPx6_ASAP7_75t_R FILLER_76_410 ();
 DECAPx2_ASAP7_75t_R FILLER_76_424 ();
 DECAPx6_ASAP7_75t_R FILLER_76_436 ();
 FILLER_ASAP7_75t_R FILLER_76_450 ();
 DECAPx10_ASAP7_75t_R FILLER_76_474 ();
 DECAPx10_ASAP7_75t_R FILLER_76_502 ();
 DECAPx1_ASAP7_75t_R FILLER_76_524 ();
 FILLER_ASAP7_75t_R FILLER_76_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_537 ();
 DECAPx10_ASAP7_75t_R FILLER_76_554 ();
 DECAPx4_ASAP7_75t_R FILLER_76_576 ();
 DECAPx10_ASAP7_75t_R FILLER_76_607 ();
 DECAPx2_ASAP7_75t_R FILLER_76_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_635 ();
 DECAPx10_ASAP7_75t_R FILLER_76_646 ();
 DECAPx10_ASAP7_75t_R FILLER_76_668 ();
 DECAPx10_ASAP7_75t_R FILLER_76_690 ();
 DECAPx10_ASAP7_75t_R FILLER_76_712 ();
 DECAPx2_ASAP7_75t_R FILLER_76_734 ();
 DECAPx10_ASAP7_75t_R FILLER_76_750 ();
 DECAPx4_ASAP7_75t_R FILLER_76_772 ();
 DECAPx10_ASAP7_75t_R FILLER_76_788 ();
 DECAPx4_ASAP7_75t_R FILLER_76_810 ();
 FILLER_ASAP7_75t_R FILLER_76_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_822 ();
 DECAPx10_ASAP7_75t_R FILLER_76_830 ();
 DECAPx10_ASAP7_75t_R FILLER_76_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_874 ();
 DECAPx10_ASAP7_75t_R FILLER_76_883 ();
 DECAPx10_ASAP7_75t_R FILLER_76_905 ();
 DECAPx10_ASAP7_75t_R FILLER_76_927 ();
 DECAPx6_ASAP7_75t_R FILLER_76_949 ();
 DECAPx2_ASAP7_75t_R FILLER_76_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_969 ();
 DECAPx10_ASAP7_75t_R FILLER_76_978 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1074 ();
 FILLER_ASAP7_75t_R FILLER_76_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1100 ();
 FILLER_ASAP7_75t_R FILLER_76_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1207 ();
 FILLER_ASAP7_75t_R FILLER_76_1221 ();
 FILLER_ASAP7_75t_R FILLER_76_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1240 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_77_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_24 ();
 DECAPx2_ASAP7_75t_R FILLER_77_33 ();
 FILLER_ASAP7_75t_R FILLER_77_57 ();
 FILLER_ASAP7_75t_R FILLER_77_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_70 ();
 DECAPx4_ASAP7_75t_R FILLER_77_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_87 ();
 FILLER_ASAP7_75t_R FILLER_77_96 ();
 FILLER_ASAP7_75t_R FILLER_77_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_115 ();
 FILLER_ASAP7_75t_R FILLER_77_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_133 ();
 DECAPx2_ASAP7_75t_R FILLER_77_153 ();
 DECAPx6_ASAP7_75t_R FILLER_77_175 ();
 DECAPx2_ASAP7_75t_R FILLER_77_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_195 ();
 FILLER_ASAP7_75t_R FILLER_77_212 ();
 FILLER_ASAP7_75t_R FILLER_77_270 ();
 FILLER_ASAP7_75t_R FILLER_77_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_280 ();
 DECAPx1_ASAP7_75t_R FILLER_77_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_293 ();
 DECAPx1_ASAP7_75t_R FILLER_77_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_305 ();
 DECAPx1_ASAP7_75t_R FILLER_77_314 ();
 DECAPx2_ASAP7_75t_R FILLER_77_328 ();
 FILLER_ASAP7_75t_R FILLER_77_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_357 ();
 DECAPx2_ASAP7_75t_R FILLER_77_368 ();
 DECAPx10_ASAP7_75t_R FILLER_77_384 ();
 DECAPx4_ASAP7_75t_R FILLER_77_406 ();
 FILLER_ASAP7_75t_R FILLER_77_428 ();
 DECAPx10_ASAP7_75t_R FILLER_77_442 ();
 DECAPx4_ASAP7_75t_R FILLER_77_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_474 ();
 DECAPx2_ASAP7_75t_R FILLER_77_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_489 ();
 DECAPx2_ASAP7_75t_R FILLER_77_503 ();
 DECAPx10_ASAP7_75t_R FILLER_77_515 ();
 DECAPx1_ASAP7_75t_R FILLER_77_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_548 ();
 FILLER_ASAP7_75t_R FILLER_77_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_557 ();
 DECAPx2_ASAP7_75t_R FILLER_77_568 ();
 FILLER_ASAP7_75t_R FILLER_77_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_576 ();
 FILLER_ASAP7_75t_R FILLER_77_598 ();
 DECAPx2_ASAP7_75t_R FILLER_77_616 ();
 FILLER_ASAP7_75t_R FILLER_77_622 ();
 DECAPx10_ASAP7_75t_R FILLER_77_652 ();
 DECAPx6_ASAP7_75t_R FILLER_77_674 ();
 DECAPx1_ASAP7_75t_R FILLER_77_688 ();
 DECAPx10_ASAP7_75t_R FILLER_77_700 ();
 DECAPx10_ASAP7_75t_R FILLER_77_722 ();
 FILLER_ASAP7_75t_R FILLER_77_744 ();
 DECAPx10_ASAP7_75t_R FILLER_77_752 ();
 DECAPx4_ASAP7_75t_R FILLER_77_774 ();
 FILLER_ASAP7_75t_R FILLER_77_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_786 ();
 DECAPx10_ASAP7_75t_R FILLER_77_793 ();
 DECAPx10_ASAP7_75t_R FILLER_77_815 ();
 DECAPx2_ASAP7_75t_R FILLER_77_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_843 ();
 DECAPx4_ASAP7_75t_R FILLER_77_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_860 ();
 DECAPx6_ASAP7_75t_R FILLER_77_877 ();
 DECAPx1_ASAP7_75t_R FILLER_77_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_895 ();
 DECAPx4_ASAP7_75t_R FILLER_77_912 ();
 FILLER_ASAP7_75t_R FILLER_77_922 ();
 FILLER_ASAP7_75t_R FILLER_77_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_928 ();
 DECAPx10_ASAP7_75t_R FILLER_77_936 ();
 DECAPx10_ASAP7_75t_R FILLER_77_958 ();
 DECAPx10_ASAP7_75t_R FILLER_77_980 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1156 ();
 FILLER_ASAP7_75t_R FILLER_77_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_77_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1202 ();
 FILLER_ASAP7_75t_R FILLER_77_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1229 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1250 ();
 FILLER_ASAP7_75t_R FILLER_77_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_78_2 ();
 DECAPx2_ASAP7_75t_R FILLER_78_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_29 ();
 DECAPx1_ASAP7_75t_R FILLER_78_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_56 ();
 DECAPx2_ASAP7_75t_R FILLER_78_67 ();
 FILLER_ASAP7_75t_R FILLER_78_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_97 ();
 DECAPx1_ASAP7_75t_R FILLER_78_112 ();
 DECAPx1_ASAP7_75t_R FILLER_78_124 ();
 DECAPx10_ASAP7_75t_R FILLER_78_157 ();
 FILLER_ASAP7_75t_R FILLER_78_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_181 ();
 DECAPx2_ASAP7_75t_R FILLER_78_188 ();
 DECAPx4_ASAP7_75t_R FILLER_78_210 ();
 FILLER_ASAP7_75t_R FILLER_78_220 ();
 DECAPx4_ASAP7_75t_R FILLER_78_228 ();
 DECAPx6_ASAP7_75t_R FILLER_78_244 ();
 DECAPx6_ASAP7_75t_R FILLER_78_270 ();
 DECAPx1_ASAP7_75t_R FILLER_78_295 ();
 DECAPx2_ASAP7_75t_R FILLER_78_305 ();
 FILLER_ASAP7_75t_R FILLER_78_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_313 ();
 DECAPx2_ASAP7_75t_R FILLER_78_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_335 ();
 FILLER_ASAP7_75t_R FILLER_78_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_390 ();
 DECAPx6_ASAP7_75t_R FILLER_78_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_411 ();
 DECAPx6_ASAP7_75t_R FILLER_78_420 ();
 DECAPx2_ASAP7_75t_R FILLER_78_434 ();
 DECAPx6_ASAP7_75t_R FILLER_78_446 ();
 FILLER_ASAP7_75t_R FILLER_78_460 ();
 DECAPx1_ASAP7_75t_R FILLER_78_476 ();
 DECAPx4_ASAP7_75t_R FILLER_78_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_500 ();
 DECAPx10_ASAP7_75t_R FILLER_78_508 ();
 DECAPx10_ASAP7_75t_R FILLER_78_530 ();
 DECAPx1_ASAP7_75t_R FILLER_78_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_556 ();
 DECAPx6_ASAP7_75t_R FILLER_78_585 ();
 DECAPx2_ASAP7_75t_R FILLER_78_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_611 ();
 FILLER_ASAP7_75t_R FILLER_78_618 ();
 DECAPx2_ASAP7_75t_R FILLER_78_626 ();
 DECAPx2_ASAP7_75t_R FILLER_78_642 ();
 DECAPx6_ASAP7_75t_R FILLER_78_672 ();
 DECAPx2_ASAP7_75t_R FILLER_78_686 ();
 DECAPx10_ASAP7_75t_R FILLER_78_699 ();
 DECAPx10_ASAP7_75t_R FILLER_78_721 ();
 DECAPx1_ASAP7_75t_R FILLER_78_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_747 ();
 DECAPx2_ASAP7_75t_R FILLER_78_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_762 ();
 DECAPx10_ASAP7_75t_R FILLER_78_769 ();
 DECAPx10_ASAP7_75t_R FILLER_78_791 ();
 DECAPx6_ASAP7_75t_R FILLER_78_813 ();
 FILLER_ASAP7_75t_R FILLER_78_827 ();
 DECAPx4_ASAP7_75t_R FILLER_78_853 ();
 DECAPx10_ASAP7_75t_R FILLER_78_869 ();
 DECAPx10_ASAP7_75t_R FILLER_78_891 ();
 DECAPx10_ASAP7_75t_R FILLER_78_913 ();
 DECAPx6_ASAP7_75t_R FILLER_78_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_949 ();
 DECAPx10_ASAP7_75t_R FILLER_78_960 ();
 DECAPx10_ASAP7_75t_R FILLER_78_982 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1125 ();
 FILLER_ASAP7_75t_R FILLER_78_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1170 ();
 FILLER_ASAP7_75t_R FILLER_78_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1255 ();
 DECAPx4_ASAP7_75t_R FILLER_78_1281 ();
 FILLER_ASAP7_75t_R FILLER_78_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_79_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_16 ();
 DECAPx6_ASAP7_75t_R FILLER_79_27 ();
 FILLER_ASAP7_75t_R FILLER_79_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_43 ();
 FILLER_ASAP7_75t_R FILLER_79_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_113 ();
 DECAPx4_ASAP7_75t_R FILLER_79_134 ();
 DECAPx2_ASAP7_75t_R FILLER_79_152 ();
 FILLER_ASAP7_75t_R FILLER_79_158 ();
 DECAPx10_ASAP7_75t_R FILLER_79_167 ();
 FILLER_ASAP7_75t_R FILLER_79_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_191 ();
 FILLER_ASAP7_75t_R FILLER_79_208 ();
 DECAPx2_ASAP7_75t_R FILLER_79_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_237 ();
 DECAPx1_ASAP7_75t_R FILLER_79_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_263 ();
 DECAPx2_ASAP7_75t_R FILLER_79_274 ();
 DECAPx10_ASAP7_75t_R FILLER_79_288 ();
 DECAPx1_ASAP7_75t_R FILLER_79_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_335 ();
 DECAPx1_ASAP7_75t_R FILLER_79_366 ();
 DECAPx2_ASAP7_75t_R FILLER_79_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_383 ();
 FILLER_ASAP7_75t_R FILLER_79_391 ();
 DECAPx10_ASAP7_75t_R FILLER_79_409 ();
 DECAPx1_ASAP7_75t_R FILLER_79_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_435 ();
 DECAPx1_ASAP7_75t_R FILLER_79_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_446 ();
 DECAPx6_ASAP7_75t_R FILLER_79_459 ();
 DECAPx2_ASAP7_75t_R FILLER_79_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_479 ();
 DECAPx6_ASAP7_75t_R FILLER_79_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_504 ();
 DECAPx1_ASAP7_75t_R FILLER_79_532 ();
 DECAPx10_ASAP7_75t_R FILLER_79_546 ();
 DECAPx2_ASAP7_75t_R FILLER_79_568 ();
 FILLER_ASAP7_75t_R FILLER_79_574 ();
 DECAPx2_ASAP7_75t_R FILLER_79_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_589 ();
 DECAPx6_ASAP7_75t_R FILLER_79_600 ();
 FILLER_ASAP7_75t_R FILLER_79_614 ();
 DECAPx10_ASAP7_75t_R FILLER_79_626 ();
 DECAPx6_ASAP7_75t_R FILLER_79_648 ();
 FILLER_ASAP7_75t_R FILLER_79_662 ();
 DECAPx10_ASAP7_75t_R FILLER_79_674 ();
 DECAPx4_ASAP7_75t_R FILLER_79_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_706 ();
 DECAPx10_ASAP7_75t_R FILLER_79_724 ();
 DECAPx10_ASAP7_75t_R FILLER_79_746 ();
 DECAPx10_ASAP7_75t_R FILLER_79_768 ();
 DECAPx10_ASAP7_75t_R FILLER_79_790 ();
 DECAPx2_ASAP7_75t_R FILLER_79_812 ();
 FILLER_ASAP7_75t_R FILLER_79_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_820 ();
 DECAPx10_ASAP7_75t_R FILLER_79_827 ();
 DECAPx10_ASAP7_75t_R FILLER_79_849 ();
 DECAPx1_ASAP7_75t_R FILLER_79_871 ();
 DECAPx10_ASAP7_75t_R FILLER_79_887 ();
 DECAPx6_ASAP7_75t_R FILLER_79_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_923 ();
 DECAPx10_ASAP7_75t_R FILLER_79_951 ();
 DECAPx4_ASAP7_75t_R FILLER_79_973 ();
 DECAPx10_ASAP7_75t_R FILLER_79_990 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1012 ();
 FILLER_ASAP7_75t_R FILLER_79_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1090 ();
 FILLER_ASAP7_75t_R FILLER_79_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1182 ();
 FILLER_ASAP7_75t_R FILLER_79_1189 ();
 FILLER_ASAP7_75t_R FILLER_79_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1268 ();
 FILLER_ASAP7_75t_R FILLER_79_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_80_2 ();
 FILLER_ASAP7_75t_R FILLER_80_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_18 ();
 DECAPx1_ASAP7_75t_R FILLER_80_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_31 ();
 DECAPx4_ASAP7_75t_R FILLER_80_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_68 ();
 DECAPx2_ASAP7_75t_R FILLER_80_83 ();
 FILLER_ASAP7_75t_R FILLER_80_89 ();
 DECAPx4_ASAP7_75t_R FILLER_80_104 ();
 FILLER_ASAP7_75t_R FILLER_80_114 ();
 FILLER_ASAP7_75t_R FILLER_80_122 ();
 DECAPx4_ASAP7_75t_R FILLER_80_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_180 ();
 DECAPx1_ASAP7_75t_R FILLER_80_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_210 ();
 DECAPx10_ASAP7_75t_R FILLER_80_236 ();
 DECAPx2_ASAP7_75t_R FILLER_80_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_264 ();
 FILLER_ASAP7_75t_R FILLER_80_275 ();
 DECAPx1_ASAP7_75t_R FILLER_80_285 ();
 FILLER_ASAP7_75t_R FILLER_80_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_313 ();
 DECAPx1_ASAP7_75t_R FILLER_80_348 ();
 FILLER_ASAP7_75t_R FILLER_80_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_364 ();
 DECAPx4_ASAP7_75t_R FILLER_80_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_452 ();
 DECAPx4_ASAP7_75t_R FILLER_80_464 ();
 FILLER_ASAP7_75t_R FILLER_80_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_476 ();
 FILLER_ASAP7_75t_R FILLER_80_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_491 ();
 DECAPx2_ASAP7_75t_R FILLER_80_500 ();
 DECAPx2_ASAP7_75t_R FILLER_80_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_533 ();
 DECAPx6_ASAP7_75t_R FILLER_80_565 ();
 DECAPx2_ASAP7_75t_R FILLER_80_579 ();
 DECAPx6_ASAP7_75t_R FILLER_80_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_627 ();
 DECAPx6_ASAP7_75t_R FILLER_80_656 ();
 DECAPx6_ASAP7_75t_R FILLER_80_676 ();
 DECAPx1_ASAP7_75t_R FILLER_80_690 ();
 DECAPx10_ASAP7_75t_R FILLER_80_708 ();
 DECAPx10_ASAP7_75t_R FILLER_80_730 ();
 DECAPx10_ASAP7_75t_R FILLER_80_752 ();
 DECAPx10_ASAP7_75t_R FILLER_80_774 ();
 FILLER_ASAP7_75t_R FILLER_80_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_798 ();
 FILLER_ASAP7_75t_R FILLER_80_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_807 ();
 DECAPx2_ASAP7_75t_R FILLER_80_814 ();
 FILLER_ASAP7_75t_R FILLER_80_820 ();
 DECAPx10_ASAP7_75t_R FILLER_80_836 ();
 DECAPx10_ASAP7_75t_R FILLER_80_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_880 ();
 DECAPx10_ASAP7_75t_R FILLER_80_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_911 ();
 DECAPx10_ASAP7_75t_R FILLER_80_926 ();
 DECAPx6_ASAP7_75t_R FILLER_80_948 ();
 FILLER_ASAP7_75t_R FILLER_80_962 ();
 DECAPx4_ASAP7_75t_R FILLER_80_974 ();
 DECAPx10_ASAP7_75t_R FILLER_80_994 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1048 ();
 FILLER_ASAP7_75t_R FILLER_80_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1131 ();
 FILLER_ASAP7_75t_R FILLER_80_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1213 ();
 DECAPx4_ASAP7_75t_R FILLER_80_1244 ();
 FILLER_ASAP7_75t_R FILLER_80_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1256 ();
 FILLER_ASAP7_75t_R FILLER_80_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1266 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1284 ();
 FILLER_ASAP7_75t_R FILLER_80_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_81_2 ();
 DECAPx2_ASAP7_75t_R FILLER_81_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_22 ();
 DECAPx10_ASAP7_75t_R FILLER_81_29 ();
 FILLER_ASAP7_75t_R FILLER_81_51 ();
 DECAPx1_ASAP7_75t_R FILLER_81_61 ();
 DECAPx2_ASAP7_75t_R FILLER_81_73 ();
 FILLER_ASAP7_75t_R FILLER_81_79 ();
 FILLER_ASAP7_75t_R FILLER_81_94 ();
 DECAPx1_ASAP7_75t_R FILLER_81_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_112 ();
 DECAPx6_ASAP7_75t_R FILLER_81_120 ();
 DECAPx1_ASAP7_75t_R FILLER_81_134 ();
 DECAPx1_ASAP7_75t_R FILLER_81_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_189 ();
 DECAPx2_ASAP7_75t_R FILLER_81_198 ();
 FILLER_ASAP7_75t_R FILLER_81_204 ();
 FILLER_ASAP7_75t_R FILLER_81_213 ();
 DECAPx4_ASAP7_75t_R FILLER_81_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_238 ();
 DECAPx10_ASAP7_75t_R FILLER_81_255 ();
 DECAPx6_ASAP7_75t_R FILLER_81_277 ();
 DECAPx2_ASAP7_75t_R FILLER_81_307 ();
 DECAPx4_ASAP7_75t_R FILLER_81_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_360 ();
 DECAPx1_ASAP7_75t_R FILLER_81_382 ();
 DECAPx1_ASAP7_75t_R FILLER_81_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_419 ();
 DECAPx6_ASAP7_75t_R FILLER_81_432 ();
 FILLER_ASAP7_75t_R FILLER_81_446 ();
 DECAPx6_ASAP7_75t_R FILLER_81_454 ();
 FILLER_ASAP7_75t_R FILLER_81_468 ();
 DECAPx1_ASAP7_75t_R FILLER_81_476 ();
 FILLER_ASAP7_75t_R FILLER_81_492 ();
 DECAPx2_ASAP7_75t_R FILLER_81_504 ();
 FILLER_ASAP7_75t_R FILLER_81_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_523 ();
 DECAPx1_ASAP7_75t_R FILLER_81_530 ();
 DECAPx1_ASAP7_75t_R FILLER_81_562 ();
 DECAPx10_ASAP7_75t_R FILLER_81_582 ();
 DECAPx10_ASAP7_75t_R FILLER_81_604 ();
 DECAPx2_ASAP7_75t_R FILLER_81_626 ();
 DECAPx1_ASAP7_75t_R FILLER_81_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_643 ();
 DECAPx10_ASAP7_75t_R FILLER_81_668 ();
 DECAPx10_ASAP7_75t_R FILLER_81_690 ();
 DECAPx10_ASAP7_75t_R FILLER_81_712 ();
 DECAPx10_ASAP7_75t_R FILLER_81_734 ();
 DECAPx10_ASAP7_75t_R FILLER_81_756 ();
 DECAPx10_ASAP7_75t_R FILLER_81_778 ();
 DECAPx10_ASAP7_75t_R FILLER_81_800 ();
 DECAPx10_ASAP7_75t_R FILLER_81_822 ();
 DECAPx10_ASAP7_75t_R FILLER_81_844 ();
 DECAPx10_ASAP7_75t_R FILLER_81_866 ();
 DECAPx10_ASAP7_75t_R FILLER_81_888 ();
 DECAPx6_ASAP7_75t_R FILLER_81_910 ();
 DECAPx10_ASAP7_75t_R FILLER_81_926 ();
 DECAPx6_ASAP7_75t_R FILLER_81_948 ();
 DECAPx1_ASAP7_75t_R FILLER_81_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_966 ();
 DECAPx4_ASAP7_75t_R FILLER_81_973 ();
 FILLER_ASAP7_75t_R FILLER_81_983 ();
 DECAPx6_ASAP7_75t_R FILLER_81_991 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1161 ();
 FILLER_ASAP7_75t_R FILLER_81_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1211 ();
 FILLER_ASAP7_75t_R FILLER_81_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1245 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_82_2 ();
 FILLER_ASAP7_75t_R FILLER_82_16 ();
 DECAPx4_ASAP7_75t_R FILLER_82_31 ();
 DECAPx2_ASAP7_75t_R FILLER_82_48 ();
 DECAPx4_ASAP7_75t_R FILLER_82_66 ();
 FILLER_ASAP7_75t_R FILLER_82_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_78 ();
 DECAPx1_ASAP7_75t_R FILLER_82_91 ();
 DECAPx4_ASAP7_75t_R FILLER_82_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_125 ();
 DECAPx2_ASAP7_75t_R FILLER_82_139 ();
 FILLER_ASAP7_75t_R FILLER_82_145 ();
 DECAPx2_ASAP7_75t_R FILLER_82_155 ();
 FILLER_ASAP7_75t_R FILLER_82_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_169 ();
 FILLER_ASAP7_75t_R FILLER_82_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_188 ();
 DECAPx4_ASAP7_75t_R FILLER_82_204 ();
 FILLER_ASAP7_75t_R FILLER_82_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_216 ();
 DECAPx4_ASAP7_75t_R FILLER_82_224 ();
 FILLER_ASAP7_75t_R FILLER_82_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_236 ();
 DECAPx6_ASAP7_75t_R FILLER_82_248 ();
 FILLER_ASAP7_75t_R FILLER_82_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_264 ();
 DECAPx1_ASAP7_75t_R FILLER_82_272 ();
 DECAPx2_ASAP7_75t_R FILLER_82_282 ();
 FILLER_ASAP7_75t_R FILLER_82_288 ();
 DECAPx6_ASAP7_75t_R FILLER_82_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_332 ();
 FILLER_ASAP7_75t_R FILLER_82_343 ();
 DECAPx10_ASAP7_75t_R FILLER_82_384 ();
 DECAPx6_ASAP7_75t_R FILLER_82_406 ();
 DECAPx2_ASAP7_75t_R FILLER_82_420 ();
 DECAPx10_ASAP7_75t_R FILLER_82_438 ();
 FILLER_ASAP7_75t_R FILLER_82_460 ();
 DECAPx1_ASAP7_75t_R FILLER_82_464 ();
 DECAPx10_ASAP7_75t_R FILLER_82_476 ();
 DECAPx4_ASAP7_75t_R FILLER_82_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_508 ();
 DECAPx2_ASAP7_75t_R FILLER_82_517 ();
 DECAPx4_ASAP7_75t_R FILLER_82_529 ();
 FILLER_ASAP7_75t_R FILLER_82_539 ();
 DECAPx1_ASAP7_75t_R FILLER_82_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_562 ();
 DECAPx2_ASAP7_75t_R FILLER_82_569 ();
 DECAPx6_ASAP7_75t_R FILLER_82_585 ();
 DECAPx1_ASAP7_75t_R FILLER_82_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_603 ();
 FILLER_ASAP7_75t_R FILLER_82_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_624 ();
 FILLER_ASAP7_75t_R FILLER_82_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_658 ();
 DECAPx10_ASAP7_75t_R FILLER_82_673 ();
 DECAPx1_ASAP7_75t_R FILLER_82_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_699 ();
 DECAPx2_ASAP7_75t_R FILLER_82_724 ();
 FILLER_ASAP7_75t_R FILLER_82_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_732 ();
 DECAPx10_ASAP7_75t_R FILLER_82_743 ();
 DECAPx4_ASAP7_75t_R FILLER_82_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_775 ();
 DECAPx10_ASAP7_75t_R FILLER_82_786 ();
 DECAPx10_ASAP7_75t_R FILLER_82_808 ();
 DECAPx6_ASAP7_75t_R FILLER_82_830 ();
 FILLER_ASAP7_75t_R FILLER_82_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_846 ();
 DECAPx10_ASAP7_75t_R FILLER_82_857 ();
 DECAPx10_ASAP7_75t_R FILLER_82_879 ();
 DECAPx6_ASAP7_75t_R FILLER_82_901 ();
 DECAPx1_ASAP7_75t_R FILLER_82_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_919 ();
 DECAPx10_ASAP7_75t_R FILLER_82_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_952 ();
 DECAPx10_ASAP7_75t_R FILLER_82_962 ();
 DECAPx10_ASAP7_75t_R FILLER_82_984 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_82_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_82_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1152 ();
 FILLER_ASAP7_75t_R FILLER_82_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1218 ();
 FILLER_ASAP7_75t_R FILLER_82_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1242 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1266 ();
 DECAPx6_ASAP7_75t_R FILLER_83_2 ();
 FILLER_ASAP7_75t_R FILLER_83_16 ();
 DECAPx2_ASAP7_75t_R FILLER_83_24 ();
 FILLER_ASAP7_75t_R FILLER_83_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_32 ();
 DECAPx1_ASAP7_75t_R FILLER_83_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_51 ();
 DECAPx2_ASAP7_75t_R FILLER_83_74 ();
 FILLER_ASAP7_75t_R FILLER_83_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_82 ();
 DECAPx1_ASAP7_75t_R FILLER_83_89 ();
 FILLER_ASAP7_75t_R FILLER_83_120 ();
 FILLER_ASAP7_75t_R FILLER_83_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_132 ();
 DECAPx2_ASAP7_75t_R FILLER_83_141 ();
 DECAPx6_ASAP7_75t_R FILLER_83_161 ();
 DECAPx2_ASAP7_75t_R FILLER_83_190 ();
 DECAPx10_ASAP7_75t_R FILLER_83_209 ();
 FILLER_ASAP7_75t_R FILLER_83_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_233 ();
 DECAPx2_ASAP7_75t_R FILLER_83_246 ();
 FILLER_ASAP7_75t_R FILLER_83_268 ();
 DECAPx10_ASAP7_75t_R FILLER_83_296 ();
 DECAPx4_ASAP7_75t_R FILLER_83_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_328 ();
 FILLER_ASAP7_75t_R FILLER_83_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_338 ();
 DECAPx6_ASAP7_75t_R FILLER_83_347 ();
 DECAPx10_ASAP7_75t_R FILLER_83_377 ();
 DECAPx4_ASAP7_75t_R FILLER_83_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_409 ();
 DECAPx1_ASAP7_75t_R FILLER_83_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_447 ();
 FILLER_ASAP7_75t_R FILLER_83_469 ();
 DECAPx6_ASAP7_75t_R FILLER_83_492 ();
 FILLER_ASAP7_75t_R FILLER_83_506 ();
 DECAPx2_ASAP7_75t_R FILLER_83_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_524 ();
 DECAPx4_ASAP7_75t_R FILLER_83_535 ();
 DECAPx1_ASAP7_75t_R FILLER_83_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_592 ();
 DECAPx6_ASAP7_75t_R FILLER_83_601 ();
 FILLER_ASAP7_75t_R FILLER_83_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_617 ();
 DECAPx10_ASAP7_75t_R FILLER_83_626 ();
 DECAPx6_ASAP7_75t_R FILLER_83_648 ();
 DECAPx1_ASAP7_75t_R FILLER_83_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_666 ();
 DECAPx10_ASAP7_75t_R FILLER_83_687 ();
 DECAPx10_ASAP7_75t_R FILLER_83_709 ();
 DECAPx10_ASAP7_75t_R FILLER_83_731 ();
 DECAPx4_ASAP7_75t_R FILLER_83_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_763 ();
 DECAPx10_ASAP7_75t_R FILLER_83_770 ();
 DECAPx10_ASAP7_75t_R FILLER_83_792 ();
 DECAPx10_ASAP7_75t_R FILLER_83_814 ();
 DECAPx10_ASAP7_75t_R FILLER_83_836 ();
 DECAPx10_ASAP7_75t_R FILLER_83_858 ();
 DECAPx4_ASAP7_75t_R FILLER_83_880 ();
 FILLER_ASAP7_75t_R FILLER_83_890 ();
 DECAPx2_ASAP7_75t_R FILLER_83_900 ();
 FILLER_ASAP7_75t_R FILLER_83_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_908 ();
 DECAPx2_ASAP7_75t_R FILLER_83_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_923 ();
 DECAPx6_ASAP7_75t_R FILLER_83_926 ();
 FILLER_ASAP7_75t_R FILLER_83_940 ();
 DECAPx4_ASAP7_75t_R FILLER_83_952 ();
 FILLER_ASAP7_75t_R FILLER_83_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_964 ();
 DECAPx10_ASAP7_75t_R FILLER_83_971 ();
 DECAPx10_ASAP7_75t_R FILLER_83_993 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1234 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_84_2 ();
 DECAPx1_ASAP7_75t_R FILLER_84_16 ();
 DECAPx4_ASAP7_75t_R FILLER_84_26 ();
 FILLER_ASAP7_75t_R FILLER_84_36 ();
 DECAPx1_ASAP7_75t_R FILLER_84_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_48 ();
 FILLER_ASAP7_75t_R FILLER_84_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_57 ();
 FILLER_ASAP7_75t_R FILLER_84_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_69 ();
 DECAPx10_ASAP7_75t_R FILLER_84_80 ();
 DECAPx2_ASAP7_75t_R FILLER_84_102 ();
 FILLER_ASAP7_75t_R FILLER_84_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_110 ();
 DECAPx4_ASAP7_75t_R FILLER_84_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_127 ();
 FILLER_ASAP7_75t_R FILLER_84_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_145 ();
 DECAPx2_ASAP7_75t_R FILLER_84_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_168 ();
 DECAPx10_ASAP7_75t_R FILLER_84_177 ();
 DECAPx4_ASAP7_75t_R FILLER_84_205 ();
 FILLER_ASAP7_75t_R FILLER_84_215 ();
 DECAPx4_ASAP7_75t_R FILLER_84_227 ();
 FILLER_ASAP7_75t_R FILLER_84_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_239 ();
 DECAPx2_ASAP7_75t_R FILLER_84_256 ();
 FILLER_ASAP7_75t_R FILLER_84_262 ();
 DECAPx10_ASAP7_75t_R FILLER_84_274 ();
 DECAPx10_ASAP7_75t_R FILLER_84_296 ();
 DECAPx4_ASAP7_75t_R FILLER_84_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_328 ();
 DECAPx4_ASAP7_75t_R FILLER_84_350 ();
 FILLER_ASAP7_75t_R FILLER_84_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_362 ();
 FILLER_ASAP7_75t_R FILLER_84_370 ();
 DECAPx2_ASAP7_75t_R FILLER_84_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_422 ();
 DECAPx1_ASAP7_75t_R FILLER_84_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_461 ();
 DECAPx1_ASAP7_75t_R FILLER_84_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_468 ();
 DECAPx2_ASAP7_75t_R FILLER_84_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_501 ();
 FILLER_ASAP7_75t_R FILLER_84_508 ();
 FILLER_ASAP7_75t_R FILLER_84_517 ();
 DECAPx4_ASAP7_75t_R FILLER_84_529 ();
 FILLER_ASAP7_75t_R FILLER_84_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_541 ();
 FILLER_ASAP7_75t_R FILLER_84_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_579 ();
 FILLER_ASAP7_75t_R FILLER_84_602 ();
 DECAPx2_ASAP7_75t_R FILLER_84_614 ();
 DECAPx10_ASAP7_75t_R FILLER_84_672 ();
 DECAPx10_ASAP7_75t_R FILLER_84_694 ();
 DECAPx10_ASAP7_75t_R FILLER_84_716 ();
 DECAPx10_ASAP7_75t_R FILLER_84_738 ();
 DECAPx10_ASAP7_75t_R FILLER_84_760 ();
 DECAPx10_ASAP7_75t_R FILLER_84_782 ();
 DECAPx10_ASAP7_75t_R FILLER_84_804 ();
 DECAPx10_ASAP7_75t_R FILLER_84_826 ();
 DECAPx10_ASAP7_75t_R FILLER_84_848 ();
 DECAPx10_ASAP7_75t_R FILLER_84_870 ();
 DECAPx10_ASAP7_75t_R FILLER_84_892 ();
 FILLER_ASAP7_75t_R FILLER_84_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_916 ();
 DECAPx6_ASAP7_75t_R FILLER_84_929 ();
 DECAPx2_ASAP7_75t_R FILLER_84_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_949 ();
 DECAPx6_ASAP7_75t_R FILLER_84_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_976 ();
 DECAPx2_ASAP7_75t_R FILLER_84_986 ();
 FILLER_ASAP7_75t_R FILLER_84_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_994 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1031 ();
 FILLER_ASAP7_75t_R FILLER_84_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1064 ();
 FILLER_ASAP7_75t_R FILLER_84_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1117 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1179 ();
 FILLER_ASAP7_75t_R FILLER_84_1187 ();
 FILLER_ASAP7_75t_R FILLER_84_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1250 ();
 FILLER_ASAP7_75t_R FILLER_84_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_85_2 ();
 DECAPx1_ASAP7_75t_R FILLER_85_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_20 ();
 DECAPx10_ASAP7_75t_R FILLER_85_39 ();
 DECAPx2_ASAP7_75t_R FILLER_85_61 ();
 FILLER_ASAP7_75t_R FILLER_85_67 ();
 DECAPx2_ASAP7_75t_R FILLER_85_75 ();
 DECAPx10_ASAP7_75t_R FILLER_85_94 ();
 DECAPx10_ASAP7_75t_R FILLER_85_116 ();
 FILLER_ASAP7_75t_R FILLER_85_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_140 ();
 FILLER_ASAP7_75t_R FILLER_85_163 ();
 DECAPx4_ASAP7_75t_R FILLER_85_193 ();
 FILLER_ASAP7_75t_R FILLER_85_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_221 ();
 FILLER_ASAP7_75t_R FILLER_85_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_248 ();
 FILLER_ASAP7_75t_R FILLER_85_259 ();
 DECAPx6_ASAP7_75t_R FILLER_85_267 ();
 DECAPx1_ASAP7_75t_R FILLER_85_281 ();
 DECAPx4_ASAP7_75t_R FILLER_85_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_305 ();
 DECAPx6_ASAP7_75t_R FILLER_85_316 ();
 DECAPx1_ASAP7_75t_R FILLER_85_330 ();
 DECAPx6_ASAP7_75t_R FILLER_85_344 ();
 FILLER_ASAP7_75t_R FILLER_85_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_360 ();
 FILLER_ASAP7_75t_R FILLER_85_382 ();
 DECAPx6_ASAP7_75t_R FILLER_85_405 ();
 DECAPx10_ASAP7_75t_R FILLER_85_457 ();
 DECAPx4_ASAP7_75t_R FILLER_85_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_489 ();
 FILLER_ASAP7_75t_R FILLER_85_499 ();
 FILLER_ASAP7_75t_R FILLER_85_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_572 ();
 DECAPx1_ASAP7_75t_R FILLER_85_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_590 ();
 DECAPx6_ASAP7_75t_R FILLER_85_597 ();
 DECAPx2_ASAP7_75t_R FILLER_85_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_635 ();
 DECAPx1_ASAP7_75t_R FILLER_85_653 ();
 DECAPx10_ASAP7_75t_R FILLER_85_669 ();
 FILLER_ASAP7_75t_R FILLER_85_691 ();
 DECAPx2_ASAP7_75t_R FILLER_85_703 ();
 FILLER_ASAP7_75t_R FILLER_85_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_711 ();
 DECAPx6_ASAP7_75t_R FILLER_85_722 ();
 DECAPx2_ASAP7_75t_R FILLER_85_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_742 ();
 DECAPx6_ASAP7_75t_R FILLER_85_763 ();
 FILLER_ASAP7_75t_R FILLER_85_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_779 ();
 DECAPx2_ASAP7_75t_R FILLER_85_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_792 ();
 DECAPx10_ASAP7_75t_R FILLER_85_800 ();
 DECAPx2_ASAP7_75t_R FILLER_85_822 ();
 FILLER_ASAP7_75t_R FILLER_85_828 ();
 DECAPx2_ASAP7_75t_R FILLER_85_836 ();
 FILLER_ASAP7_75t_R FILLER_85_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_844 ();
 DECAPx4_ASAP7_75t_R FILLER_85_855 ();
 DECAPx6_ASAP7_75t_R FILLER_85_873 ();
 DECAPx1_ASAP7_75t_R FILLER_85_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_891 ();
 DECAPx10_ASAP7_75t_R FILLER_85_902 ();
 DECAPx10_ASAP7_75t_R FILLER_85_926 ();
 DECAPx10_ASAP7_75t_R FILLER_85_948 ();
 DECAPx10_ASAP7_75t_R FILLER_85_970 ();
 FILLER_ASAP7_75t_R FILLER_85_992 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1032 ();
 FILLER_ASAP7_75t_R FILLER_85_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1080 ();
 FILLER_ASAP7_75t_R FILLER_85_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1184 ();
 FILLER_ASAP7_75t_R FILLER_85_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1220 ();
 FILLER_ASAP7_75t_R FILLER_85_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_86_2 ();
 DECAPx4_ASAP7_75t_R FILLER_86_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_34 ();
 DECAPx6_ASAP7_75t_R FILLER_86_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_61 ();
 DECAPx1_ASAP7_75t_R FILLER_86_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_96 ();
 FILLER_ASAP7_75t_R FILLER_86_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_105 ();
 FILLER_ASAP7_75t_R FILLER_86_137 ();
 DECAPx2_ASAP7_75t_R FILLER_86_153 ();
 FILLER_ASAP7_75t_R FILLER_86_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_161 ();
 FILLER_ASAP7_75t_R FILLER_86_174 ();
 FILLER_ASAP7_75t_R FILLER_86_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_228 ();
 DECAPx1_ASAP7_75t_R FILLER_86_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_241 ();
 FILLER_ASAP7_75t_R FILLER_86_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_258 ();
 DECAPx2_ASAP7_75t_R FILLER_86_269 ();
 FILLER_ASAP7_75t_R FILLER_86_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_277 ();
 DECAPx6_ASAP7_75t_R FILLER_86_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_300 ();
 DECAPx4_ASAP7_75t_R FILLER_86_311 ();
 FILLER_ASAP7_75t_R FILLER_86_321 ();
 FILLER_ASAP7_75t_R FILLER_86_351 ();
 DECAPx4_ASAP7_75t_R FILLER_86_363 ();
 FILLER_ASAP7_75t_R FILLER_86_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_383 ();
 DECAPx2_ASAP7_75t_R FILLER_86_401 ();
 FILLER_ASAP7_75t_R FILLER_86_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_440 ();
 DECAPx4_ASAP7_75t_R FILLER_86_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_461 ();
 DECAPx10_ASAP7_75t_R FILLER_86_464 ();
 FILLER_ASAP7_75t_R FILLER_86_486 ();
 DECAPx10_ASAP7_75t_R FILLER_86_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_531 ();
 DECAPx4_ASAP7_75t_R FILLER_86_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_557 ();
 DECAPx2_ASAP7_75t_R FILLER_86_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_574 ();
 DECAPx2_ASAP7_75t_R FILLER_86_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_598 ();
 DECAPx10_ASAP7_75t_R FILLER_86_627 ();
 FILLER_ASAP7_75t_R FILLER_86_649 ();
 DECAPx6_ASAP7_75t_R FILLER_86_657 ();
 FILLER_ASAP7_75t_R FILLER_86_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_673 ();
 DECAPx10_ASAP7_75t_R FILLER_86_682 ();
 DECAPx2_ASAP7_75t_R FILLER_86_704 ();
 FILLER_ASAP7_75t_R FILLER_86_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_730 ();
 DECAPx6_ASAP7_75t_R FILLER_86_741 ();
 DECAPx1_ASAP7_75t_R FILLER_86_755 ();
 DECAPx6_ASAP7_75t_R FILLER_86_767 ();
 DECAPx1_ASAP7_75t_R FILLER_86_781 ();
 DECAPx10_ASAP7_75t_R FILLER_86_792 ();
 DECAPx6_ASAP7_75t_R FILLER_86_814 ();
 FILLER_ASAP7_75t_R FILLER_86_828 ();
 DECAPx10_ASAP7_75t_R FILLER_86_838 ();
 DECAPx10_ASAP7_75t_R FILLER_86_860 ();
 DECAPx10_ASAP7_75t_R FILLER_86_882 ();
 DECAPx10_ASAP7_75t_R FILLER_86_904 ();
 DECAPx6_ASAP7_75t_R FILLER_86_926 ();
 FILLER_ASAP7_75t_R FILLER_86_940 ();
 DECAPx10_ASAP7_75t_R FILLER_86_951 ();
 DECAPx10_ASAP7_75t_R FILLER_86_973 ();
 DECAPx1_ASAP7_75t_R FILLER_86_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_999 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1118 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1152 ();
 FILLER_ASAP7_75t_R FILLER_86_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1204 ();
 FILLER_ASAP7_75t_R FILLER_86_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1236 ();
 FILLER_ASAP7_75t_R FILLER_86_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1248 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1256 ();
 FILLER_ASAP7_75t_R FILLER_86_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_87_2 ();
 FILLER_ASAP7_75t_R FILLER_87_24 ();
 DECAPx2_ASAP7_75t_R FILLER_87_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_40 ();
 DECAPx10_ASAP7_75t_R FILLER_87_55 ();
 DECAPx2_ASAP7_75t_R FILLER_87_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_83 ();
 DECAPx1_ASAP7_75t_R FILLER_87_105 ();
 DECAPx6_ASAP7_75t_R FILLER_87_115 ();
 DECAPx6_ASAP7_75t_R FILLER_87_151 ();
 DECAPx1_ASAP7_75t_R FILLER_87_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_169 ();
 DECAPx4_ASAP7_75t_R FILLER_87_193 ();
 FILLER_ASAP7_75t_R FILLER_87_211 ();
 DECAPx10_ASAP7_75t_R FILLER_87_220 ();
 DECAPx10_ASAP7_75t_R FILLER_87_251 ();
 DECAPx10_ASAP7_75t_R FILLER_87_273 ();
 DECAPx10_ASAP7_75t_R FILLER_87_295 ();
 DECAPx4_ASAP7_75t_R FILLER_87_317 ();
 FILLER_ASAP7_75t_R FILLER_87_327 ();
 DECAPx1_ASAP7_75t_R FILLER_87_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_340 ();
 DECAPx10_ASAP7_75t_R FILLER_87_362 ();
 DECAPx4_ASAP7_75t_R FILLER_87_384 ();
 FILLER_ASAP7_75t_R FILLER_87_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_406 ();
 DECAPx6_ASAP7_75t_R FILLER_87_414 ();
 FILLER_ASAP7_75t_R FILLER_87_428 ();
 DECAPx2_ASAP7_75t_R FILLER_87_458 ();
 FILLER_ASAP7_75t_R FILLER_87_464 ();
 DECAPx10_ASAP7_75t_R FILLER_87_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_494 ();
 FILLER_ASAP7_75t_R FILLER_87_502 ();
 DECAPx2_ASAP7_75t_R FILLER_87_514 ();
 FILLER_ASAP7_75t_R FILLER_87_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_540 ();
 DECAPx1_ASAP7_75t_R FILLER_87_551 ();
 FILLER_ASAP7_75t_R FILLER_87_597 ();
 DECAPx10_ASAP7_75t_R FILLER_87_609 ();
 DECAPx10_ASAP7_75t_R FILLER_87_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_653 ();
 DECAPx10_ASAP7_75t_R FILLER_87_669 ();
 DECAPx6_ASAP7_75t_R FILLER_87_691 ();
 DECAPx1_ASAP7_75t_R FILLER_87_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_709 ();
 DECAPx10_ASAP7_75t_R FILLER_87_720 ();
 DECAPx10_ASAP7_75t_R FILLER_87_742 ();
 DECAPx4_ASAP7_75t_R FILLER_87_764 ();
 DECAPx10_ASAP7_75t_R FILLER_87_780 ();
 DECAPx10_ASAP7_75t_R FILLER_87_802 ();
 DECAPx2_ASAP7_75t_R FILLER_87_824 ();
 FILLER_ASAP7_75t_R FILLER_87_830 ();
 DECAPx10_ASAP7_75t_R FILLER_87_838 ();
 FILLER_ASAP7_75t_R FILLER_87_860 ();
 DECAPx10_ASAP7_75t_R FILLER_87_869 ();
 DECAPx10_ASAP7_75t_R FILLER_87_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_913 ();
 DECAPx10_ASAP7_75t_R FILLER_87_926 ();
 DECAPx10_ASAP7_75t_R FILLER_87_948 ();
 DECAPx10_ASAP7_75t_R FILLER_87_970 ();
 DECAPx1_ASAP7_75t_R FILLER_87_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_996 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1220 ();
 FILLER_ASAP7_75t_R FILLER_87_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1241 ();
 DECAPx6_ASAP7_75t_R FILLER_88_2 ();
 DECAPx2_ASAP7_75t_R FILLER_88_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_28 ();
 FILLER_ASAP7_75t_R FILLER_88_35 ();
 FILLER_ASAP7_75t_R FILLER_88_69 ();
 DECAPx2_ASAP7_75t_R FILLER_88_93 ();
 FILLER_ASAP7_75t_R FILLER_88_99 ();
 DECAPx1_ASAP7_75t_R FILLER_88_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_150 ();
 FILLER_ASAP7_75t_R FILLER_88_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_173 ();
 DECAPx1_ASAP7_75t_R FILLER_88_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_184 ();
 FILLER_ASAP7_75t_R FILLER_88_191 ();
 DECAPx4_ASAP7_75t_R FILLER_88_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_229 ();
 DECAPx2_ASAP7_75t_R FILLER_88_258 ();
 DECAPx10_ASAP7_75t_R FILLER_88_276 ();
 DECAPx6_ASAP7_75t_R FILLER_88_298 ();
 FILLER_ASAP7_75t_R FILLER_88_312 ();
 DECAPx6_ASAP7_75t_R FILLER_88_339 ();
 FILLER_ASAP7_75t_R FILLER_88_353 ();
 DECAPx2_ASAP7_75t_R FILLER_88_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_378 ();
 DECAPx6_ASAP7_75t_R FILLER_88_400 ();
 DECAPx2_ASAP7_75t_R FILLER_88_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_420 ();
 DECAPx10_ASAP7_75t_R FILLER_88_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_451 ();
 DECAPx6_ASAP7_75t_R FILLER_88_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_484 ();
 DECAPx10_ASAP7_75t_R FILLER_88_495 ();
 DECAPx2_ASAP7_75t_R FILLER_88_517 ();
 FILLER_ASAP7_75t_R FILLER_88_523 ();
 DECAPx1_ASAP7_75t_R FILLER_88_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_535 ();
 DECAPx10_ASAP7_75t_R FILLER_88_564 ();
 DECAPx2_ASAP7_75t_R FILLER_88_586 ();
 FILLER_ASAP7_75t_R FILLER_88_592 ();
 DECAPx1_ASAP7_75t_R FILLER_88_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_619 ();
 DECAPx10_ASAP7_75t_R FILLER_88_641 ();
 DECAPx10_ASAP7_75t_R FILLER_88_677 ();
 DECAPx10_ASAP7_75t_R FILLER_88_699 ();
 DECAPx10_ASAP7_75t_R FILLER_88_721 ();
 DECAPx10_ASAP7_75t_R FILLER_88_743 ();
 DECAPx6_ASAP7_75t_R FILLER_88_765 ();
 DECAPx1_ASAP7_75t_R FILLER_88_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_790 ();
 DECAPx10_ASAP7_75t_R FILLER_88_801 ();
 DECAPx6_ASAP7_75t_R FILLER_88_823 ();
 DECAPx4_ASAP7_75t_R FILLER_88_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_856 ();
 DECAPx1_ASAP7_75t_R FILLER_88_877 ();
 DECAPx10_ASAP7_75t_R FILLER_88_897 ();
 DECAPx2_ASAP7_75t_R FILLER_88_919 ();
 FILLER_ASAP7_75t_R FILLER_88_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_927 ();
 DECAPx6_ASAP7_75t_R FILLER_88_939 ();
 DECAPx2_ASAP7_75t_R FILLER_88_953 ();
 DECAPx10_ASAP7_75t_R FILLER_88_962 ();
 DECAPx1_ASAP7_75t_R FILLER_88_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_988 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1003 ();
 FILLER_ASAP7_75t_R FILLER_88_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1065 ();
 FILLER_ASAP7_75t_R FILLER_88_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1095 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1168 ();
 FILLER_ASAP7_75t_R FILLER_88_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1213 ();
 FILLER_ASAP7_75t_R FILLER_88_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1264 ();
 FILLER_ASAP7_75t_R FILLER_88_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1280 ();
 FILLER_ASAP7_75t_R FILLER_88_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_89_2 ();
 DECAPx2_ASAP7_75t_R FILLER_89_16 ();
 FILLER_ASAP7_75t_R FILLER_89_43 ();
 DECAPx4_ASAP7_75t_R FILLER_89_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_67 ();
 DECAPx2_ASAP7_75t_R FILLER_89_75 ();
 FILLER_ASAP7_75t_R FILLER_89_81 ();
 FILLER_ASAP7_75t_R FILLER_89_95 ();
 DECAPx1_ASAP7_75t_R FILLER_89_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_147 ();
 FILLER_ASAP7_75t_R FILLER_89_156 ();
 FILLER_ASAP7_75t_R FILLER_89_166 ();
 DECAPx6_ASAP7_75t_R FILLER_89_180 ();
 DECAPx1_ASAP7_75t_R FILLER_89_194 ();
 DECAPx10_ASAP7_75t_R FILLER_89_206 ();
 DECAPx2_ASAP7_75t_R FILLER_89_246 ();
 FILLER_ASAP7_75t_R FILLER_89_262 ();
 DECAPx2_ASAP7_75t_R FILLER_89_276 ();
 FILLER_ASAP7_75t_R FILLER_89_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_284 ();
 DECAPx10_ASAP7_75t_R FILLER_89_301 ();
 DECAPx4_ASAP7_75t_R FILLER_89_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_333 ();
 DECAPx2_ASAP7_75t_R FILLER_89_344 ();
 FILLER_ASAP7_75t_R FILLER_89_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_352 ();
 FILLER_ASAP7_75t_R FILLER_89_374 ();
 DECAPx1_ASAP7_75t_R FILLER_89_393 ();
 DECAPx1_ASAP7_75t_R FILLER_89_407 ();
 DECAPx2_ASAP7_75t_R FILLER_89_417 ();
 FILLER_ASAP7_75t_R FILLER_89_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_451 ();
 DECAPx6_ASAP7_75t_R FILLER_89_462 ();
 DECAPx1_ASAP7_75t_R FILLER_89_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_480 ();
 DECAPx10_ASAP7_75t_R FILLER_89_489 ();
 DECAPx2_ASAP7_75t_R FILLER_89_511 ();
 FILLER_ASAP7_75t_R FILLER_89_517 ();
 DECAPx10_ASAP7_75t_R FILLER_89_545 ();
 DECAPx4_ASAP7_75t_R FILLER_89_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_577 ();
 DECAPx4_ASAP7_75t_R FILLER_89_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_596 ();
 DECAPx6_ASAP7_75t_R FILLER_89_604 ();
 DECAPx2_ASAP7_75t_R FILLER_89_618 ();
 DECAPx1_ASAP7_75t_R FILLER_89_634 ();
 DECAPx2_ASAP7_75t_R FILLER_89_655 ();
 FILLER_ASAP7_75t_R FILLER_89_661 ();
 DECAPx4_ASAP7_75t_R FILLER_89_675 ();
 FILLER_ASAP7_75t_R FILLER_89_685 ();
 DECAPx10_ASAP7_75t_R FILLER_89_697 ();
 DECAPx10_ASAP7_75t_R FILLER_89_719 ();
 DECAPx6_ASAP7_75t_R FILLER_89_741 ();
 DECAPx1_ASAP7_75t_R FILLER_89_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_759 ();
 DECAPx1_ASAP7_75t_R FILLER_89_770 ();
 DECAPx10_ASAP7_75t_R FILLER_89_784 ();
 DECAPx10_ASAP7_75t_R FILLER_89_806 ();
 DECAPx10_ASAP7_75t_R FILLER_89_828 ();
 DECAPx10_ASAP7_75t_R FILLER_89_850 ();
 DECAPx10_ASAP7_75t_R FILLER_89_872 ();
 DECAPx10_ASAP7_75t_R FILLER_89_894 ();
 DECAPx2_ASAP7_75t_R FILLER_89_916 ();
 FILLER_ASAP7_75t_R FILLER_89_922 ();
 DECAPx2_ASAP7_75t_R FILLER_89_926 ();
 DECAPx6_ASAP7_75t_R FILLER_89_938 ();
 DECAPx1_ASAP7_75t_R FILLER_89_952 ();
 FILLER_ASAP7_75t_R FILLER_89_965 ();
 DECAPx6_ASAP7_75t_R FILLER_89_975 ();
 FILLER_ASAP7_75t_R FILLER_89_989 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1063 ();
 FILLER_ASAP7_75t_R FILLER_89_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1075 ();
 FILLER_ASAP7_75t_R FILLER_89_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1190 ();
 FILLER_ASAP7_75t_R FILLER_89_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1216 ();
 FILLER_ASAP7_75t_R FILLER_89_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1260 ();
 FILLER_ASAP7_75t_R FILLER_89_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_89_1280 ();
 FILLER_ASAP7_75t_R FILLER_89_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_90_2 ();
 DECAPx2_ASAP7_75t_R FILLER_90_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_38 ();
 FILLER_ASAP7_75t_R FILLER_90_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_55 ();
 DECAPx2_ASAP7_75t_R FILLER_90_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_69 ();
 DECAPx6_ASAP7_75t_R FILLER_90_77 ();
 DECAPx2_ASAP7_75t_R FILLER_90_91 ();
 DECAPx4_ASAP7_75t_R FILLER_90_105 ();
 FILLER_ASAP7_75t_R FILLER_90_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_124 ();
 DECAPx1_ASAP7_75t_R FILLER_90_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_166 ();
 DECAPx1_ASAP7_75t_R FILLER_90_181 ();
 DECAPx10_ASAP7_75t_R FILLER_90_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_231 ();
 DECAPx10_ASAP7_75t_R FILLER_90_252 ();
 DECAPx10_ASAP7_75t_R FILLER_90_274 ();
 DECAPx10_ASAP7_75t_R FILLER_90_296 ();
 DECAPx2_ASAP7_75t_R FILLER_90_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_324 ();
 FILLER_ASAP7_75t_R FILLER_90_411 ();
 DECAPx1_ASAP7_75t_R FILLER_90_425 ();
 DECAPx2_ASAP7_75t_R FILLER_90_435 ();
 DECAPx10_ASAP7_75t_R FILLER_90_464 ();
 DECAPx2_ASAP7_75t_R FILLER_90_486 ();
 DECAPx1_ASAP7_75t_R FILLER_90_502 ();
 FILLER_ASAP7_75t_R FILLER_90_513 ();
 FILLER_ASAP7_75t_R FILLER_90_525 ();
 FILLER_ASAP7_75t_R FILLER_90_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_535 ();
 FILLER_ASAP7_75t_R FILLER_90_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_545 ();
 DECAPx4_ASAP7_75t_R FILLER_90_567 ();
 FILLER_ASAP7_75t_R FILLER_90_577 ();
 DECAPx1_ASAP7_75t_R FILLER_90_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_593 ();
 DECAPx6_ASAP7_75t_R FILLER_90_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_643 ();
 DECAPx10_ASAP7_75t_R FILLER_90_686 ();
 DECAPx1_ASAP7_75t_R FILLER_90_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_712 ();
 DECAPx10_ASAP7_75t_R FILLER_90_719 ();
 DECAPx6_ASAP7_75t_R FILLER_90_741 ();
 DECAPx6_ASAP7_75t_R FILLER_90_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_777 ();
 DECAPx10_ASAP7_75t_R FILLER_90_784 ();
 DECAPx10_ASAP7_75t_R FILLER_90_806 ();
 DECAPx10_ASAP7_75t_R FILLER_90_828 ();
 DECAPx10_ASAP7_75t_R FILLER_90_850 ();
 DECAPx10_ASAP7_75t_R FILLER_90_872 ();
 DECAPx10_ASAP7_75t_R FILLER_90_894 ();
 DECAPx10_ASAP7_75t_R FILLER_90_916 ();
 DECAPx2_ASAP7_75t_R FILLER_90_938 ();
 FILLER_ASAP7_75t_R FILLER_90_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_946 ();
 DECAPx10_ASAP7_75t_R FILLER_90_959 ();
 DECAPx10_ASAP7_75t_R FILLER_90_981 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1025 ();
 FILLER_ASAP7_75t_R FILLER_90_1037 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1163 ();
 FILLER_ASAP7_75t_R FILLER_90_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1204 ();
 FILLER_ASAP7_75t_R FILLER_90_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_90_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1247 ();
 DECAPx6_ASAP7_75t_R FILLER_91_2 ();
 DECAPx1_ASAP7_75t_R FILLER_91_16 ();
 DECAPx1_ASAP7_75t_R FILLER_91_26 ();
 FILLER_ASAP7_75t_R FILLER_91_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_39 ();
 DECAPx6_ASAP7_75t_R FILLER_91_52 ();
 DECAPx2_ASAP7_75t_R FILLER_91_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_72 ();
 DECAPx1_ASAP7_75t_R FILLER_91_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_84 ();
 DECAPx10_ASAP7_75t_R FILLER_91_101 ();
 DECAPx6_ASAP7_75t_R FILLER_91_123 ();
 FILLER_ASAP7_75t_R FILLER_91_137 ();
 DECAPx1_ASAP7_75t_R FILLER_91_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_171 ();
 FILLER_ASAP7_75t_R FILLER_91_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_180 ();
 FILLER_ASAP7_75t_R FILLER_91_203 ();
 FILLER_ASAP7_75t_R FILLER_91_211 ();
 FILLER_ASAP7_75t_R FILLER_91_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_231 ();
 DECAPx4_ASAP7_75t_R FILLER_91_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_262 ();
 DECAPx2_ASAP7_75t_R FILLER_91_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_281 ();
 DECAPx10_ASAP7_75t_R FILLER_91_300 ();
 DECAPx6_ASAP7_75t_R FILLER_91_322 ();
 DECAPx2_ASAP7_75t_R FILLER_91_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_364 ();
 FILLER_ASAP7_75t_R FILLER_91_386 ();
 DECAPx6_ASAP7_75t_R FILLER_91_422 ();
 FILLER_ASAP7_75t_R FILLER_91_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_438 ();
 DECAPx10_ASAP7_75t_R FILLER_91_461 ();
 FILLER_ASAP7_75t_R FILLER_91_483 ();
 DECAPx4_ASAP7_75t_R FILLER_91_533 ();
 FILLER_ASAP7_75t_R FILLER_91_543 ();
 DECAPx6_ASAP7_75t_R FILLER_91_562 ();
 DECAPx6_ASAP7_75t_R FILLER_91_582 ();
 FILLER_ASAP7_75t_R FILLER_91_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_598 ();
 DECAPx10_ASAP7_75t_R FILLER_91_609 ();
 FILLER_ASAP7_75t_R FILLER_91_631 ();
 DECAPx6_ASAP7_75t_R FILLER_91_643 ();
 DECAPx2_ASAP7_75t_R FILLER_91_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_663 ();
 DECAPx10_ASAP7_75t_R FILLER_91_674 ();
 DECAPx6_ASAP7_75t_R FILLER_91_696 ();
 FILLER_ASAP7_75t_R FILLER_91_710 ();
 DECAPx4_ASAP7_75t_R FILLER_91_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_728 ();
 DECAPx10_ASAP7_75t_R FILLER_91_735 ();
 DECAPx10_ASAP7_75t_R FILLER_91_757 ();
 DECAPx10_ASAP7_75t_R FILLER_91_779 ();
 DECAPx10_ASAP7_75t_R FILLER_91_801 ();
 DECAPx10_ASAP7_75t_R FILLER_91_823 ();
 DECAPx10_ASAP7_75t_R FILLER_91_845 ();
 DECAPx10_ASAP7_75t_R FILLER_91_867 ();
 DECAPx1_ASAP7_75t_R FILLER_91_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_893 ();
 DECAPx10_ASAP7_75t_R FILLER_91_900 ();
 FILLER_ASAP7_75t_R FILLER_91_922 ();
 DECAPx10_ASAP7_75t_R FILLER_91_926 ();
 DECAPx10_ASAP7_75t_R FILLER_91_948 ();
 DECAPx10_ASAP7_75t_R FILLER_91_970 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1204 ();
 FILLER_ASAP7_75t_R FILLER_91_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1272 ();
 FILLER_ASAP7_75t_R FILLER_91_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1280 ();
 FILLER_ASAP7_75t_R FILLER_91_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_92_2 ();
 DECAPx4_ASAP7_75t_R FILLER_92_24 ();
 DECAPx2_ASAP7_75t_R FILLER_92_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_47 ();
 DECAPx1_ASAP7_75t_R FILLER_92_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_58 ();
 DECAPx6_ASAP7_75t_R FILLER_92_82 ();
 FILLER_ASAP7_75t_R FILLER_92_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_110 ();
 DECAPx1_ASAP7_75t_R FILLER_92_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_121 ();
 DECAPx1_ASAP7_75t_R FILLER_92_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_134 ();
 DECAPx10_ASAP7_75t_R FILLER_92_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_176 ();
 DECAPx4_ASAP7_75t_R FILLER_92_193 ();
 DECAPx4_ASAP7_75t_R FILLER_92_209 ();
 DECAPx4_ASAP7_75t_R FILLER_92_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_243 ();
 DECAPx6_ASAP7_75t_R FILLER_92_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_272 ();
 DECAPx4_ASAP7_75t_R FILLER_92_283 ();
 FILLER_ASAP7_75t_R FILLER_92_293 ();
 DECAPx4_ASAP7_75t_R FILLER_92_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_326 ();
 DECAPx2_ASAP7_75t_R FILLER_92_333 ();
 DECAPx2_ASAP7_75t_R FILLER_92_360 ();
 FILLER_ASAP7_75t_R FILLER_92_366 ();
 DECAPx1_ASAP7_75t_R FILLER_92_412 ();
 DECAPx6_ASAP7_75t_R FILLER_92_423 ();
 FILLER_ASAP7_75t_R FILLER_92_443 ();
 FILLER_ASAP7_75t_R FILLER_92_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_454 ();
 DECAPx1_ASAP7_75t_R FILLER_92_485 ();
 DECAPx6_ASAP7_75t_R FILLER_92_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_510 ();
 FILLER_ASAP7_75t_R FILLER_92_518 ();
 DECAPx10_ASAP7_75t_R FILLER_92_530 ();
 DECAPx10_ASAP7_75t_R FILLER_92_552 ();
 DECAPx10_ASAP7_75t_R FILLER_92_574 ();
 DECAPx1_ASAP7_75t_R FILLER_92_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_600 ();
 DECAPx10_ASAP7_75t_R FILLER_92_608 ();
 DECAPx10_ASAP7_75t_R FILLER_92_630 ();
 DECAPx4_ASAP7_75t_R FILLER_92_652 ();
 FILLER_ASAP7_75t_R FILLER_92_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_664 ();
 DECAPx10_ASAP7_75t_R FILLER_92_672 ();
 DECAPx10_ASAP7_75t_R FILLER_92_694 ();
 DECAPx6_ASAP7_75t_R FILLER_92_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_730 ();
 DECAPx10_ASAP7_75t_R FILLER_92_737 ();
 DECAPx10_ASAP7_75t_R FILLER_92_759 ();
 DECAPx10_ASAP7_75t_R FILLER_92_781 ();
 DECAPx1_ASAP7_75t_R FILLER_92_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_807 ();
 DECAPx6_ASAP7_75t_R FILLER_92_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_828 ();
 DECAPx10_ASAP7_75t_R FILLER_92_841 ();
 DECAPx10_ASAP7_75t_R FILLER_92_863 ();
 DECAPx2_ASAP7_75t_R FILLER_92_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_891 ();
 DECAPx10_ASAP7_75t_R FILLER_92_906 ();
 DECAPx10_ASAP7_75t_R FILLER_92_928 ();
 DECAPx10_ASAP7_75t_R FILLER_92_950 ();
 DECAPx10_ASAP7_75t_R FILLER_92_972 ();
 DECAPx6_ASAP7_75t_R FILLER_92_994 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_92_1084 ();
 FILLER_ASAP7_75t_R FILLER_92_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1167 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1191 ();
 FILLER_ASAP7_75t_R FILLER_92_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1199 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1280 ();
 FILLER_ASAP7_75t_R FILLER_92_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_93_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_16 ();
 DECAPx2_ASAP7_75t_R FILLER_93_39 ();
 FILLER_ASAP7_75t_R FILLER_93_45 ();
 DECAPx4_ASAP7_75t_R FILLER_93_57 ();
 FILLER_ASAP7_75t_R FILLER_93_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_69 ();
 FILLER_ASAP7_75t_R FILLER_93_84 ();
 FILLER_ASAP7_75t_R FILLER_93_92 ();
 DECAPx4_ASAP7_75t_R FILLER_93_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_111 ();
 DECAPx1_ASAP7_75t_R FILLER_93_126 ();
 DECAPx1_ASAP7_75t_R FILLER_93_136 ();
 DECAPx2_ASAP7_75t_R FILLER_93_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_152 ();
 DECAPx2_ASAP7_75t_R FILLER_93_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_167 ();
 DECAPx1_ASAP7_75t_R FILLER_93_176 ();
 FILLER_ASAP7_75t_R FILLER_93_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_195 ();
 DECAPx4_ASAP7_75t_R FILLER_93_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_213 ();
 DECAPx10_ASAP7_75t_R FILLER_93_230 ();
 DECAPx10_ASAP7_75t_R FILLER_93_252 ();
 DECAPx2_ASAP7_75t_R FILLER_93_274 ();
 FILLER_ASAP7_75t_R FILLER_93_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_282 ();
 DECAPx10_ASAP7_75t_R FILLER_93_303 ();
 DECAPx1_ASAP7_75t_R FILLER_93_325 ();
 FILLER_ASAP7_75t_R FILLER_93_336 ();
 DECAPx6_ASAP7_75t_R FILLER_93_348 ();
 FILLER_ASAP7_75t_R FILLER_93_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_374 ();
 FILLER_ASAP7_75t_R FILLER_93_383 ();
 FILLER_ASAP7_75t_R FILLER_93_395 ();
 DECAPx1_ASAP7_75t_R FILLER_93_404 ();
 DECAPx2_ASAP7_75t_R FILLER_93_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_435 ();
 DECAPx2_ASAP7_75t_R FILLER_93_442 ();
 FILLER_ASAP7_75t_R FILLER_93_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_450 ();
 DECAPx2_ASAP7_75t_R FILLER_93_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_477 ();
 DECAPx4_ASAP7_75t_R FILLER_93_499 ();
 DECAPx10_ASAP7_75t_R FILLER_93_530 ();
 DECAPx6_ASAP7_75t_R FILLER_93_562 ();
 DECAPx10_ASAP7_75t_R FILLER_93_588 ();
 DECAPx10_ASAP7_75t_R FILLER_93_610 ();
 DECAPx10_ASAP7_75t_R FILLER_93_632 ();
 DECAPx2_ASAP7_75t_R FILLER_93_654 ();
 DECAPx4_ASAP7_75t_R FILLER_93_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_680 ();
 DECAPx2_ASAP7_75t_R FILLER_93_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_697 ();
 DECAPx4_ASAP7_75t_R FILLER_93_704 ();
 DECAPx10_ASAP7_75t_R FILLER_93_724 ();
 DECAPx1_ASAP7_75t_R FILLER_93_746 ();
 DECAPx10_ASAP7_75t_R FILLER_93_764 ();
 DECAPx10_ASAP7_75t_R FILLER_93_786 ();
 DECAPx10_ASAP7_75t_R FILLER_93_808 ();
 FILLER_ASAP7_75t_R FILLER_93_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_832 ();
 DECAPx10_ASAP7_75t_R FILLER_93_839 ();
 DECAPx10_ASAP7_75t_R FILLER_93_861 ();
 DECAPx10_ASAP7_75t_R FILLER_93_883 ();
 DECAPx6_ASAP7_75t_R FILLER_93_905 ();
 DECAPx1_ASAP7_75t_R FILLER_93_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_923 ();
 DECAPx10_ASAP7_75t_R FILLER_93_926 ();
 DECAPx10_ASAP7_75t_R FILLER_93_948 ();
 DECAPx2_ASAP7_75t_R FILLER_93_970 ();
 FILLER_ASAP7_75t_R FILLER_93_976 ();
 DECAPx2_ASAP7_75t_R FILLER_93_984 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_93_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1144 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1192 ();
 FILLER_ASAP7_75t_R FILLER_93_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1206 ();
 FILLER_ASAP7_75t_R FILLER_93_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1247 ();
 FILLER_ASAP7_75t_R FILLER_93_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1277 ();
 FILLER_ASAP7_75t_R FILLER_93_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_94_2 ();
 FILLER_ASAP7_75t_R FILLER_94_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_23 ();
 DECAPx4_ASAP7_75t_R FILLER_94_42 ();
 FILLER_ASAP7_75t_R FILLER_94_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_60 ();
 DECAPx6_ASAP7_75t_R FILLER_94_73 ();
 DECAPx1_ASAP7_75t_R FILLER_94_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_91 ();
 DECAPx2_ASAP7_75t_R FILLER_94_106 ();
 FILLER_ASAP7_75t_R FILLER_94_122 ();
 DECAPx4_ASAP7_75t_R FILLER_94_139 ();
 DECAPx4_ASAP7_75t_R FILLER_94_157 ();
 DECAPx6_ASAP7_75t_R FILLER_94_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_189 ();
 FILLER_ASAP7_75t_R FILLER_94_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_222 ();
 FILLER_ASAP7_75t_R FILLER_94_229 ();
 FILLER_ASAP7_75t_R FILLER_94_241 ();
 DECAPx2_ASAP7_75t_R FILLER_94_255 ();
 FILLER_ASAP7_75t_R FILLER_94_261 ();
 DECAPx4_ASAP7_75t_R FILLER_94_275 ();
 FILLER_ASAP7_75t_R FILLER_94_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_302 ();
 DECAPx6_ASAP7_75t_R FILLER_94_309 ();
 FILLER_ASAP7_75t_R FILLER_94_323 ();
 FILLER_ASAP7_75t_R FILLER_94_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_348 ();
 DECAPx1_ASAP7_75t_R FILLER_94_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_374 ();
 DECAPx1_ASAP7_75t_R FILLER_94_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_400 ();
 DECAPx1_ASAP7_75t_R FILLER_94_411 ();
 DECAPx1_ASAP7_75t_R FILLER_94_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_435 ();
 DECAPx4_ASAP7_75t_R FILLER_94_452 ();
 DECAPx2_ASAP7_75t_R FILLER_94_464 ();
 FILLER_ASAP7_75t_R FILLER_94_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_472 ();
 DECAPx4_ASAP7_75t_R FILLER_94_490 ();
 DECAPx2_ASAP7_75t_R FILLER_94_510 ();
 DECAPx10_ASAP7_75t_R FILLER_94_523 ();
 DECAPx2_ASAP7_75t_R FILLER_94_545 ();
 DECAPx2_ASAP7_75t_R FILLER_94_557 ();
 DECAPx6_ASAP7_75t_R FILLER_94_570 ();
 DECAPx6_ASAP7_75t_R FILLER_94_590 ();
 FILLER_ASAP7_75t_R FILLER_94_604 ();
 DECAPx10_ASAP7_75t_R FILLER_94_612 ();
 DECAPx2_ASAP7_75t_R FILLER_94_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_640 ();
 DECAPx10_ASAP7_75t_R FILLER_94_651 ();
 DECAPx6_ASAP7_75t_R FILLER_94_683 ();
 FILLER_ASAP7_75t_R FILLER_94_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_699 ();
 DECAPx1_ASAP7_75t_R FILLER_94_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_710 ();
 DECAPx10_ASAP7_75t_R FILLER_94_717 ();
 DECAPx10_ASAP7_75t_R FILLER_94_739 ();
 DECAPx10_ASAP7_75t_R FILLER_94_761 ();
 DECAPx6_ASAP7_75t_R FILLER_94_783 ();
 DECAPx1_ASAP7_75t_R FILLER_94_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_801 ();
 DECAPx10_ASAP7_75t_R FILLER_94_808 ();
 DECAPx10_ASAP7_75t_R FILLER_94_830 ();
 DECAPx6_ASAP7_75t_R FILLER_94_852 ();
 FILLER_ASAP7_75t_R FILLER_94_866 ();
 DECAPx4_ASAP7_75t_R FILLER_94_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_888 ();
 DECAPx6_ASAP7_75t_R FILLER_94_899 ();
 DECAPx10_ASAP7_75t_R FILLER_94_927 ();
 DECAPx4_ASAP7_75t_R FILLER_94_949 ();
 DECAPx2_ASAP7_75t_R FILLER_94_975 ();
 DECAPx1_ASAP7_75t_R FILLER_94_998 ();
 FILLER_ASAP7_75t_R FILLER_94_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1021 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1053 ();
 FILLER_ASAP7_75t_R FILLER_94_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1150 ();
 FILLER_ASAP7_75t_R FILLER_94_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1179 ();
 FILLER_ASAP7_75t_R FILLER_94_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1222 ();
 FILLER_ASAP7_75t_R FILLER_94_1228 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_95_2 ();
 FILLER_ASAP7_75t_R FILLER_95_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_27 ();
 DECAPx2_ASAP7_75t_R FILLER_95_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_50 ();
 DECAPx1_ASAP7_75t_R FILLER_95_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_61 ();
 DECAPx4_ASAP7_75t_R FILLER_95_105 ();
 FILLER_ASAP7_75t_R FILLER_95_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_117 ();
 FILLER_ASAP7_75t_R FILLER_95_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_143 ();
 FILLER_ASAP7_75t_R FILLER_95_166 ();
 DECAPx4_ASAP7_75t_R FILLER_95_176 ();
 FILLER_ASAP7_75t_R FILLER_95_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_188 ();
 DECAPx6_ASAP7_75t_R FILLER_95_209 ();
 DECAPx2_ASAP7_75t_R FILLER_95_223 ();
 DECAPx10_ASAP7_75t_R FILLER_95_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_281 ();
 DECAPx1_ASAP7_75t_R FILLER_95_296 ();
 DECAPx10_ASAP7_75t_R FILLER_95_311 ();
 DECAPx4_ASAP7_75t_R FILLER_95_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_343 ();
 DECAPx2_ASAP7_75t_R FILLER_95_382 ();
 FILLER_ASAP7_75t_R FILLER_95_388 ();
 DECAPx6_ASAP7_75t_R FILLER_95_407 ();
 DECAPx2_ASAP7_75t_R FILLER_95_433 ();
 DECAPx2_ASAP7_75t_R FILLER_95_482 ();
 FILLER_ASAP7_75t_R FILLER_95_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_490 ();
 DECAPx10_ASAP7_75t_R FILLER_95_518 ();
 DECAPx6_ASAP7_75t_R FILLER_95_540 ();
 DECAPx1_ASAP7_75t_R FILLER_95_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_558 ();
 FILLER_ASAP7_75t_R FILLER_95_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_567 ();
 DECAPx10_ASAP7_75t_R FILLER_95_575 ();
 DECAPx10_ASAP7_75t_R FILLER_95_597 ();
 DECAPx10_ASAP7_75t_R FILLER_95_619 ();
 DECAPx6_ASAP7_75t_R FILLER_95_641 ();
 DECAPx1_ASAP7_75t_R FILLER_95_655 ();
 DECAPx2_ASAP7_75t_R FILLER_95_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_701 ();
 DECAPx10_ASAP7_75t_R FILLER_95_709 ();
 DECAPx10_ASAP7_75t_R FILLER_95_731 ();
 DECAPx10_ASAP7_75t_R FILLER_95_753 ();
 DECAPx10_ASAP7_75t_R FILLER_95_775 ();
 DECAPx2_ASAP7_75t_R FILLER_95_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_803 ();
 DECAPx10_ASAP7_75t_R FILLER_95_814 ();
 DECAPx10_ASAP7_75t_R FILLER_95_836 ();
 DECAPx10_ASAP7_75t_R FILLER_95_858 ();
 DECAPx2_ASAP7_75t_R FILLER_95_880 ();
 DECAPx10_ASAP7_75t_R FILLER_95_900 ();
 FILLER_ASAP7_75t_R FILLER_95_922 ();
 DECAPx10_ASAP7_75t_R FILLER_95_926 ();
 DECAPx10_ASAP7_75t_R FILLER_95_948 ();
 DECAPx10_ASAP7_75t_R FILLER_95_970 ();
 DECAPx10_ASAP7_75t_R FILLER_95_992 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1112 ();
 FILLER_ASAP7_75t_R FILLER_95_1118 ();
 FILLER_ASAP7_75t_R FILLER_95_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1129 ();
 FILLER_ASAP7_75t_R FILLER_95_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1161 ();
 FILLER_ASAP7_75t_R FILLER_95_1175 ();
 FILLER_ASAP7_75t_R FILLER_95_1213 ();
 DECAPx4_ASAP7_75t_R FILLER_95_1221 ();
 FILLER_ASAP7_75t_R FILLER_95_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1233 ();
 FILLER_ASAP7_75t_R FILLER_95_1251 ();
 DECAPx4_ASAP7_75t_R FILLER_95_1260 ();
 FILLER_ASAP7_75t_R FILLER_95_1270 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_96_2 ();
 DECAPx1_ASAP7_75t_R FILLER_96_19 ();
 DECAPx2_ASAP7_75t_R FILLER_96_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_56 ();
 DECAPx1_ASAP7_75t_R FILLER_96_67 ();
 DECAPx4_ASAP7_75t_R FILLER_96_77 ();
 FILLER_ASAP7_75t_R FILLER_96_87 ();
 DECAPx6_ASAP7_75t_R FILLER_96_95 ();
 DECAPx1_ASAP7_75t_R FILLER_96_109 ();
 DECAPx2_ASAP7_75t_R FILLER_96_119 ();
 FILLER_ASAP7_75t_R FILLER_96_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_139 ();
 DECAPx4_ASAP7_75t_R FILLER_96_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_173 ();
 FILLER_ASAP7_75t_R FILLER_96_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_191 ();
 FILLER_ASAP7_75t_R FILLER_96_198 ();
 DECAPx6_ASAP7_75t_R FILLER_96_214 ();
 FILLER_ASAP7_75t_R FILLER_96_228 ();
 DECAPx10_ASAP7_75t_R FILLER_96_240 ();
 DECAPx10_ASAP7_75t_R FILLER_96_262 ();
 FILLER_ASAP7_75t_R FILLER_96_298 ();
 FILLER_ASAP7_75t_R FILLER_96_310 ();
 FILLER_ASAP7_75t_R FILLER_96_329 ();
 DECAPx10_ASAP7_75t_R FILLER_96_347 ();
 DECAPx4_ASAP7_75t_R FILLER_96_369 ();
 FILLER_ASAP7_75t_R FILLER_96_379 ();
 DECAPx6_ASAP7_75t_R FILLER_96_402 ();
 DECAPx1_ASAP7_75t_R FILLER_96_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_420 ();
 DECAPx10_ASAP7_75t_R FILLER_96_427 ();
 DECAPx2_ASAP7_75t_R FILLER_96_449 ();
 FILLER_ASAP7_75t_R FILLER_96_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_494 ();
 DECAPx1_ASAP7_75t_R FILLER_96_502 ();
 DECAPx10_ASAP7_75t_R FILLER_96_524 ();
 DECAPx10_ASAP7_75t_R FILLER_96_546 ();
 DECAPx4_ASAP7_75t_R FILLER_96_568 ();
 FILLER_ASAP7_75t_R FILLER_96_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_580 ();
 DECAPx10_ASAP7_75t_R FILLER_96_591 ();
 DECAPx10_ASAP7_75t_R FILLER_96_613 ();
 DECAPx6_ASAP7_75t_R FILLER_96_635 ();
 DECAPx2_ASAP7_75t_R FILLER_96_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_655 ();
 DECAPx10_ASAP7_75t_R FILLER_96_666 ();
 DECAPx2_ASAP7_75t_R FILLER_96_688 ();
 FILLER_ASAP7_75t_R FILLER_96_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_696 ();
 DECAPx10_ASAP7_75t_R FILLER_96_707 ();
 DECAPx2_ASAP7_75t_R FILLER_96_729 ();
 DECAPx10_ASAP7_75t_R FILLER_96_741 ();
 DECAPx10_ASAP7_75t_R FILLER_96_763 ();
 DECAPx10_ASAP7_75t_R FILLER_96_785 ();
 DECAPx10_ASAP7_75t_R FILLER_96_807 ();
 DECAPx10_ASAP7_75t_R FILLER_96_829 ();
 DECAPx4_ASAP7_75t_R FILLER_96_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_861 ();
 DECAPx10_ASAP7_75t_R FILLER_96_868 ();
 DECAPx10_ASAP7_75t_R FILLER_96_890 ();
 DECAPx4_ASAP7_75t_R FILLER_96_912 ();
 FILLER_ASAP7_75t_R FILLER_96_922 ();
 DECAPx6_ASAP7_75t_R FILLER_96_934 ();
 FILLER_ASAP7_75t_R FILLER_96_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_950 ();
 DECAPx2_ASAP7_75t_R FILLER_96_957 ();
 FILLER_ASAP7_75t_R FILLER_96_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_965 ();
 DECAPx10_ASAP7_75t_R FILLER_96_976 ();
 DECAPx1_ASAP7_75t_R FILLER_96_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1060 ();
 FILLER_ASAP7_75t_R FILLER_96_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1110 ();
 FILLER_ASAP7_75t_R FILLER_96_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1156 ();
 FILLER_ASAP7_75t_R FILLER_96_1165 ();
 FILLER_ASAP7_75t_R FILLER_96_1175 ();
 FILLER_ASAP7_75t_R FILLER_96_1187 ();
 FILLER_ASAP7_75t_R FILLER_96_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1231 ();
 FILLER_ASAP7_75t_R FILLER_96_1245 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_97_2 ();
 FILLER_ASAP7_75t_R FILLER_97_8 ();
 FILLER_ASAP7_75t_R FILLER_97_37 ();
 FILLER_ASAP7_75t_R FILLER_97_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_56 ();
 FILLER_ASAP7_75t_R FILLER_97_65 ();
 FILLER_ASAP7_75t_R FILLER_97_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_77 ();
 FILLER_ASAP7_75t_R FILLER_97_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_90 ();
 FILLER_ASAP7_75t_R FILLER_97_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_99 ();
 DECAPx6_ASAP7_75t_R FILLER_97_106 ();
 FILLER_ASAP7_75t_R FILLER_97_120 ();
 DECAPx4_ASAP7_75t_R FILLER_97_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_147 ();
 DECAPx4_ASAP7_75t_R FILLER_97_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_166 ();
 DECAPx2_ASAP7_75t_R FILLER_97_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_180 ();
 DECAPx2_ASAP7_75t_R FILLER_97_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_194 ();
 DECAPx10_ASAP7_75t_R FILLER_97_202 ();
 DECAPx6_ASAP7_75t_R FILLER_97_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_238 ();
 DECAPx6_ASAP7_75t_R FILLER_97_259 ();
 DECAPx2_ASAP7_75t_R FILLER_97_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_310 ();
 FILLER_ASAP7_75t_R FILLER_97_317 ();
 DECAPx10_ASAP7_75t_R FILLER_97_327 ();
 DECAPx10_ASAP7_75t_R FILLER_97_349 ();
 DECAPx4_ASAP7_75t_R FILLER_97_371 ();
 DECAPx2_ASAP7_75t_R FILLER_97_402 ();
 FILLER_ASAP7_75t_R FILLER_97_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_410 ();
 DECAPx1_ASAP7_75t_R FILLER_97_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_432 ();
 DECAPx6_ASAP7_75t_R FILLER_97_490 ();
 DECAPx1_ASAP7_75t_R FILLER_97_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_508 ();
 DECAPx4_ASAP7_75t_R FILLER_97_527 ();
 FILLER_ASAP7_75t_R FILLER_97_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_539 ();
 FILLER_ASAP7_75t_R FILLER_97_554 ();
 DECAPx10_ASAP7_75t_R FILLER_97_565 ();
 DECAPx6_ASAP7_75t_R FILLER_97_587 ();
 FILLER_ASAP7_75t_R FILLER_97_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_603 ();
 DECAPx6_ASAP7_75t_R FILLER_97_621 ();
 FILLER_ASAP7_75t_R FILLER_97_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_637 ();
 DECAPx1_ASAP7_75t_R FILLER_97_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_648 ();
 DECAPx10_ASAP7_75t_R FILLER_97_661 ();
 DECAPx6_ASAP7_75t_R FILLER_97_683 ();
 FILLER_ASAP7_75t_R FILLER_97_697 ();
 FILLER_ASAP7_75t_R FILLER_97_728 ();
 DECAPx10_ASAP7_75t_R FILLER_97_740 ();
 FILLER_ASAP7_75t_R FILLER_97_762 ();
 DECAPx10_ASAP7_75t_R FILLER_97_780 ();
 DECAPx10_ASAP7_75t_R FILLER_97_802 ();
 DECAPx2_ASAP7_75t_R FILLER_97_824 ();
 FILLER_ASAP7_75t_R FILLER_97_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_832 ();
 DECAPx10_ASAP7_75t_R FILLER_97_847 ();
 DECAPx10_ASAP7_75t_R FILLER_97_869 ();
 DECAPx6_ASAP7_75t_R FILLER_97_891 ();
 DECAPx4_ASAP7_75t_R FILLER_97_911 ();
 FILLER_ASAP7_75t_R FILLER_97_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_923 ();
 DECAPx6_ASAP7_75t_R FILLER_97_926 ();
 DECAPx1_ASAP7_75t_R FILLER_97_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_944 ();
 DECAPx10_ASAP7_75t_R FILLER_97_959 ();
 FILLER_ASAP7_75t_R FILLER_97_981 ();
 DECAPx2_ASAP7_75t_R FILLER_97_993 ();
 FILLER_ASAP7_75t_R FILLER_97_999 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1203 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1254 ();
 FILLER_ASAP7_75t_R FILLER_97_1260 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_98_2 ();
 FILLER_ASAP7_75t_R FILLER_98_8 ();
 FILLER_ASAP7_75t_R FILLER_98_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_28 ();
 DECAPx2_ASAP7_75t_R FILLER_98_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_67 ();
 DECAPx2_ASAP7_75t_R FILLER_98_74 ();
 FILLER_ASAP7_75t_R FILLER_98_80 ();
 DECAPx1_ASAP7_75t_R FILLER_98_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_99 ();
 DECAPx4_ASAP7_75t_R FILLER_98_122 ();
 DECAPx10_ASAP7_75t_R FILLER_98_147 ();
 FILLER_ASAP7_75t_R FILLER_98_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_194 ();
 DECAPx2_ASAP7_75t_R FILLER_98_201 ();
 FILLER_ASAP7_75t_R FILLER_98_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_209 ();
 DECAPx4_ASAP7_75t_R FILLER_98_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_230 ();
 DECAPx10_ASAP7_75t_R FILLER_98_241 ();
 FILLER_ASAP7_75t_R FILLER_98_263 ();
 FILLER_ASAP7_75t_R FILLER_98_287 ();
 DECAPx1_ASAP7_75t_R FILLER_98_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_299 ();
 FILLER_ASAP7_75t_R FILLER_98_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_309 ();
 FILLER_ASAP7_75t_R FILLER_98_318 ();
 FILLER_ASAP7_75t_R FILLER_98_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_328 ();
 FILLER_ASAP7_75t_R FILLER_98_335 ();
 DECAPx1_ASAP7_75t_R FILLER_98_345 ();
 DECAPx4_ASAP7_75t_R FILLER_98_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_365 ();
 DECAPx1_ASAP7_75t_R FILLER_98_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_380 ();
 DECAPx2_ASAP7_75t_R FILLER_98_388 ();
 FILLER_ASAP7_75t_R FILLER_98_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_396 ();
 FILLER_ASAP7_75t_R FILLER_98_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_409 ();
 DECAPx6_ASAP7_75t_R FILLER_98_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_445 ();
 DECAPx2_ASAP7_75t_R FILLER_98_456 ();
 DECAPx1_ASAP7_75t_R FILLER_98_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_476 ();
 DECAPx4_ASAP7_75t_R FILLER_98_498 ();
 FILLER_ASAP7_75t_R FILLER_98_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_510 ();
 DECAPx10_ASAP7_75t_R FILLER_98_533 ();
 DECAPx10_ASAP7_75t_R FILLER_98_555 ();
 DECAPx2_ASAP7_75t_R FILLER_98_577 ();
 FILLER_ASAP7_75t_R FILLER_98_583 ();
 DECAPx10_ASAP7_75t_R FILLER_98_591 ();
 DECAPx1_ASAP7_75t_R FILLER_98_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_668 ();
 DECAPx4_ASAP7_75t_R FILLER_98_690 ();
 FILLER_ASAP7_75t_R FILLER_98_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_731 ();
 DECAPx10_ASAP7_75t_R FILLER_98_738 ();
 DECAPx10_ASAP7_75t_R FILLER_98_760 ();
 DECAPx6_ASAP7_75t_R FILLER_98_782 ();
 DECAPx2_ASAP7_75t_R FILLER_98_796 ();
 DECAPx10_ASAP7_75t_R FILLER_98_812 ();
 DECAPx10_ASAP7_75t_R FILLER_98_834 ();
 DECAPx10_ASAP7_75t_R FILLER_98_856 ();
 DECAPx6_ASAP7_75t_R FILLER_98_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_892 ();
 DECAPx2_ASAP7_75t_R FILLER_98_901 ();
 DECAPx10_ASAP7_75t_R FILLER_98_913 ();
 DECAPx10_ASAP7_75t_R FILLER_98_935 ();
 DECAPx10_ASAP7_75t_R FILLER_98_957 ();
 DECAPx4_ASAP7_75t_R FILLER_98_979 ();
 FILLER_ASAP7_75t_R FILLER_98_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_991 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1157 ();
 FILLER_ASAP7_75t_R FILLER_98_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1212 ();
 FILLER_ASAP7_75t_R FILLER_98_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1244 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1276 ();
 FILLER_ASAP7_75t_R FILLER_98_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_99_2 ();
 FILLER_ASAP7_75t_R FILLER_99_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_18 ();
 DECAPx4_ASAP7_75t_R FILLER_99_25 ();
 DECAPx2_ASAP7_75t_R FILLER_99_41 ();
 FILLER_ASAP7_75t_R FILLER_99_47 ();
 DECAPx1_ASAP7_75t_R FILLER_99_67 ();
 DECAPx10_ASAP7_75t_R FILLER_99_77 ();
 DECAPx2_ASAP7_75t_R FILLER_99_99 ();
 FILLER_ASAP7_75t_R FILLER_99_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_115 ();
 FILLER_ASAP7_75t_R FILLER_99_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_131 ();
 DECAPx2_ASAP7_75t_R FILLER_99_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_145 ();
 DECAPx1_ASAP7_75t_R FILLER_99_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_156 ();
 DECAPx4_ASAP7_75t_R FILLER_99_173 ();
 DECAPx6_ASAP7_75t_R FILLER_99_201 ();
 DECAPx1_ASAP7_75t_R FILLER_99_215 ();
 FILLER_ASAP7_75t_R FILLER_99_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_263 ();
 FILLER_ASAP7_75t_R FILLER_99_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_273 ();
 DECAPx1_ASAP7_75t_R FILLER_99_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_298 ();
 DECAPx2_ASAP7_75t_R FILLER_99_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_330 ();
 DECAPx6_ASAP7_75t_R FILLER_99_339 ();
 DECAPx2_ASAP7_75t_R FILLER_99_353 ();
 DECAPx1_ASAP7_75t_R FILLER_99_377 ();
 DECAPx1_ASAP7_75t_R FILLER_99_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_395 ();
 DECAPx2_ASAP7_75t_R FILLER_99_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_409 ();
 FILLER_ASAP7_75t_R FILLER_99_431 ();
 FILLER_ASAP7_75t_R FILLER_99_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_464 ();
 FILLER_ASAP7_75t_R FILLER_99_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_517 ();
 DECAPx10_ASAP7_75t_R FILLER_99_528 ();
 DECAPx4_ASAP7_75t_R FILLER_99_550 ();
 FILLER_ASAP7_75t_R FILLER_99_566 ();
 DECAPx10_ASAP7_75t_R FILLER_99_575 ();
 DECAPx10_ASAP7_75t_R FILLER_99_597 ();
 DECAPx4_ASAP7_75t_R FILLER_99_619 ();
 FILLER_ASAP7_75t_R FILLER_99_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_631 ();
 DECAPx2_ASAP7_75t_R FILLER_99_662 ();
 DECAPx4_ASAP7_75t_R FILLER_99_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_688 ();
 DECAPx1_ASAP7_75t_R FILLER_99_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_699 ();
 FILLER_ASAP7_75t_R FILLER_99_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_726 ();
 DECAPx10_ASAP7_75t_R FILLER_99_742 ();
 DECAPx2_ASAP7_75t_R FILLER_99_764 ();
 FILLER_ASAP7_75t_R FILLER_99_770 ();
 DECAPx10_ASAP7_75t_R FILLER_99_778 ();
 DECAPx10_ASAP7_75t_R FILLER_99_800 ();
 DECAPx10_ASAP7_75t_R FILLER_99_822 ();
 DECAPx10_ASAP7_75t_R FILLER_99_844 ();
 DECAPx10_ASAP7_75t_R FILLER_99_866 ();
 DECAPx10_ASAP7_75t_R FILLER_99_888 ();
 DECAPx6_ASAP7_75t_R FILLER_99_910 ();
 DECAPx10_ASAP7_75t_R FILLER_99_926 ();
 DECAPx10_ASAP7_75t_R FILLER_99_948 ();
 DECAPx10_ASAP7_75t_R FILLER_99_970 ();
 DECAPx6_ASAP7_75t_R FILLER_99_992 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1040 ();
 FILLER_ASAP7_75t_R FILLER_99_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1110 ();
 FILLER_ASAP7_75t_R FILLER_99_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_99_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_99_1203 ();
 FILLER_ASAP7_75t_R FILLER_99_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1241 ();
 FILLER_ASAP7_75t_R FILLER_99_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1283 ();
 DECAPx4_ASAP7_75t_R FILLER_100_2 ();
 FILLER_ASAP7_75t_R FILLER_100_12 ();
 DECAPx1_ASAP7_75t_R FILLER_100_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_55 ();
 FILLER_ASAP7_75t_R FILLER_100_62 ();
 DECAPx1_ASAP7_75t_R FILLER_100_71 ();
 FILLER_ASAP7_75t_R FILLER_100_83 ();
 FILLER_ASAP7_75t_R FILLER_100_99 ();
 DECAPx2_ASAP7_75t_R FILLER_100_107 ();
 FILLER_ASAP7_75t_R FILLER_100_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_130 ();
 DECAPx1_ASAP7_75t_R FILLER_100_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_149 ();
 FILLER_ASAP7_75t_R FILLER_100_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_159 ();
 DECAPx4_ASAP7_75t_R FILLER_100_182 ();
 DECAPx6_ASAP7_75t_R FILLER_100_200 ();
 DECAPx1_ASAP7_75t_R FILLER_100_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_218 ();
 DECAPx4_ASAP7_75t_R FILLER_100_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_250 ();
 FILLER_ASAP7_75t_R FILLER_100_261 ();
 DECAPx2_ASAP7_75t_R FILLER_100_269 ();
 FILLER_ASAP7_75t_R FILLER_100_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_297 ();
 FILLER_ASAP7_75t_R FILLER_100_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_318 ();
 FILLER_ASAP7_75t_R FILLER_100_325 ();
 DECAPx10_ASAP7_75t_R FILLER_100_333 ();
 DECAPx10_ASAP7_75t_R FILLER_100_355 ();
 DECAPx4_ASAP7_75t_R FILLER_100_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_387 ();
 DECAPx6_ASAP7_75t_R FILLER_100_426 ();
 DECAPx1_ASAP7_75t_R FILLER_100_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_464 ();
 DECAPx6_ASAP7_75t_R FILLER_100_475 ();
 DECAPx1_ASAP7_75t_R FILLER_100_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_493 ();
 DECAPx6_ASAP7_75t_R FILLER_100_515 ();
 DECAPx10_ASAP7_75t_R FILLER_100_535 ();
 DECAPx6_ASAP7_75t_R FILLER_100_557 ();
 DECAPx1_ASAP7_75t_R FILLER_100_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_575 ();
 DECAPx10_ASAP7_75t_R FILLER_100_588 ();
 FILLER_ASAP7_75t_R FILLER_100_610 ();
 DECAPx10_ASAP7_75t_R FILLER_100_618 ();
 DECAPx10_ASAP7_75t_R FILLER_100_640 ();
 DECAPx2_ASAP7_75t_R FILLER_100_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_668 ();
 DECAPx4_ASAP7_75t_R FILLER_100_676 ();
 FILLER_ASAP7_75t_R FILLER_100_686 ();
 DECAPx1_ASAP7_75t_R FILLER_100_694 ();
 DECAPx10_ASAP7_75t_R FILLER_100_715 ();
 DECAPx10_ASAP7_75t_R FILLER_100_737 ();
 DECAPx10_ASAP7_75t_R FILLER_100_759 ();
 DECAPx10_ASAP7_75t_R FILLER_100_781 ();
 DECAPx10_ASAP7_75t_R FILLER_100_803 ();
 DECAPx6_ASAP7_75t_R FILLER_100_825 ();
 FILLER_ASAP7_75t_R FILLER_100_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_841 ();
 DECAPx10_ASAP7_75t_R FILLER_100_848 ();
 DECAPx6_ASAP7_75t_R FILLER_100_870 ();
 DECAPx2_ASAP7_75t_R FILLER_100_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_897 ();
 DECAPx4_ASAP7_75t_R FILLER_100_930 ();
 FILLER_ASAP7_75t_R FILLER_100_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_942 ();
 DECAPx10_ASAP7_75t_R FILLER_100_959 ();
 DECAPx10_ASAP7_75t_R FILLER_100_981 ();
 FILLER_ASAP7_75t_R FILLER_100_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1085 ();
 FILLER_ASAP7_75t_R FILLER_100_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1173 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1207 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_101_2 ();
 DECAPx6_ASAP7_75t_R FILLER_101_24 ();
 DECAPx1_ASAP7_75t_R FILLER_101_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_48 ();
 FILLER_ASAP7_75t_R FILLER_101_55 ();
 DECAPx2_ASAP7_75t_R FILLER_101_63 ();
 FILLER_ASAP7_75t_R FILLER_101_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_71 ();
 DECAPx4_ASAP7_75t_R FILLER_101_82 ();
 FILLER_ASAP7_75t_R FILLER_101_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_130 ();
 DECAPx2_ASAP7_75t_R FILLER_101_139 ();
 FILLER_ASAP7_75t_R FILLER_101_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_147 ();
 FILLER_ASAP7_75t_R FILLER_101_156 ();
 FILLER_ASAP7_75t_R FILLER_101_168 ();
 FILLER_ASAP7_75t_R FILLER_101_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_179 ();
 DECAPx1_ASAP7_75t_R FILLER_101_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_223 ();
 DECAPx6_ASAP7_75t_R FILLER_101_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_287 ();
 DECAPx4_ASAP7_75t_R FILLER_101_294 ();
 FILLER_ASAP7_75t_R FILLER_101_316 ();
 FILLER_ASAP7_75t_R FILLER_101_324 ();
 DECAPx2_ASAP7_75t_R FILLER_101_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_338 ();
 FILLER_ASAP7_75t_R FILLER_101_346 ();
 DECAPx6_ASAP7_75t_R FILLER_101_368 ();
 DECAPx2_ASAP7_75t_R FILLER_101_392 ();
 FILLER_ASAP7_75t_R FILLER_101_398 ();
 DECAPx6_ASAP7_75t_R FILLER_101_410 ();
 DECAPx2_ASAP7_75t_R FILLER_101_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_430 ();
 DECAPx6_ASAP7_75t_R FILLER_101_448 ();
 DECAPx4_ASAP7_75t_R FILLER_101_483 ();
 FILLER_ASAP7_75t_R FILLER_101_493 ();
 DECAPx4_ASAP7_75t_R FILLER_101_516 ();
 FILLER_ASAP7_75t_R FILLER_101_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_528 ();
 DECAPx10_ASAP7_75t_R FILLER_101_535 ();
 DECAPx1_ASAP7_75t_R FILLER_101_557 ();
 DECAPx10_ASAP7_75t_R FILLER_101_568 ();
 DECAPx10_ASAP7_75t_R FILLER_101_590 ();
 DECAPx6_ASAP7_75t_R FILLER_101_612 ();
 DECAPx2_ASAP7_75t_R FILLER_101_626 ();
 DECAPx4_ASAP7_75t_R FILLER_101_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_663 ();
 DECAPx10_ASAP7_75t_R FILLER_101_670 ();
 DECAPx10_ASAP7_75t_R FILLER_101_692 ();
 DECAPx2_ASAP7_75t_R FILLER_101_714 ();
 DECAPx10_ASAP7_75t_R FILLER_101_730 ();
 DECAPx10_ASAP7_75t_R FILLER_101_752 ();
 DECAPx1_ASAP7_75t_R FILLER_101_774 ();
 DECAPx10_ASAP7_75t_R FILLER_101_788 ();
 DECAPx4_ASAP7_75t_R FILLER_101_810 ();
 DECAPx4_ASAP7_75t_R FILLER_101_828 ();
 FILLER_ASAP7_75t_R FILLER_101_838 ();
 DECAPx4_ASAP7_75t_R FILLER_101_850 ();
 DECAPx10_ASAP7_75t_R FILLER_101_868 ();
 DECAPx10_ASAP7_75t_R FILLER_101_890 ();
 DECAPx4_ASAP7_75t_R FILLER_101_912 ();
 FILLER_ASAP7_75t_R FILLER_101_922 ();
 DECAPx10_ASAP7_75t_R FILLER_101_926 ();
 DECAPx10_ASAP7_75t_R FILLER_101_948 ();
 DECAPx1_ASAP7_75t_R FILLER_101_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_974 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1001 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1023 ();
 FILLER_ASAP7_75t_R FILLER_101_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1068 ();
 FILLER_ASAP7_75t_R FILLER_101_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1134 ();
 FILLER_ASAP7_75t_R FILLER_101_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1149 ();
 FILLER_ASAP7_75t_R FILLER_101_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1224 ();
 FILLER_ASAP7_75t_R FILLER_101_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1236 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_102_2 ();
 DECAPx1_ASAP7_75t_R FILLER_102_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_28 ();
 DECAPx1_ASAP7_75t_R FILLER_102_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_53 ();
 DECAPx10_ASAP7_75t_R FILLER_102_68 ();
 DECAPx1_ASAP7_75t_R FILLER_102_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_94 ();
 DECAPx4_ASAP7_75t_R FILLER_102_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_151 ();
 DECAPx2_ASAP7_75t_R FILLER_102_176 ();
 FILLER_ASAP7_75t_R FILLER_102_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_184 ();
 DECAPx6_ASAP7_75t_R FILLER_102_195 ();
 FILLER_ASAP7_75t_R FILLER_102_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_211 ();
 DECAPx6_ASAP7_75t_R FILLER_102_222 ();
 FILLER_ASAP7_75t_R FILLER_102_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_238 ();
 FILLER_ASAP7_75t_R FILLER_102_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_293 ();
 DECAPx4_ASAP7_75t_R FILLER_102_302 ();
 DECAPx1_ASAP7_75t_R FILLER_102_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_328 ();
 DECAPx1_ASAP7_75t_R FILLER_102_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_346 ();
 FILLER_ASAP7_75t_R FILLER_102_369 ();
 DECAPx4_ASAP7_75t_R FILLER_102_381 ();
 FILLER_ASAP7_75t_R FILLER_102_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_400 ();
 DECAPx1_ASAP7_75t_R FILLER_102_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_412 ();
 DECAPx1_ASAP7_75t_R FILLER_102_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_427 ();
 FILLER_ASAP7_75t_R FILLER_102_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_451 ();
 DECAPx1_ASAP7_75t_R FILLER_102_464 ();
 DECAPx2_ASAP7_75t_R FILLER_102_489 ();
 FILLER_ASAP7_75t_R FILLER_102_495 ();
 FILLER_ASAP7_75t_R FILLER_102_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_509 ();
 DECAPx2_ASAP7_75t_R FILLER_102_527 ();
 FILLER_ASAP7_75t_R FILLER_102_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_546 ();
 DECAPx10_ASAP7_75t_R FILLER_102_557 ();
 FILLER_ASAP7_75t_R FILLER_102_579 ();
 DECAPx10_ASAP7_75t_R FILLER_102_587 ();
 DECAPx2_ASAP7_75t_R FILLER_102_609 ();
 FILLER_ASAP7_75t_R FILLER_102_615 ();
 DECAPx1_ASAP7_75t_R FILLER_102_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_635 ();
 FILLER_ASAP7_75t_R FILLER_102_653 ();
 DECAPx10_ASAP7_75t_R FILLER_102_675 ();
 DECAPx4_ASAP7_75t_R FILLER_102_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_707 ();
 DECAPx2_ASAP7_75t_R FILLER_102_714 ();
 DECAPx2_ASAP7_75t_R FILLER_102_750 ();
 FILLER_ASAP7_75t_R FILLER_102_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_758 ();
 DECAPx10_ASAP7_75t_R FILLER_102_769 ();
 DECAPx10_ASAP7_75t_R FILLER_102_791 ();
 DECAPx10_ASAP7_75t_R FILLER_102_813 ();
 DECAPx10_ASAP7_75t_R FILLER_102_835 ();
 DECAPx10_ASAP7_75t_R FILLER_102_857 ();
 DECAPx10_ASAP7_75t_R FILLER_102_879 ();
 DECAPx10_ASAP7_75t_R FILLER_102_901 ();
 DECAPx10_ASAP7_75t_R FILLER_102_923 ();
 DECAPx10_ASAP7_75t_R FILLER_102_945 ();
 DECAPx10_ASAP7_75t_R FILLER_102_967 ();
 DECAPx10_ASAP7_75t_R FILLER_102_989 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1114 ();
 FILLER_ASAP7_75t_R FILLER_102_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1152 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_102_1245 ();
 FILLER_ASAP7_75t_R FILLER_102_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_103_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_19 ();
 DECAPx6_ASAP7_75t_R FILLER_103_45 ();
 DECAPx4_ASAP7_75t_R FILLER_103_65 ();
 FILLER_ASAP7_75t_R FILLER_103_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_77 ();
 DECAPx10_ASAP7_75t_R FILLER_103_84 ();
 DECAPx10_ASAP7_75t_R FILLER_103_106 ();
 FILLER_ASAP7_75t_R FILLER_103_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_130 ();
 DECAPx1_ASAP7_75t_R FILLER_103_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_151 ();
 DECAPx2_ASAP7_75t_R FILLER_103_160 ();
 FILLER_ASAP7_75t_R FILLER_103_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_168 ();
 DECAPx10_ASAP7_75t_R FILLER_103_193 ();
 DECAPx10_ASAP7_75t_R FILLER_103_215 ();
 DECAPx10_ASAP7_75t_R FILLER_103_237 ();
 DECAPx10_ASAP7_75t_R FILLER_103_259 ();
 DECAPx6_ASAP7_75t_R FILLER_103_281 ();
 FILLER_ASAP7_75t_R FILLER_103_295 ();
 DECAPx1_ASAP7_75t_R FILLER_103_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_329 ();
 FILLER_ASAP7_75t_R FILLER_103_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_367 ();
 DECAPx4_ASAP7_75t_R FILLER_103_376 ();
 FILLER_ASAP7_75t_R FILLER_103_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_410 ();
 FILLER_ASAP7_75t_R FILLER_103_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_420 ();
 DECAPx4_ASAP7_75t_R FILLER_103_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_469 ();
 DECAPx10_ASAP7_75t_R FILLER_103_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_509 ();
 DECAPx2_ASAP7_75t_R FILLER_103_531 ();
 DECAPx10_ASAP7_75t_R FILLER_103_544 ();
 DECAPx4_ASAP7_75t_R FILLER_103_566 ();
 DECAPx6_ASAP7_75t_R FILLER_103_600 ();
 DECAPx1_ASAP7_75t_R FILLER_103_614 ();
 DECAPx4_ASAP7_75t_R FILLER_103_627 ();
 FILLER_ASAP7_75t_R FILLER_103_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_639 ();
 DECAPx6_ASAP7_75t_R FILLER_103_678 ();
 DECAPx1_ASAP7_75t_R FILLER_103_692 ();
 FILLER_ASAP7_75t_R FILLER_103_716 ();
 FILLER_ASAP7_75t_R FILLER_103_728 ();
 DECAPx6_ASAP7_75t_R FILLER_103_736 ();
 DECAPx2_ASAP7_75t_R FILLER_103_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_756 ();
 DECAPx10_ASAP7_75t_R FILLER_103_769 ();
 DECAPx10_ASAP7_75t_R FILLER_103_791 ();
 DECAPx10_ASAP7_75t_R FILLER_103_813 ();
 DECAPx10_ASAP7_75t_R FILLER_103_835 ();
 DECAPx10_ASAP7_75t_R FILLER_103_857 ();
 DECAPx10_ASAP7_75t_R FILLER_103_879 ();
 DECAPx10_ASAP7_75t_R FILLER_103_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_923 ();
 DECAPx1_ASAP7_75t_R FILLER_103_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_930 ();
 DECAPx10_ASAP7_75t_R FILLER_103_937 ();
 DECAPx10_ASAP7_75t_R FILLER_103_959 ();
 DECAPx10_ASAP7_75t_R FILLER_103_981 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1066 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_103_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1186 ();
 FILLER_ASAP7_75t_R FILLER_103_1221 ();
 FILLER_ASAP7_75t_R FILLER_103_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1247 ();
 FILLER_ASAP7_75t_R FILLER_103_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_104_2 ();
 FILLER_ASAP7_75t_R FILLER_104_16 ();
 DECAPx6_ASAP7_75t_R FILLER_104_24 ();
 FILLER_ASAP7_75t_R FILLER_104_38 ();
 DECAPx2_ASAP7_75t_R FILLER_104_50 ();
 FILLER_ASAP7_75t_R FILLER_104_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_58 ();
 FILLER_ASAP7_75t_R FILLER_104_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_68 ();
 DECAPx1_ASAP7_75t_R FILLER_104_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_81 ();
 DECAPx2_ASAP7_75t_R FILLER_104_90 ();
 FILLER_ASAP7_75t_R FILLER_104_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_98 ();
 DECAPx2_ASAP7_75t_R FILLER_104_106 ();
 FILLER_ASAP7_75t_R FILLER_104_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_114 ();
 DECAPx2_ASAP7_75t_R FILLER_104_123 ();
 DECAPx1_ASAP7_75t_R FILLER_104_137 ();
 DECAPx10_ASAP7_75t_R FILLER_104_148 ();
 FILLER_ASAP7_75t_R FILLER_104_170 ();
 DECAPx4_ASAP7_75t_R FILLER_104_208 ();
 FILLER_ASAP7_75t_R FILLER_104_218 ();
 DECAPx10_ASAP7_75t_R FILLER_104_230 ();
 DECAPx10_ASAP7_75t_R FILLER_104_252 ();
 DECAPx4_ASAP7_75t_R FILLER_104_274 ();
 FILLER_ASAP7_75t_R FILLER_104_284 ();
 DECAPx6_ASAP7_75t_R FILLER_104_293 ();
 FILLER_ASAP7_75t_R FILLER_104_307 ();
 FILLER_ASAP7_75t_R FILLER_104_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_317 ();
 DECAPx2_ASAP7_75t_R FILLER_104_332 ();
 FILLER_ASAP7_75t_R FILLER_104_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_340 ();
 FILLER_ASAP7_75t_R FILLER_104_347 ();
 FILLER_ASAP7_75t_R FILLER_104_361 ();
 DECAPx6_ASAP7_75t_R FILLER_104_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_385 ();
 DECAPx1_ASAP7_75t_R FILLER_104_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_440 ();
 FILLER_ASAP7_75t_R FILLER_104_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_483 ();
 DECAPx6_ASAP7_75t_R FILLER_104_494 ();
 FILLER_ASAP7_75t_R FILLER_104_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_517 ();
 DECAPx2_ASAP7_75t_R FILLER_104_528 ();
 FILLER_ASAP7_75t_R FILLER_104_534 ();
 DECAPx4_ASAP7_75t_R FILLER_104_557 ();
 FILLER_ASAP7_75t_R FILLER_104_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_569 ();
 DECAPx6_ASAP7_75t_R FILLER_104_580 ();
 DECAPx2_ASAP7_75t_R FILLER_104_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_621 ();
 DECAPx6_ASAP7_75t_R FILLER_104_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_680 ();
 DECAPx1_ASAP7_75t_R FILLER_104_698 ();
 DECAPx10_ASAP7_75t_R FILLER_104_735 ();
 FILLER_ASAP7_75t_R FILLER_104_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_759 ();
 DECAPx1_ASAP7_75t_R FILLER_104_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_774 ();
 DECAPx10_ASAP7_75t_R FILLER_104_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_807 ();
 DECAPx10_ASAP7_75t_R FILLER_104_814 ();
 DECAPx10_ASAP7_75t_R FILLER_104_836 ();
 DECAPx10_ASAP7_75t_R FILLER_104_858 ();
 DECAPx10_ASAP7_75t_R FILLER_104_880 ();
 DECAPx10_ASAP7_75t_R FILLER_104_902 ();
 DECAPx10_ASAP7_75t_R FILLER_104_924 ();
 DECAPx6_ASAP7_75t_R FILLER_104_946 ();
 FILLER_ASAP7_75t_R FILLER_104_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_962 ();
 DECAPx1_ASAP7_75t_R FILLER_104_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_973 ();
 DECAPx2_ASAP7_75t_R FILLER_104_982 ();
 DECAPx4_ASAP7_75t_R FILLER_104_998 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1014 ();
 FILLER_ASAP7_75t_R FILLER_104_1030 ();
 FILLER_ASAP7_75t_R FILLER_104_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1093 ();
 FILLER_ASAP7_75t_R FILLER_104_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1182 ();
 FILLER_ASAP7_75t_R FILLER_104_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1197 ();
 FILLER_ASAP7_75t_R FILLER_104_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1212 ();
 FILLER_ASAP7_75t_R FILLER_104_1223 ();
 FILLER_ASAP7_75t_R FILLER_104_1270 ();
 DECAPx4_ASAP7_75t_R FILLER_105_2 ();
 FILLER_ASAP7_75t_R FILLER_105_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_14 ();
 DECAPx1_ASAP7_75t_R FILLER_105_27 ();
 DECAPx1_ASAP7_75t_R FILLER_105_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_68 ();
 FILLER_ASAP7_75t_R FILLER_105_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_89 ();
 DECAPx4_ASAP7_75t_R FILLER_105_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_107 ();
 DECAPx10_ASAP7_75t_R FILLER_105_128 ();
 DECAPx1_ASAP7_75t_R FILLER_105_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_154 ();
 DECAPx1_ASAP7_75t_R FILLER_105_169 ();
 DECAPx10_ASAP7_75t_R FILLER_105_210 ();
 DECAPx10_ASAP7_75t_R FILLER_105_232 ();
 DECAPx10_ASAP7_75t_R FILLER_105_254 ();
 DECAPx6_ASAP7_75t_R FILLER_105_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_290 ();
 DECAPx6_ASAP7_75t_R FILLER_105_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_338 ();
 FILLER_ASAP7_75t_R FILLER_105_345 ();
 DECAPx2_ASAP7_75t_R FILLER_105_353 ();
 FILLER_ASAP7_75t_R FILLER_105_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_361 ();
 DECAPx6_ASAP7_75t_R FILLER_105_384 ();
 DECAPx1_ASAP7_75t_R FILLER_105_398 ();
 DECAPx10_ASAP7_75t_R FILLER_105_412 ();
 FILLER_ASAP7_75t_R FILLER_105_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_436 ();
 DECAPx2_ASAP7_75t_R FILLER_105_468 ();
 FILLER_ASAP7_75t_R FILLER_105_495 ();
 DECAPx1_ASAP7_75t_R FILLER_105_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_518 ();
 DECAPx6_ASAP7_75t_R FILLER_105_529 ();
 DECAPx6_ASAP7_75t_R FILLER_105_553 ();
 FILLER_ASAP7_75t_R FILLER_105_567 ();
 DECAPx2_ASAP7_75t_R FILLER_105_581 ();
 FILLER_ASAP7_75t_R FILLER_105_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_589 ();
 DECAPx2_ASAP7_75t_R FILLER_105_597 ();
 FILLER_ASAP7_75t_R FILLER_105_603 ();
 FILLER_ASAP7_75t_R FILLER_105_612 ();
 FILLER_ASAP7_75t_R FILLER_105_624 ();
 DECAPx6_ASAP7_75t_R FILLER_105_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_646 ();
 FILLER_ASAP7_75t_R FILLER_105_657 ();
 DECAPx2_ASAP7_75t_R FILLER_105_676 ();
 FILLER_ASAP7_75t_R FILLER_105_710 ();
 DECAPx2_ASAP7_75t_R FILLER_105_718 ();
 DECAPx10_ASAP7_75t_R FILLER_105_738 ();
 DECAPx10_ASAP7_75t_R FILLER_105_760 ();
 DECAPx10_ASAP7_75t_R FILLER_105_782 ();
 DECAPx1_ASAP7_75t_R FILLER_105_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_808 ();
 FILLER_ASAP7_75t_R FILLER_105_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_817 ();
 DECAPx6_ASAP7_75t_R FILLER_105_828 ();
 DECAPx2_ASAP7_75t_R FILLER_105_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_848 ();
 DECAPx10_ASAP7_75t_R FILLER_105_855 ();
 FILLER_ASAP7_75t_R FILLER_105_877 ();
 DECAPx10_ASAP7_75t_R FILLER_105_898 ();
 DECAPx1_ASAP7_75t_R FILLER_105_920 ();
 DECAPx6_ASAP7_75t_R FILLER_105_926 ();
 FILLER_ASAP7_75t_R FILLER_105_940 ();
 DECAPx10_ASAP7_75t_R FILLER_105_950 ();
 DECAPx10_ASAP7_75t_R FILLER_105_972 ();
 DECAPx10_ASAP7_75t_R FILLER_105_994 ();
 FILLER_ASAP7_75t_R FILLER_105_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1068 ();
 FILLER_ASAP7_75t_R FILLER_105_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1099 ();
 FILLER_ASAP7_75t_R FILLER_105_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1107 ();
 FILLER_ASAP7_75t_R FILLER_105_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1135 ();
 FILLER_ASAP7_75t_R FILLER_105_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1150 ();
 FILLER_ASAP7_75t_R FILLER_105_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_105_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_105_1218 ();
 FILLER_ASAP7_75t_R FILLER_105_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1234 ();
 FILLER_ASAP7_75t_R FILLER_105_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1285 ();
 FILLER_ASAP7_75t_R FILLER_105_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_106_2 ();
 DECAPx2_ASAP7_75t_R FILLER_106_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_22 ();
 DECAPx2_ASAP7_75t_R FILLER_106_29 ();
 FILLER_ASAP7_75t_R FILLER_106_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_44 ();
 DECAPx1_ASAP7_75t_R FILLER_106_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_66 ();
 DECAPx6_ASAP7_75t_R FILLER_106_80 ();
 DECAPx4_ASAP7_75t_R FILLER_106_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_118 ();
 DECAPx4_ASAP7_75t_R FILLER_106_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_136 ();
 FILLER_ASAP7_75t_R FILLER_106_151 ();
 DECAPx1_ASAP7_75t_R FILLER_106_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_178 ();
 DECAPx10_ASAP7_75t_R FILLER_106_186 ();
 DECAPx10_ASAP7_75t_R FILLER_106_208 ();
 DECAPx6_ASAP7_75t_R FILLER_106_230 ();
 DECAPx4_ASAP7_75t_R FILLER_106_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_264 ();
 FILLER_ASAP7_75t_R FILLER_106_275 ();
 DECAPx6_ASAP7_75t_R FILLER_106_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_297 ();
 DECAPx6_ASAP7_75t_R FILLER_106_305 ();
 DECAPx1_ASAP7_75t_R FILLER_106_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_323 ();
 DECAPx4_ASAP7_75t_R FILLER_106_330 ();
 DECAPx10_ASAP7_75t_R FILLER_106_354 ();
 DECAPx6_ASAP7_75t_R FILLER_106_376 ();
 DECAPx2_ASAP7_75t_R FILLER_106_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_396 ();
 DECAPx2_ASAP7_75t_R FILLER_106_407 ();
 FILLER_ASAP7_75t_R FILLER_106_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_415 ();
 DECAPx2_ASAP7_75t_R FILLER_106_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_432 ();
 DECAPx2_ASAP7_75t_R FILLER_106_445 ();
 FILLER_ASAP7_75t_R FILLER_106_451 ();
 FILLER_ASAP7_75t_R FILLER_106_460 ();
 DECAPx2_ASAP7_75t_R FILLER_106_464 ();
 FILLER_ASAP7_75t_R FILLER_106_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_472 ();
 DECAPx1_ASAP7_75t_R FILLER_106_491 ();
 DECAPx6_ASAP7_75t_R FILLER_106_516 ();
 FILLER_ASAP7_75t_R FILLER_106_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_532 ();
 FILLER_ASAP7_75t_R FILLER_106_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_556 ();
 DECAPx1_ASAP7_75t_R FILLER_106_564 ();
 DECAPx6_ASAP7_75t_R FILLER_106_578 ();
 DECAPx2_ASAP7_75t_R FILLER_106_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_598 ();
 FILLER_ASAP7_75t_R FILLER_106_613 ();
 DECAPx2_ASAP7_75t_R FILLER_106_621 ();
 DECAPx4_ASAP7_75t_R FILLER_106_633 ();
 FILLER_ASAP7_75t_R FILLER_106_643 ();
 DECAPx4_ASAP7_75t_R FILLER_106_652 ();
 FILLER_ASAP7_75t_R FILLER_106_689 ();
 DECAPx1_ASAP7_75t_R FILLER_106_701 ();
 DECAPx10_ASAP7_75t_R FILLER_106_715 ();
 DECAPx10_ASAP7_75t_R FILLER_106_737 ();
 DECAPx10_ASAP7_75t_R FILLER_106_759 ();
 DECAPx10_ASAP7_75t_R FILLER_106_781 ();
 DECAPx10_ASAP7_75t_R FILLER_106_803 ();
 DECAPx10_ASAP7_75t_R FILLER_106_825 ();
 DECAPx10_ASAP7_75t_R FILLER_106_847 ();
 DECAPx10_ASAP7_75t_R FILLER_106_869 ();
 DECAPx2_ASAP7_75t_R FILLER_106_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_897 ();
 DECAPx4_ASAP7_75t_R FILLER_106_908 ();
 DECAPx10_ASAP7_75t_R FILLER_106_928 ();
 DECAPx10_ASAP7_75t_R FILLER_106_950 ();
 DECAPx6_ASAP7_75t_R FILLER_106_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_986 ();
 DECAPx10_ASAP7_75t_R FILLER_106_993 ();
 FILLER_ASAP7_75t_R FILLER_106_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1023 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1071 ();
 FILLER_ASAP7_75t_R FILLER_106_1081 ();
 FILLER_ASAP7_75t_R FILLER_106_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1163 ();
 FILLER_ASAP7_75t_R FILLER_106_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1197 ();
 FILLER_ASAP7_75t_R FILLER_106_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1234 ();
 FILLER_ASAP7_75t_R FILLER_106_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_107_2 ();
 DECAPx4_ASAP7_75t_R FILLER_107_24 ();
 FILLER_ASAP7_75t_R FILLER_107_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_36 ();
 DECAPx2_ASAP7_75t_R FILLER_107_45 ();
 FILLER_ASAP7_75t_R FILLER_107_51 ();
 DECAPx4_ASAP7_75t_R FILLER_107_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_70 ();
 DECAPx4_ASAP7_75t_R FILLER_107_77 ();
 FILLER_ASAP7_75t_R FILLER_107_87 ();
 FILLER_ASAP7_75t_R FILLER_107_113 ();
 FILLER_ASAP7_75t_R FILLER_107_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_141 ();
 FILLER_ASAP7_75t_R FILLER_107_158 ();
 FILLER_ASAP7_75t_R FILLER_107_166 ();
 FILLER_ASAP7_75t_R FILLER_107_174 ();
 DECAPx6_ASAP7_75t_R FILLER_107_200 ();
 DECAPx1_ASAP7_75t_R FILLER_107_214 ();
 DECAPx6_ASAP7_75t_R FILLER_107_228 ();
 DECAPx1_ASAP7_75t_R FILLER_107_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_246 ();
 DECAPx10_ASAP7_75t_R FILLER_107_257 ();
 DECAPx1_ASAP7_75t_R FILLER_107_279 ();
 FILLER_ASAP7_75t_R FILLER_107_293 ();
 DECAPx10_ASAP7_75t_R FILLER_107_302 ();
 DECAPx6_ASAP7_75t_R FILLER_107_324 ();
 FILLER_ASAP7_75t_R FILLER_107_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_340 ();
 DECAPx10_ASAP7_75t_R FILLER_107_370 ();
 DECAPx10_ASAP7_75t_R FILLER_107_392 ();
 DECAPx2_ASAP7_75t_R FILLER_107_421 ();
 DECAPx10_ASAP7_75t_R FILLER_107_449 ();
 DECAPx4_ASAP7_75t_R FILLER_107_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_481 ();
 DECAPx1_ASAP7_75t_R FILLER_107_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_507 ();
 DECAPx2_ASAP7_75t_R FILLER_107_515 ();
 FILLER_ASAP7_75t_R FILLER_107_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_523 ();
 DECAPx2_ASAP7_75t_R FILLER_107_534 ();
 FILLER_ASAP7_75t_R FILLER_107_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_542 ();
 DECAPx2_ASAP7_75t_R FILLER_107_550 ();
 DECAPx2_ASAP7_75t_R FILLER_107_587 ();
 FILLER_ASAP7_75t_R FILLER_107_593 ();
 DECAPx1_ASAP7_75t_R FILLER_107_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_615 ();
 DECAPx10_ASAP7_75t_R FILLER_107_622 ();
 FILLER_ASAP7_75t_R FILLER_107_644 ();
 DECAPx4_ASAP7_75t_R FILLER_107_667 ();
 FILLER_ASAP7_75t_R FILLER_107_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_715 ();
 DECAPx10_ASAP7_75t_R FILLER_107_737 ();
 DECAPx10_ASAP7_75t_R FILLER_107_759 ();
 DECAPx10_ASAP7_75t_R FILLER_107_781 ();
 DECAPx1_ASAP7_75t_R FILLER_107_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_807 ();
 DECAPx10_ASAP7_75t_R FILLER_107_822 ();
 DECAPx10_ASAP7_75t_R FILLER_107_844 ();
 DECAPx2_ASAP7_75t_R FILLER_107_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_872 ();
 DECAPx10_ASAP7_75t_R FILLER_107_880 ();
 DECAPx10_ASAP7_75t_R FILLER_107_902 ();
 DECAPx6_ASAP7_75t_R FILLER_107_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_940 ();
 DECAPx10_ASAP7_75t_R FILLER_107_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_971 ();
 DECAPx2_ASAP7_75t_R FILLER_107_982 ();
 FILLER_ASAP7_75t_R FILLER_107_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_990 ();
 DECAPx10_ASAP7_75t_R FILLER_107_999 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1021 ();
 FILLER_ASAP7_75t_R FILLER_107_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1097 ();
 FILLER_ASAP7_75t_R FILLER_107_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_107_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1184 ();
 FILLER_ASAP7_75t_R FILLER_107_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1233 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_108_2 ();
 DECAPx2_ASAP7_75t_R FILLER_108_24 ();
 FILLER_ASAP7_75t_R FILLER_108_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_32 ();
 DECAPx6_ASAP7_75t_R FILLER_108_54 ();
 DECAPx1_ASAP7_75t_R FILLER_108_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_72 ();
 DECAPx2_ASAP7_75t_R FILLER_108_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_103 ();
 DECAPx6_ASAP7_75t_R FILLER_108_129 ();
 DECAPx2_ASAP7_75t_R FILLER_108_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_156 ();
 DECAPx4_ASAP7_75t_R FILLER_108_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_175 ();
 DECAPx10_ASAP7_75t_R FILLER_108_194 ();
 FILLER_ASAP7_75t_R FILLER_108_216 ();
 DECAPx2_ASAP7_75t_R FILLER_108_221 ();
 FILLER_ASAP7_75t_R FILLER_108_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_229 ();
 DECAPx6_ASAP7_75t_R FILLER_108_256 ();
 FILLER_ASAP7_75t_R FILLER_108_270 ();
 FILLER_ASAP7_75t_R FILLER_108_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_280 ();
 DECAPx10_ASAP7_75t_R FILLER_108_291 ();
 DECAPx1_ASAP7_75t_R FILLER_108_313 ();
 DECAPx10_ASAP7_75t_R FILLER_108_324 ();
 DECAPx10_ASAP7_75t_R FILLER_108_346 ();
 DECAPx10_ASAP7_75t_R FILLER_108_368 ();
 DECAPx2_ASAP7_75t_R FILLER_108_390 ();
 FILLER_ASAP7_75t_R FILLER_108_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_405 ();
 FILLER_ASAP7_75t_R FILLER_108_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_439 ();
 DECAPx1_ASAP7_75t_R FILLER_108_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_454 ();
 DECAPx6_ASAP7_75t_R FILLER_108_464 ();
 FILLER_ASAP7_75t_R FILLER_108_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_480 ();
 DECAPx2_ASAP7_75t_R FILLER_108_498 ();
 FILLER_ASAP7_75t_R FILLER_108_504 ();
 DECAPx4_ASAP7_75t_R FILLER_108_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_558 ();
 DECAPx1_ASAP7_75t_R FILLER_108_611 ();
 DECAPx4_ASAP7_75t_R FILLER_108_625 ();
 DECAPx10_ASAP7_75t_R FILLER_108_655 ();
 DECAPx10_ASAP7_75t_R FILLER_108_677 ();
 DECAPx10_ASAP7_75t_R FILLER_108_699 ();
 DECAPx10_ASAP7_75t_R FILLER_108_721 ();
 DECAPx10_ASAP7_75t_R FILLER_108_757 ();
 DECAPx10_ASAP7_75t_R FILLER_108_779 ();
 DECAPx10_ASAP7_75t_R FILLER_108_801 ();
 DECAPx10_ASAP7_75t_R FILLER_108_823 ();
 DECAPx10_ASAP7_75t_R FILLER_108_845 ();
 DECAPx6_ASAP7_75t_R FILLER_108_867 ();
 DECAPx2_ASAP7_75t_R FILLER_108_881 ();
 DECAPx10_ASAP7_75t_R FILLER_108_893 ();
 DECAPx10_ASAP7_75t_R FILLER_108_915 ();
 DECAPx6_ASAP7_75t_R FILLER_108_937 ();
 DECAPx2_ASAP7_75t_R FILLER_108_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_957 ();
 DECAPx10_ASAP7_75t_R FILLER_108_968 ();
 DECAPx4_ASAP7_75t_R FILLER_108_990 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1020 ();
 FILLER_ASAP7_75t_R FILLER_108_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1110 ();
 FILLER_ASAP7_75t_R FILLER_108_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1137 ();
 FILLER_ASAP7_75t_R FILLER_108_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_109_2 ();
 FILLER_ASAP7_75t_R FILLER_109_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_62 ();
 DECAPx1_ASAP7_75t_R FILLER_109_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_95 ();
 FILLER_ASAP7_75t_R FILLER_109_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_117 ();
 DECAPx2_ASAP7_75t_R FILLER_109_125 ();
 FILLER_ASAP7_75t_R FILLER_109_131 ();
 FILLER_ASAP7_75t_R FILLER_109_146 ();
 DECAPx1_ASAP7_75t_R FILLER_109_156 ();
 FILLER_ASAP7_75t_R FILLER_109_168 ();
 DECAPx10_ASAP7_75t_R FILLER_109_190 ();
 DECAPx4_ASAP7_75t_R FILLER_109_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_222 ();
 DECAPx4_ASAP7_75t_R FILLER_109_233 ();
 FILLER_ASAP7_75t_R FILLER_109_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_252 ();
 DECAPx2_ASAP7_75t_R FILLER_109_259 ();
 DECAPx2_ASAP7_75t_R FILLER_109_275 ();
 DECAPx4_ASAP7_75t_R FILLER_109_293 ();
 DECAPx10_ASAP7_75t_R FILLER_109_310 ();
 DECAPx6_ASAP7_75t_R FILLER_109_332 ();
 DECAPx1_ASAP7_75t_R FILLER_109_346 ();
 DECAPx10_ASAP7_75t_R FILLER_109_355 ();
 DECAPx10_ASAP7_75t_R FILLER_109_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_399 ();
 DECAPx4_ASAP7_75t_R FILLER_109_421 ();
 DECAPx1_ASAP7_75t_R FILLER_109_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_452 ();
 FILLER_ASAP7_75t_R FILLER_109_474 ();
 DECAPx1_ASAP7_75t_R FILLER_109_497 ();
 DECAPx1_ASAP7_75t_R FILLER_109_518 ();
 DECAPx6_ASAP7_75t_R FILLER_109_536 ();
 FILLER_ASAP7_75t_R FILLER_109_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_581 ();
 DECAPx4_ASAP7_75t_R FILLER_109_599 ();
 DECAPx6_ASAP7_75t_R FILLER_109_643 ();
 DECAPx1_ASAP7_75t_R FILLER_109_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_674 ();
 DECAPx10_ASAP7_75t_R FILLER_109_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_703 ();
 FILLER_ASAP7_75t_R FILLER_109_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_720 ();
 DECAPx6_ASAP7_75t_R FILLER_109_729 ();
 DECAPx4_ASAP7_75t_R FILLER_109_749 ();
 DECAPx10_ASAP7_75t_R FILLER_109_769 ();
 DECAPx10_ASAP7_75t_R FILLER_109_791 ();
 DECAPx10_ASAP7_75t_R FILLER_109_813 ();
 DECAPx4_ASAP7_75t_R FILLER_109_835 ();
 DECAPx6_ASAP7_75t_R FILLER_109_853 ();
 FILLER_ASAP7_75t_R FILLER_109_867 ();
 FILLER_ASAP7_75t_R FILLER_109_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_888 ();
 DECAPx6_ASAP7_75t_R FILLER_109_895 ();
 DECAPx2_ASAP7_75t_R FILLER_109_909 ();
 FILLER_ASAP7_75t_R FILLER_109_926 ();
 FILLER_ASAP7_75t_R FILLER_109_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_940 ();
 FILLER_ASAP7_75t_R FILLER_109_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_951 ();
 FILLER_ASAP7_75t_R FILLER_109_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_960 ();
 DECAPx2_ASAP7_75t_R FILLER_109_970 ();
 DECAPx10_ASAP7_75t_R FILLER_109_993 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1015 ();
 FILLER_ASAP7_75t_R FILLER_109_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1078 ();
 FILLER_ASAP7_75t_R FILLER_109_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1135 ();
 FILLER_ASAP7_75t_R FILLER_109_1141 ();
 FILLER_ASAP7_75t_R FILLER_109_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1205 ();
 FILLER_ASAP7_75t_R FILLER_109_1215 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1249 ();
 FILLER_ASAP7_75t_R FILLER_109_1255 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1285 ();
 FILLER_ASAP7_75t_R FILLER_109_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_110_2 ();
 DECAPx2_ASAP7_75t_R FILLER_110_24 ();
 FILLER_ASAP7_75t_R FILLER_110_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_32 ();
 DECAPx2_ASAP7_75t_R FILLER_110_53 ();
 FILLER_ASAP7_75t_R FILLER_110_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_79 ();
 DECAPx2_ASAP7_75t_R FILLER_110_86 ();
 FILLER_ASAP7_75t_R FILLER_110_92 ();
 DECAPx2_ASAP7_75t_R FILLER_110_106 ();
 FILLER_ASAP7_75t_R FILLER_110_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_136 ();
 FILLER_ASAP7_75t_R FILLER_110_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_146 ();
 DECAPx2_ASAP7_75t_R FILLER_110_169 ();
 FILLER_ASAP7_75t_R FILLER_110_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_187 ();
 DECAPx10_ASAP7_75t_R FILLER_110_191 ();
 DECAPx2_ASAP7_75t_R FILLER_110_213 ();
 FILLER_ASAP7_75t_R FILLER_110_219 ();
 DECAPx2_ASAP7_75t_R FILLER_110_241 ();
 DECAPx2_ASAP7_75t_R FILLER_110_257 ();
 FILLER_ASAP7_75t_R FILLER_110_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_265 ();
 DECAPx1_ASAP7_75t_R FILLER_110_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_296 ();
 DECAPx2_ASAP7_75t_R FILLER_110_311 ();
 FILLER_ASAP7_75t_R FILLER_110_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_319 ();
 DECAPx1_ASAP7_75t_R FILLER_110_330 ();
 FILLER_ASAP7_75t_R FILLER_110_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_350 ();
 DECAPx10_ASAP7_75t_R FILLER_110_361 ();
 DECAPx4_ASAP7_75t_R FILLER_110_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_393 ();
 DECAPx4_ASAP7_75t_R FILLER_110_418 ();
 FILLER_ASAP7_75t_R FILLER_110_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_430 ();
 FILLER_ASAP7_75t_R FILLER_110_474 ();
 DECAPx1_ASAP7_75t_R FILLER_110_483 ();
 DECAPx1_ASAP7_75t_R FILLER_110_541 ();
 DECAPx10_ASAP7_75t_R FILLER_110_568 ();
 DECAPx6_ASAP7_75t_R FILLER_110_590 ();
 FILLER_ASAP7_75t_R FILLER_110_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_606 ();
 DECAPx4_ASAP7_75t_R FILLER_110_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_634 ();
 DECAPx10_ASAP7_75t_R FILLER_110_641 ();
 DECAPx10_ASAP7_75t_R FILLER_110_663 ();
 DECAPx10_ASAP7_75t_R FILLER_110_685 ();
 DECAPx10_ASAP7_75t_R FILLER_110_707 ();
 DECAPx10_ASAP7_75t_R FILLER_110_729 ();
 DECAPx10_ASAP7_75t_R FILLER_110_751 ();
 DECAPx10_ASAP7_75t_R FILLER_110_773 ();
 DECAPx2_ASAP7_75t_R FILLER_110_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_801 ();
 FILLER_ASAP7_75t_R FILLER_110_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_810 ();
 DECAPx1_ASAP7_75t_R FILLER_110_823 ();
 DECAPx10_ASAP7_75t_R FILLER_110_837 ();
 DECAPx1_ASAP7_75t_R FILLER_110_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_863 ();
 DECAPx10_ASAP7_75t_R FILLER_110_885 ();
 DECAPx6_ASAP7_75t_R FILLER_110_907 ();
 FILLER_ASAP7_75t_R FILLER_110_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_923 ();
 DECAPx10_ASAP7_75t_R FILLER_110_930 ();
 DECAPx10_ASAP7_75t_R FILLER_110_952 ();
 DECAPx6_ASAP7_75t_R FILLER_110_974 ();
 DECAPx1_ASAP7_75t_R FILLER_110_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_992 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1053 ();
 FILLER_ASAP7_75t_R FILLER_110_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1061 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1068 ();
 FILLER_ASAP7_75t_R FILLER_110_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1090 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1097 ();
 FILLER_ASAP7_75t_R FILLER_110_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1178 ();
 FILLER_ASAP7_75t_R FILLER_110_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_111_2 ();
 FILLER_ASAP7_75t_R FILLER_111_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_43 ();
 DECAPx10_ASAP7_75t_R FILLER_111_51 ();
 DECAPx6_ASAP7_75t_R FILLER_111_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_87 ();
 DECAPx2_ASAP7_75t_R FILLER_111_114 ();
 FILLER_ASAP7_75t_R FILLER_111_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_135 ();
 DECAPx6_ASAP7_75t_R FILLER_111_143 ();
 DECAPx10_ASAP7_75t_R FILLER_111_181 ();
 DECAPx4_ASAP7_75t_R FILLER_111_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_213 ();
 DECAPx10_ASAP7_75t_R FILLER_111_224 ();
 DECAPx1_ASAP7_75t_R FILLER_111_246 ();
 DECAPx4_ASAP7_75t_R FILLER_111_266 ();
 DECAPx4_ASAP7_75t_R FILLER_111_292 ();
 FILLER_ASAP7_75t_R FILLER_111_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_304 ();
 DECAPx6_ASAP7_75t_R FILLER_111_328 ();
 FILLER_ASAP7_75t_R FILLER_111_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_344 ();
 DECAPx4_ASAP7_75t_R FILLER_111_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_369 ();
 DECAPx10_ASAP7_75t_R FILLER_111_396 ();
 DECAPx6_ASAP7_75t_R FILLER_111_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_432 ();
 DECAPx2_ASAP7_75t_R FILLER_111_449 ();
 FILLER_ASAP7_75t_R FILLER_111_455 ();
 DECAPx1_ASAP7_75t_R FILLER_111_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_482 ();
 DECAPx2_ASAP7_75t_R FILLER_111_493 ();
 FILLER_ASAP7_75t_R FILLER_111_499 ();
 FILLER_ASAP7_75t_R FILLER_111_552 ();
 DECAPx10_ASAP7_75t_R FILLER_111_566 ();
 DECAPx6_ASAP7_75t_R FILLER_111_588 ();
 DECAPx10_ASAP7_75t_R FILLER_111_633 ();
 DECAPx10_ASAP7_75t_R FILLER_111_655 ();
 DECAPx6_ASAP7_75t_R FILLER_111_677 ();
 FILLER_ASAP7_75t_R FILLER_111_691 ();
 FILLER_ASAP7_75t_R FILLER_111_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_716 ();
 DECAPx2_ASAP7_75t_R FILLER_111_724 ();
 FILLER_ASAP7_75t_R FILLER_111_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_732 ();
 DECAPx10_ASAP7_75t_R FILLER_111_741 ();
 DECAPx10_ASAP7_75t_R FILLER_111_763 ();
 DECAPx10_ASAP7_75t_R FILLER_111_785 ();
 DECAPx4_ASAP7_75t_R FILLER_111_807 ();
 DECAPx10_ASAP7_75t_R FILLER_111_823 ();
 DECAPx10_ASAP7_75t_R FILLER_111_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_867 ();
 FILLER_ASAP7_75t_R FILLER_111_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_884 ();
 DECAPx4_ASAP7_75t_R FILLER_111_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_901 ();
 DECAPx10_ASAP7_75t_R FILLER_111_926 ();
 DECAPx10_ASAP7_75t_R FILLER_111_948 ();
 DECAPx10_ASAP7_75t_R FILLER_111_970 ();
 DECAPx6_ASAP7_75t_R FILLER_111_992 ();
 FILLER_ASAP7_75t_R FILLER_111_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1045 ();
 FILLER_ASAP7_75t_R FILLER_111_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1069 ();
 FILLER_ASAP7_75t_R FILLER_111_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1085 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1099 ();
 FILLER_ASAP7_75t_R FILLER_111_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1111 ();
 FILLER_ASAP7_75t_R FILLER_111_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1216 ();
 FILLER_ASAP7_75t_R FILLER_111_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1242 ();
 FILLER_ASAP7_75t_R FILLER_111_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1277 ();
 FILLER_ASAP7_75t_R FILLER_111_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_112_2 ();
 DECAPx4_ASAP7_75t_R FILLER_112_24 ();
 DECAPx1_ASAP7_75t_R FILLER_112_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_69 ();
 DECAPx1_ASAP7_75t_R FILLER_112_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_82 ();
 DECAPx10_ASAP7_75t_R FILLER_112_96 ();
 DECAPx1_ASAP7_75t_R FILLER_112_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_122 ();
 DECAPx2_ASAP7_75t_R FILLER_112_129 ();
 DECAPx1_ASAP7_75t_R FILLER_112_141 ();
 DECAPx2_ASAP7_75t_R FILLER_112_167 ();
 FILLER_ASAP7_75t_R FILLER_112_173 ();
 DECAPx4_ASAP7_75t_R FILLER_112_186 ();
 DECAPx2_ASAP7_75t_R FILLER_112_202 ();
 FILLER_ASAP7_75t_R FILLER_112_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_210 ();
 DECAPx2_ASAP7_75t_R FILLER_112_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_234 ();
 DECAPx2_ASAP7_75t_R FILLER_112_255 ();
 FILLER_ASAP7_75t_R FILLER_112_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_263 ();
 DECAPx2_ASAP7_75t_R FILLER_112_277 ();
 DECAPx1_ASAP7_75t_R FILLER_112_290 ();
 FILLER_ASAP7_75t_R FILLER_112_304 ();
 DECAPx1_ASAP7_75t_R FILLER_112_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_323 ();
 DECAPx10_ASAP7_75t_R FILLER_112_341 ();
 DECAPx4_ASAP7_75t_R FILLER_112_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_373 ();
 DECAPx4_ASAP7_75t_R FILLER_112_384 ();
 DECAPx2_ASAP7_75t_R FILLER_112_404 ();
 FILLER_ASAP7_75t_R FILLER_112_410 ();
 DECAPx10_ASAP7_75t_R FILLER_112_422 ();
 DECAPx4_ASAP7_75t_R FILLER_112_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_454 ();
 DECAPx10_ASAP7_75t_R FILLER_112_464 ();
 DECAPx2_ASAP7_75t_R FILLER_112_486 ();
 FILLER_ASAP7_75t_R FILLER_112_492 ();
 DECAPx10_ASAP7_75t_R FILLER_112_532 ();
 DECAPx10_ASAP7_75t_R FILLER_112_554 ();
 DECAPx6_ASAP7_75t_R FILLER_112_576 ();
 DECAPx1_ASAP7_75t_R FILLER_112_590 ();
 FILLER_ASAP7_75t_R FILLER_112_601 ();
 DECAPx10_ASAP7_75t_R FILLER_112_610 ();
 DECAPx4_ASAP7_75t_R FILLER_112_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_642 ();
 FILLER_ASAP7_75t_R FILLER_112_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_663 ();
 DECAPx4_ASAP7_75t_R FILLER_112_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_680 ();
 FILLER_ASAP7_75t_R FILLER_112_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_693 ();
 DECAPx10_ASAP7_75t_R FILLER_112_724 ();
 DECAPx10_ASAP7_75t_R FILLER_112_746 ();
 FILLER_ASAP7_75t_R FILLER_112_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_770 ();
 DECAPx10_ASAP7_75t_R FILLER_112_777 ();
 DECAPx10_ASAP7_75t_R FILLER_112_799 ();
 DECAPx6_ASAP7_75t_R FILLER_112_821 ();
 FILLER_ASAP7_75t_R FILLER_112_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_837 ();
 DECAPx2_ASAP7_75t_R FILLER_112_854 ();
 FILLER_ASAP7_75t_R FILLER_112_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_862 ();
 DECAPx10_ASAP7_75t_R FILLER_112_873 ();
 FILLER_ASAP7_75t_R FILLER_112_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_897 ();
 DECAPx10_ASAP7_75t_R FILLER_112_912 ();
 DECAPx10_ASAP7_75t_R FILLER_112_934 ();
 DECAPx6_ASAP7_75t_R FILLER_112_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_970 ();
 DECAPx1_ASAP7_75t_R FILLER_112_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1078 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_112_1124 ();
 FILLER_ASAP7_75t_R FILLER_112_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1211 ();
 FILLER_ASAP7_75t_R FILLER_112_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1230 ();
 FILLER_ASAP7_75t_R FILLER_112_1236 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1245 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_113_2 ();
 DECAPx4_ASAP7_75t_R FILLER_113_24 ();
 FILLER_ASAP7_75t_R FILLER_113_34 ();
 DECAPx2_ASAP7_75t_R FILLER_113_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_75 ();
 DECAPx1_ASAP7_75t_R FILLER_113_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_88 ();
 DECAPx2_ASAP7_75t_R FILLER_113_103 ();
 FILLER_ASAP7_75t_R FILLER_113_109 ();
 FILLER_ASAP7_75t_R FILLER_113_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_119 ();
 DECAPx6_ASAP7_75t_R FILLER_113_126 ();
 DECAPx1_ASAP7_75t_R FILLER_113_140 ();
 DECAPx1_ASAP7_75t_R FILLER_113_152 ();
 DECAPx1_ASAP7_75t_R FILLER_113_164 ();
 FILLER_ASAP7_75t_R FILLER_113_174 ();
 DECAPx2_ASAP7_75t_R FILLER_113_195 ();
 DECAPx4_ASAP7_75t_R FILLER_113_204 ();
 FILLER_ASAP7_75t_R FILLER_113_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_216 ();
 FILLER_ASAP7_75t_R FILLER_113_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_222 ();
 DECAPx1_ASAP7_75t_R FILLER_113_243 ();
 FILLER_ASAP7_75t_R FILLER_113_257 ();
 FILLER_ASAP7_75t_R FILLER_113_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_283 ();
 DECAPx2_ASAP7_75t_R FILLER_113_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_306 ();
 DECAPx2_ASAP7_75t_R FILLER_113_314 ();
 FILLER_ASAP7_75t_R FILLER_113_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_322 ();
 FILLER_ASAP7_75t_R FILLER_113_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_331 ();
 DECAPx10_ASAP7_75t_R FILLER_113_354 ();
 DECAPx4_ASAP7_75t_R FILLER_113_386 ();
 DECAPx2_ASAP7_75t_R FILLER_113_402 ();
 DECAPx10_ASAP7_75t_R FILLER_113_418 ();
 DECAPx10_ASAP7_75t_R FILLER_113_440 ();
 DECAPx6_ASAP7_75t_R FILLER_113_462 ();
 DECAPx2_ASAP7_75t_R FILLER_113_476 ();
 FILLER_ASAP7_75t_R FILLER_113_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_505 ();
 FILLER_ASAP7_75t_R FILLER_113_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_515 ();
 DECAPx6_ASAP7_75t_R FILLER_113_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_551 ();
 DECAPx10_ASAP7_75t_R FILLER_113_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_584 ();
 DECAPx2_ASAP7_75t_R FILLER_113_595 ();
 FILLER_ASAP7_75t_R FILLER_113_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_603 ();
 DECAPx6_ASAP7_75t_R FILLER_113_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_624 ();
 FILLER_ASAP7_75t_R FILLER_113_649 ();
 DECAPx10_ASAP7_75t_R FILLER_113_663 ();
 DECAPx10_ASAP7_75t_R FILLER_113_685 ();
 DECAPx4_ASAP7_75t_R FILLER_113_707 ();
 DECAPx4_ASAP7_75t_R FILLER_113_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_733 ();
 DECAPx6_ASAP7_75t_R FILLER_113_746 ();
 DECAPx1_ASAP7_75t_R FILLER_113_760 ();
 DECAPx10_ASAP7_75t_R FILLER_113_770 ();
 DECAPx10_ASAP7_75t_R FILLER_113_792 ();
 DECAPx10_ASAP7_75t_R FILLER_113_814 ();
 DECAPx1_ASAP7_75t_R FILLER_113_836 ();
 DECAPx10_ASAP7_75t_R FILLER_113_849 ();
 DECAPx10_ASAP7_75t_R FILLER_113_871 ();
 DECAPx4_ASAP7_75t_R FILLER_113_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_903 ();
 DECAPx6_ASAP7_75t_R FILLER_113_907 ();
 FILLER_ASAP7_75t_R FILLER_113_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_923 ();
 DECAPx4_ASAP7_75t_R FILLER_113_926 ();
 DECAPx10_ASAP7_75t_R FILLER_113_942 ();
 DECAPx10_ASAP7_75t_R FILLER_113_964 ();
 DECAPx6_ASAP7_75t_R FILLER_113_986 ();
 FILLER_ASAP7_75t_R FILLER_113_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1030 ();
 FILLER_ASAP7_75t_R FILLER_113_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1086 ();
 FILLER_ASAP7_75t_R FILLER_113_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1150 ();
 FILLER_ASAP7_75t_R FILLER_113_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1200 ();
 FILLER_ASAP7_75t_R FILLER_113_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1252 ();
 FILLER_ASAP7_75t_R FILLER_113_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_114_2 ();
 DECAPx2_ASAP7_75t_R FILLER_114_16 ();
 DECAPx2_ASAP7_75t_R FILLER_114_30 ();
 FILLER_ASAP7_75t_R FILLER_114_36 ();
 DECAPx1_ASAP7_75t_R FILLER_114_92 ();
 FILLER_ASAP7_75t_R FILLER_114_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_167 ();
 DECAPx2_ASAP7_75t_R FILLER_114_174 ();
 FILLER_ASAP7_75t_R FILLER_114_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_182 ();
 DECAPx4_ASAP7_75t_R FILLER_114_186 ();
 DECAPx6_ASAP7_75t_R FILLER_114_199 ();
 DECAPx2_ASAP7_75t_R FILLER_114_213 ();
 DECAPx6_ASAP7_75t_R FILLER_114_222 ();
 FILLER_ASAP7_75t_R FILLER_114_236 ();
 DECAPx10_ASAP7_75t_R FILLER_114_244 ();
 FILLER_ASAP7_75t_R FILLER_114_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_268 ();
 DECAPx10_ASAP7_75t_R FILLER_114_276 ();
 DECAPx10_ASAP7_75t_R FILLER_114_298 ();
 DECAPx6_ASAP7_75t_R FILLER_114_320 ();
 DECAPx2_ASAP7_75t_R FILLER_114_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_340 ();
 FILLER_ASAP7_75t_R FILLER_114_348 ();
 DECAPx1_ASAP7_75t_R FILLER_114_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_360 ();
 FILLER_ASAP7_75t_R FILLER_114_379 ();
 DECAPx10_ASAP7_75t_R FILLER_114_411 ();
 DECAPx4_ASAP7_75t_R FILLER_114_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_443 ();
 DECAPx6_ASAP7_75t_R FILLER_114_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_478 ();
 DECAPx1_ASAP7_75t_R FILLER_114_489 ();
 FILLER_ASAP7_75t_R FILLER_114_514 ();
 DECAPx6_ASAP7_75t_R FILLER_114_533 ();
 DECAPx2_ASAP7_75t_R FILLER_114_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_553 ();
 DECAPx10_ASAP7_75t_R FILLER_114_566 ();
 DECAPx10_ASAP7_75t_R FILLER_114_588 ();
 DECAPx2_ASAP7_75t_R FILLER_114_610 ();
 FILLER_ASAP7_75t_R FILLER_114_616 ();
 DECAPx10_ASAP7_75t_R FILLER_114_628 ();
 DECAPx10_ASAP7_75t_R FILLER_114_650 ();
 DECAPx10_ASAP7_75t_R FILLER_114_672 ();
 DECAPx10_ASAP7_75t_R FILLER_114_694 ();
 DECAPx10_ASAP7_75t_R FILLER_114_716 ();
 DECAPx10_ASAP7_75t_R FILLER_114_738 ();
 DECAPx10_ASAP7_75t_R FILLER_114_760 ();
 FILLER_ASAP7_75t_R FILLER_114_782 ();
 DECAPx1_ASAP7_75t_R FILLER_114_790 ();
 DECAPx6_ASAP7_75t_R FILLER_114_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_814 ();
 DECAPx10_ASAP7_75t_R FILLER_114_821 ();
 DECAPx1_ASAP7_75t_R FILLER_114_843 ();
 DECAPx2_ASAP7_75t_R FILLER_114_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_859 ();
 DECAPx2_ASAP7_75t_R FILLER_114_868 ();
 FILLER_ASAP7_75t_R FILLER_114_874 ();
 DECAPx10_ASAP7_75t_R FILLER_114_890 ();
 DECAPx10_ASAP7_75t_R FILLER_114_912 ();
 DECAPx2_ASAP7_75t_R FILLER_114_934 ();
 DECAPx6_ASAP7_75t_R FILLER_114_948 ();
 DECAPx1_ASAP7_75t_R FILLER_114_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_966 ();
 DECAPx4_ASAP7_75t_R FILLER_114_973 ();
 DECAPx6_ASAP7_75t_R FILLER_114_989 ();
 FILLER_ASAP7_75t_R FILLER_114_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1013 ();
 FILLER_ASAP7_75t_R FILLER_114_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1225 ();
 FILLER_ASAP7_75t_R FILLER_114_1235 ();
 FILLER_ASAP7_75t_R FILLER_114_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1270 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_115_2 ();
 DECAPx10_ASAP7_75t_R FILLER_115_24 ();
 DECAPx10_ASAP7_75t_R FILLER_115_46 ();
 DECAPx6_ASAP7_75t_R FILLER_115_68 ();
 FILLER_ASAP7_75t_R FILLER_115_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_84 ();
 FILLER_ASAP7_75t_R FILLER_115_106 ();
 DECAPx2_ASAP7_75t_R FILLER_115_126 ();
 DECAPx10_ASAP7_75t_R FILLER_115_160 ();
 DECAPx10_ASAP7_75t_R FILLER_115_182 ();
 DECAPx10_ASAP7_75t_R FILLER_115_207 ();
 DECAPx6_ASAP7_75t_R FILLER_115_229 ();
 DECAPx1_ASAP7_75t_R FILLER_115_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_247 ();
 DECAPx1_ASAP7_75t_R FILLER_115_264 ();
 DECAPx2_ASAP7_75t_R FILLER_115_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_288 ();
 DECAPx10_ASAP7_75t_R FILLER_115_296 ();
 DECAPx2_ASAP7_75t_R FILLER_115_318 ();
 FILLER_ASAP7_75t_R FILLER_115_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_336 ();
 DECAPx10_ASAP7_75t_R FILLER_115_356 ();
 DECAPx2_ASAP7_75t_R FILLER_115_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_384 ();
 FILLER_ASAP7_75t_R FILLER_115_395 ();
 DECAPx4_ASAP7_75t_R FILLER_115_407 ();
 DECAPx10_ASAP7_75t_R FILLER_115_437 ();
 DECAPx6_ASAP7_75t_R FILLER_115_459 ();
 DECAPx2_ASAP7_75t_R FILLER_115_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_505 ();
 DECAPx4_ASAP7_75t_R FILLER_115_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_526 ();
 DECAPx10_ASAP7_75t_R FILLER_115_537 ();
 DECAPx10_ASAP7_75t_R FILLER_115_559 ();
 FILLER_ASAP7_75t_R FILLER_115_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_583 ();
 DECAPx10_ASAP7_75t_R FILLER_115_590 ();
 DECAPx2_ASAP7_75t_R FILLER_115_612 ();
 FILLER_ASAP7_75t_R FILLER_115_618 ();
 DECAPx4_ASAP7_75t_R FILLER_115_626 ();
 FILLER_ASAP7_75t_R FILLER_115_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_638 ();
 DECAPx10_ASAP7_75t_R FILLER_115_651 ();
 DECAPx10_ASAP7_75t_R FILLER_115_673 ();
 DECAPx6_ASAP7_75t_R FILLER_115_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_709 ();
 DECAPx2_ASAP7_75t_R FILLER_115_716 ();
 FILLER_ASAP7_75t_R FILLER_115_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_724 ();
 DECAPx10_ASAP7_75t_R FILLER_115_731 ();
 DECAPx10_ASAP7_75t_R FILLER_115_753 ();
 DECAPx4_ASAP7_75t_R FILLER_115_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_785 ();
 DECAPx6_ASAP7_75t_R FILLER_115_792 ();
 DECAPx10_ASAP7_75t_R FILLER_115_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_834 ();
 DECAPx2_ASAP7_75t_R FILLER_115_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_859 ();
 DECAPx10_ASAP7_75t_R FILLER_115_866 ();
 FILLER_ASAP7_75t_R FILLER_115_895 ();
 DECAPx2_ASAP7_75t_R FILLER_115_936 ();
 FILLER_ASAP7_75t_R FILLER_115_942 ();
 DECAPx1_ASAP7_75t_R FILLER_115_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_960 ();
 DECAPx10_ASAP7_75t_R FILLER_115_971 ();
 DECAPx10_ASAP7_75t_R FILLER_115_993 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1015 ();
 FILLER_ASAP7_75t_R FILLER_115_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_115_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1090 ();
 FILLER_ASAP7_75t_R FILLER_115_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1122 ();
 FILLER_ASAP7_75t_R FILLER_115_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1150 ();
 FILLER_ASAP7_75t_R FILLER_115_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1162 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1197 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1226 ();
 FILLER_ASAP7_75t_R FILLER_115_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1250 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_116_2 ();
 DECAPx10_ASAP7_75t_R FILLER_116_24 ();
 DECAPx10_ASAP7_75t_R FILLER_116_46 ();
 DECAPx10_ASAP7_75t_R FILLER_116_68 ();
 DECAPx10_ASAP7_75t_R FILLER_116_90 ();
 DECAPx6_ASAP7_75t_R FILLER_116_112 ();
 DECAPx2_ASAP7_75t_R FILLER_116_134 ();
 FILLER_ASAP7_75t_R FILLER_116_140 ();
 DECAPx10_ASAP7_75t_R FILLER_116_150 ();
 DECAPx1_ASAP7_75t_R FILLER_116_172 ();
 DECAPx4_ASAP7_75t_R FILLER_116_179 ();
 DECAPx6_ASAP7_75t_R FILLER_116_202 ();
 FILLER_ASAP7_75t_R FILLER_116_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_255 ();
 FILLER_ASAP7_75t_R FILLER_116_266 ();
 FILLER_ASAP7_75t_R FILLER_116_278 ();
 DECAPx6_ASAP7_75t_R FILLER_116_294 ();
 FILLER_ASAP7_75t_R FILLER_116_315 ();
 DECAPx6_ASAP7_75t_R FILLER_116_329 ();
 FILLER_ASAP7_75t_R FILLER_116_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_345 ();
 FILLER_ASAP7_75t_R FILLER_116_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_355 ();
 DECAPx2_ASAP7_75t_R FILLER_116_364 ();
 FILLER_ASAP7_75t_R FILLER_116_370 ();
 FILLER_ASAP7_75t_R FILLER_116_382 ();
 DECAPx2_ASAP7_75t_R FILLER_116_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_426 ();
 DECAPx10_ASAP7_75t_R FILLER_116_437 ();
 FILLER_ASAP7_75t_R FILLER_116_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_461 ();
 DECAPx10_ASAP7_75t_R FILLER_116_464 ();
 DECAPx6_ASAP7_75t_R FILLER_116_486 ();
 DECAPx1_ASAP7_75t_R FILLER_116_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_504 ();
 DECAPx10_ASAP7_75t_R FILLER_116_533 ();
 DECAPx10_ASAP7_75t_R FILLER_116_555 ();
 FILLER_ASAP7_75t_R FILLER_116_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_592 ();
 DECAPx4_ASAP7_75t_R FILLER_116_599 ();
 FILLER_ASAP7_75t_R FILLER_116_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_611 ();
 DECAPx2_ASAP7_75t_R FILLER_116_633 ();
 FILLER_ASAP7_75t_R FILLER_116_639 ();
 DECAPx2_ASAP7_75t_R FILLER_116_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_668 ();
 DECAPx10_ASAP7_75t_R FILLER_116_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_734 ();
 DECAPx10_ASAP7_75t_R FILLER_116_741 ();
 DECAPx10_ASAP7_75t_R FILLER_116_763 ();
 DECAPx10_ASAP7_75t_R FILLER_116_785 ();
 DECAPx10_ASAP7_75t_R FILLER_116_807 ();
 DECAPx1_ASAP7_75t_R FILLER_116_829 ();
 DECAPx10_ASAP7_75t_R FILLER_116_857 ();
 DECAPx6_ASAP7_75t_R FILLER_116_879 ();
 DECAPx1_ASAP7_75t_R FILLER_116_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_897 ();
 DECAPx1_ASAP7_75t_R FILLER_116_910 ();
 DECAPx10_ASAP7_75t_R FILLER_116_923 ();
 DECAPx10_ASAP7_75t_R FILLER_116_945 ();
 DECAPx6_ASAP7_75t_R FILLER_116_967 ();
 DECAPx1_ASAP7_75t_R FILLER_116_981 ();
 DECAPx2_ASAP7_75t_R FILLER_116_995 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1029 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1077 ();
 FILLER_ASAP7_75t_R FILLER_116_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1111 ();
 FILLER_ASAP7_75t_R FILLER_116_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1216 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1238 ();
 FILLER_ASAP7_75t_R FILLER_116_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_117_2 ();
 DECAPx10_ASAP7_75t_R FILLER_117_24 ();
 DECAPx10_ASAP7_75t_R FILLER_117_46 ();
 DECAPx10_ASAP7_75t_R FILLER_117_68 ();
 DECAPx10_ASAP7_75t_R FILLER_117_90 ();
 DECAPx6_ASAP7_75t_R FILLER_117_112 ();
 DECAPx1_ASAP7_75t_R FILLER_117_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_130 ();
 DECAPx2_ASAP7_75t_R FILLER_117_159 ();
 FILLER_ASAP7_75t_R FILLER_117_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_167 ();
 DECAPx2_ASAP7_75t_R FILLER_117_171 ();
 FILLER_ASAP7_75t_R FILLER_117_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_179 ();
 FILLER_ASAP7_75t_R FILLER_117_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_185 ();
 DECAPx2_ASAP7_75t_R FILLER_117_208 ();
 FILLER_ASAP7_75t_R FILLER_117_214 ();
 DECAPx2_ASAP7_75t_R FILLER_117_226 ();
 DECAPx4_ASAP7_75t_R FILLER_117_248 ();
 FILLER_ASAP7_75t_R FILLER_117_258 ();
 DECAPx10_ASAP7_75t_R FILLER_117_282 ();
 FILLER_ASAP7_75t_R FILLER_117_304 ();
 DECAPx10_ASAP7_75t_R FILLER_117_316 ();
 DECAPx2_ASAP7_75t_R FILLER_117_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_344 ();
 FILLER_ASAP7_75t_R FILLER_117_352 ();
 DECAPx2_ASAP7_75t_R FILLER_117_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_427 ();
 DECAPx1_ASAP7_75t_R FILLER_117_438 ();
 DECAPx6_ASAP7_75t_R FILLER_117_464 ();
 FILLER_ASAP7_75t_R FILLER_117_478 ();
 DECAPx10_ASAP7_75t_R FILLER_117_498 ();
 DECAPx2_ASAP7_75t_R FILLER_117_520 ();
 DECAPx6_ASAP7_75t_R FILLER_117_547 ();
 DECAPx2_ASAP7_75t_R FILLER_117_561 ();
 DECAPx1_ASAP7_75t_R FILLER_117_615 ();
 DECAPx6_ASAP7_75t_R FILLER_117_625 ();
 DECAPx1_ASAP7_75t_R FILLER_117_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_643 ();
 DECAPx4_ASAP7_75t_R FILLER_117_656 ();
 FILLER_ASAP7_75t_R FILLER_117_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_706 ();
 DECAPx10_ASAP7_75t_R FILLER_117_737 ();
 DECAPx10_ASAP7_75t_R FILLER_117_759 ();
 DECAPx10_ASAP7_75t_R FILLER_117_781 ();
 DECAPx10_ASAP7_75t_R FILLER_117_803 ();
 DECAPx6_ASAP7_75t_R FILLER_117_825 ();
 DECAPx2_ASAP7_75t_R FILLER_117_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_845 ();
 DECAPx6_ASAP7_75t_R FILLER_117_858 ();
 DECAPx2_ASAP7_75t_R FILLER_117_872 ();
 DECAPx2_ASAP7_75t_R FILLER_117_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_902 ();
 DECAPx10_ASAP7_75t_R FILLER_117_926 ();
 DECAPx6_ASAP7_75t_R FILLER_117_948 ();
 FILLER_ASAP7_75t_R FILLER_117_962 ();
 DECAPx4_ASAP7_75t_R FILLER_117_972 ();
 FILLER_ASAP7_75t_R FILLER_117_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_996 ();
 FILLER_ASAP7_75t_R FILLER_117_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1142 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1167 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1248 ();
 FILLER_ASAP7_75t_R FILLER_117_1270 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_118_2 ();
 DECAPx10_ASAP7_75t_R FILLER_118_24 ();
 DECAPx10_ASAP7_75t_R FILLER_118_46 ();
 DECAPx10_ASAP7_75t_R FILLER_118_68 ();
 DECAPx10_ASAP7_75t_R FILLER_118_90 ();
 DECAPx10_ASAP7_75t_R FILLER_118_112 ();
 DECAPx10_ASAP7_75t_R FILLER_118_134 ();
 DECAPx10_ASAP7_75t_R FILLER_118_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_178 ();
 DECAPx2_ASAP7_75t_R FILLER_118_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_188 ();
 DECAPx2_ASAP7_75t_R FILLER_118_198 ();
 FILLER_ASAP7_75t_R FILLER_118_224 ();
 DECAPx2_ASAP7_75t_R FILLER_118_232 ();
 DECAPx1_ASAP7_75t_R FILLER_118_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_264 ();
 DECAPx2_ASAP7_75t_R FILLER_118_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_293 ();
 DECAPx2_ASAP7_75t_R FILLER_118_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_317 ();
 DECAPx4_ASAP7_75t_R FILLER_118_324 ();
 DECAPx2_ASAP7_75t_R FILLER_118_341 ();
 DECAPx10_ASAP7_75t_R FILLER_118_357 ();
 DECAPx6_ASAP7_75t_R FILLER_118_379 ();
 DECAPx2_ASAP7_75t_R FILLER_118_393 ();
 DECAPx10_ASAP7_75t_R FILLER_118_423 ();
 DECAPx6_ASAP7_75t_R FILLER_118_445 ();
 FILLER_ASAP7_75t_R FILLER_118_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_461 ();
 FILLER_ASAP7_75t_R FILLER_118_464 ();
 DECAPx1_ASAP7_75t_R FILLER_118_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_496 ();
 DECAPx4_ASAP7_75t_R FILLER_118_512 ();
 DECAPx6_ASAP7_75t_R FILLER_118_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_550 ();
 DECAPx1_ASAP7_75t_R FILLER_118_572 ();
 FILLER_ASAP7_75t_R FILLER_118_606 ();
 DECAPx6_ASAP7_75t_R FILLER_118_620 ();
 FILLER_ASAP7_75t_R FILLER_118_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_657 ();
 DECAPx10_ASAP7_75t_R FILLER_118_679 ();
 DECAPx10_ASAP7_75t_R FILLER_118_701 ();
 DECAPx10_ASAP7_75t_R FILLER_118_723 ();
 DECAPx6_ASAP7_75t_R FILLER_118_745 ();
 FILLER_ASAP7_75t_R FILLER_118_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_761 ();
 DECAPx2_ASAP7_75t_R FILLER_118_772 ();
 FILLER_ASAP7_75t_R FILLER_118_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_780 ();
 DECAPx10_ASAP7_75t_R FILLER_118_787 ();
 DECAPx10_ASAP7_75t_R FILLER_118_809 ();
 DECAPx10_ASAP7_75t_R FILLER_118_831 ();
 DECAPx4_ASAP7_75t_R FILLER_118_853 ();
 FILLER_ASAP7_75t_R FILLER_118_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_865 ();
 DECAPx2_ASAP7_75t_R FILLER_118_872 ();
 FILLER_ASAP7_75t_R FILLER_118_902 ();
 DECAPx10_ASAP7_75t_R FILLER_118_916 ();
 DECAPx10_ASAP7_75t_R FILLER_118_938 ();
 DECAPx1_ASAP7_75t_R FILLER_118_960 ();
 DECAPx2_ASAP7_75t_R FILLER_118_980 ();
 FILLER_ASAP7_75t_R FILLER_118_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_988 ();
 FILLER_ASAP7_75t_R FILLER_118_995 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1100 ();
 FILLER_ASAP7_75t_R FILLER_118_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1144 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1167 ();
 FILLER_ASAP7_75t_R FILLER_118_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1186 ();
 FILLER_ASAP7_75t_R FILLER_118_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1212 ();
 FILLER_ASAP7_75t_R FILLER_118_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1285 ();
 FILLER_ASAP7_75t_R FILLER_118_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_119_2 ();
 DECAPx10_ASAP7_75t_R FILLER_119_24 ();
 DECAPx10_ASAP7_75t_R FILLER_119_46 ();
 DECAPx10_ASAP7_75t_R FILLER_119_68 ();
 DECAPx10_ASAP7_75t_R FILLER_119_90 ();
 DECAPx10_ASAP7_75t_R FILLER_119_112 ();
 DECAPx10_ASAP7_75t_R FILLER_119_134 ();
 DECAPx6_ASAP7_75t_R FILLER_119_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_170 ();
 DECAPx10_ASAP7_75t_R FILLER_119_174 ();
 DECAPx10_ASAP7_75t_R FILLER_119_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_218 ();
 DECAPx10_ASAP7_75t_R FILLER_119_225 ();
 DECAPx10_ASAP7_75t_R FILLER_119_247 ();
 DECAPx4_ASAP7_75t_R FILLER_119_269 ();
 FILLER_ASAP7_75t_R FILLER_119_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_281 ();
 DECAPx10_ASAP7_75t_R FILLER_119_285 ();
 DECAPx2_ASAP7_75t_R FILLER_119_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_313 ();
 DECAPx10_ASAP7_75t_R FILLER_119_351 ();
 DECAPx10_ASAP7_75t_R FILLER_119_373 ();
 DECAPx6_ASAP7_75t_R FILLER_119_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_409 ();
 DECAPx10_ASAP7_75t_R FILLER_119_430 ();
 DECAPx10_ASAP7_75t_R FILLER_119_452 ();
 DECAPx10_ASAP7_75t_R FILLER_119_474 ();
 DECAPx10_ASAP7_75t_R FILLER_119_496 ();
 DECAPx1_ASAP7_75t_R FILLER_119_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_522 ();
 DECAPx6_ASAP7_75t_R FILLER_119_533 ();
 FILLER_ASAP7_75t_R FILLER_119_547 ();
 DECAPx4_ASAP7_75t_R FILLER_119_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_624 ();
 FILLER_ASAP7_75t_R FILLER_119_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_657 ();
 DECAPx6_ASAP7_75t_R FILLER_119_670 ();
 DECAPx2_ASAP7_75t_R FILLER_119_722 ();
 FILLER_ASAP7_75t_R FILLER_119_728 ();
 DECAPx1_ASAP7_75t_R FILLER_119_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_761 ();
 DECAPx4_ASAP7_75t_R FILLER_119_772 ();
 FILLER_ASAP7_75t_R FILLER_119_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_784 ();
 DECAPx6_ASAP7_75t_R FILLER_119_808 ();
 FILLER_ASAP7_75t_R FILLER_119_822 ();
 DECAPx10_ASAP7_75t_R FILLER_119_832 ();
 DECAPx10_ASAP7_75t_R FILLER_119_854 ();
 DECAPx6_ASAP7_75t_R FILLER_119_904 ();
 DECAPx2_ASAP7_75t_R FILLER_119_918 ();
 DECAPx2_ASAP7_75t_R FILLER_119_926 ();
 FILLER_ASAP7_75t_R FILLER_119_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_934 ();
 DECAPx10_ASAP7_75t_R FILLER_119_947 ();
 FILLER_ASAP7_75t_R FILLER_119_969 ();
 DECAPx10_ASAP7_75t_R FILLER_119_977 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1049 ();
 FILLER_ASAP7_75t_R FILLER_119_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_119_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1113 ();
 FILLER_ASAP7_75t_R FILLER_119_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1138 ();
 FILLER_ASAP7_75t_R FILLER_119_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1146 ();
 FILLER_ASAP7_75t_R FILLER_119_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1228 ();
 FILLER_ASAP7_75t_R FILLER_119_1242 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_120_2 ();
 DECAPx10_ASAP7_75t_R FILLER_120_24 ();
 DECAPx10_ASAP7_75t_R FILLER_120_46 ();
 DECAPx10_ASAP7_75t_R FILLER_120_68 ();
 DECAPx10_ASAP7_75t_R FILLER_120_90 ();
 DECAPx10_ASAP7_75t_R FILLER_120_112 ();
 DECAPx10_ASAP7_75t_R FILLER_120_134 ();
 DECAPx10_ASAP7_75t_R FILLER_120_156 ();
 DECAPx6_ASAP7_75t_R FILLER_120_178 ();
 FILLER_ASAP7_75t_R FILLER_120_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_194 ();
 DECAPx10_ASAP7_75t_R FILLER_120_198 ();
 DECAPx10_ASAP7_75t_R FILLER_120_220 ();
 DECAPx10_ASAP7_75t_R FILLER_120_242 ();
 DECAPx10_ASAP7_75t_R FILLER_120_264 ();
 DECAPx4_ASAP7_75t_R FILLER_120_286 ();
 FILLER_ASAP7_75t_R FILLER_120_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_327 ();
 DECAPx10_ASAP7_75t_R FILLER_120_338 ();
 DECAPx2_ASAP7_75t_R FILLER_120_360 ();
 FILLER_ASAP7_75t_R FILLER_120_366 ();
 DECAPx10_ASAP7_75t_R FILLER_120_398 ();
 DECAPx10_ASAP7_75t_R FILLER_120_420 ();
 DECAPx6_ASAP7_75t_R FILLER_120_442 ();
 DECAPx2_ASAP7_75t_R FILLER_120_456 ();
 DECAPx10_ASAP7_75t_R FILLER_120_464 ();
 DECAPx10_ASAP7_75t_R FILLER_120_486 ();
 DECAPx6_ASAP7_75t_R FILLER_120_508 ();
 DECAPx2_ASAP7_75t_R FILLER_120_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_528 ();
 DECAPx2_ASAP7_75t_R FILLER_120_591 ();
 FILLER_ASAP7_75t_R FILLER_120_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_599 ();
 DECAPx6_ASAP7_75t_R FILLER_120_621 ();
 DECAPx1_ASAP7_75t_R FILLER_120_635 ();
 DECAPx6_ASAP7_75t_R FILLER_120_655 ();
 FILLER_ASAP7_75t_R FILLER_120_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_671 ();
 DECAPx6_ASAP7_75t_R FILLER_120_688 ();
 FILLER_ASAP7_75t_R FILLER_120_702 ();
 DECAPx1_ASAP7_75t_R FILLER_120_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_729 ();
 DECAPx2_ASAP7_75t_R FILLER_120_742 ();
 FILLER_ASAP7_75t_R FILLER_120_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_750 ();
 FILLER_ASAP7_75t_R FILLER_120_757 ();
 DECAPx4_ASAP7_75t_R FILLER_120_771 ();
 FILLER_ASAP7_75t_R FILLER_120_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_789 ();
 DECAPx6_ASAP7_75t_R FILLER_120_800 ();
 DECAPx2_ASAP7_75t_R FILLER_120_814 ();
 DECAPx6_ASAP7_75t_R FILLER_120_840 ();
 DECAPx2_ASAP7_75t_R FILLER_120_854 ();
 DECAPx6_ASAP7_75t_R FILLER_120_866 ();
 DECAPx10_ASAP7_75t_R FILLER_120_908 ();
 DECAPx4_ASAP7_75t_R FILLER_120_930 ();
 FILLER_ASAP7_75t_R FILLER_120_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_942 ();
 DECAPx10_ASAP7_75t_R FILLER_120_952 ();
 DECAPx6_ASAP7_75t_R FILLER_120_974 ();
 FILLER_ASAP7_75t_R FILLER_120_988 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1032 ();
 FILLER_ASAP7_75t_R FILLER_120_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1067 ();
 FILLER_ASAP7_75t_R FILLER_120_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1090 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1140 ();
 FILLER_ASAP7_75t_R FILLER_120_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1178 ();
 DECAPx6_ASAP7_75t_R FILLER_120_1189 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1216 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_121_2 ();
 DECAPx10_ASAP7_75t_R FILLER_121_24 ();
 DECAPx10_ASAP7_75t_R FILLER_121_46 ();
 DECAPx10_ASAP7_75t_R FILLER_121_68 ();
 DECAPx10_ASAP7_75t_R FILLER_121_90 ();
 DECAPx10_ASAP7_75t_R FILLER_121_112 ();
 DECAPx10_ASAP7_75t_R FILLER_121_134 ();
 DECAPx10_ASAP7_75t_R FILLER_121_156 ();
 DECAPx10_ASAP7_75t_R FILLER_121_178 ();
 DECAPx1_ASAP7_75t_R FILLER_121_200 ();
 DECAPx10_ASAP7_75t_R FILLER_121_207 ();
 DECAPx6_ASAP7_75t_R FILLER_121_229 ();
 DECAPx2_ASAP7_75t_R FILLER_121_243 ();
 DECAPx4_ASAP7_75t_R FILLER_121_252 ();
 FILLER_ASAP7_75t_R FILLER_121_262 ();
 DECAPx10_ASAP7_75t_R FILLER_121_285 ();
 DECAPx4_ASAP7_75t_R FILLER_121_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_317 ();
 DECAPx2_ASAP7_75t_R FILLER_121_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_330 ();
 DECAPx10_ASAP7_75t_R FILLER_121_337 ();
 DECAPx6_ASAP7_75t_R FILLER_121_359 ();
 DECAPx2_ASAP7_75t_R FILLER_121_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_379 ();
 DECAPx10_ASAP7_75t_R FILLER_121_390 ();
 DECAPx10_ASAP7_75t_R FILLER_121_412 ();
 DECAPx10_ASAP7_75t_R FILLER_121_434 ();
 DECAPx10_ASAP7_75t_R FILLER_121_456 ();
 DECAPx10_ASAP7_75t_R FILLER_121_478 ();
 DECAPx10_ASAP7_75t_R FILLER_121_500 ();
 DECAPx10_ASAP7_75t_R FILLER_121_522 ();
 DECAPx10_ASAP7_75t_R FILLER_121_544 ();
 DECAPx1_ASAP7_75t_R FILLER_121_566 ();
 DECAPx10_ASAP7_75t_R FILLER_121_576 ();
 DECAPx2_ASAP7_75t_R FILLER_121_598 ();
 FILLER_ASAP7_75t_R FILLER_121_604 ();
 DECAPx10_ASAP7_75t_R FILLER_121_612 ();
 DECAPx4_ASAP7_75t_R FILLER_121_634 ();
 FILLER_ASAP7_75t_R FILLER_121_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_646 ();
 DECAPx10_ASAP7_75t_R FILLER_121_659 ();
 DECAPx10_ASAP7_75t_R FILLER_121_681 ();
 DECAPx4_ASAP7_75t_R FILLER_121_703 ();
 FILLER_ASAP7_75t_R FILLER_121_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_715 ();
 DECAPx10_ASAP7_75t_R FILLER_121_728 ();
 DECAPx10_ASAP7_75t_R FILLER_121_750 ();
 DECAPx10_ASAP7_75t_R FILLER_121_772 ();
 DECAPx6_ASAP7_75t_R FILLER_121_794 ();
 DECAPx1_ASAP7_75t_R FILLER_121_808 ();
 DECAPx10_ASAP7_75t_R FILLER_121_826 ();
 DECAPx6_ASAP7_75t_R FILLER_121_848 ();
 DECAPx2_ASAP7_75t_R FILLER_121_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_868 ();
 DECAPx2_ASAP7_75t_R FILLER_121_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_889 ();
 DECAPx1_ASAP7_75t_R FILLER_121_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_901 ();
 DECAPx1_ASAP7_75t_R FILLER_121_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_923 ();
 DECAPx10_ASAP7_75t_R FILLER_121_938 ();
 DECAPx10_ASAP7_75t_R FILLER_121_960 ();
 DECAPx2_ASAP7_75t_R FILLER_121_988 ();
 FILLER_ASAP7_75t_R FILLER_121_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_996 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1013 ();
 FILLER_ASAP7_75t_R FILLER_121_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1074 ();
 FILLER_ASAP7_75t_R FILLER_121_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1198 ();
 FILLER_ASAP7_75t_R FILLER_121_1204 ();
 FILLER_ASAP7_75t_R FILLER_121_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_121_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_122_2 ();
 DECAPx10_ASAP7_75t_R FILLER_122_24 ();
 DECAPx10_ASAP7_75t_R FILLER_122_46 ();
 DECAPx10_ASAP7_75t_R FILLER_122_68 ();
 DECAPx10_ASAP7_75t_R FILLER_122_90 ();
 DECAPx10_ASAP7_75t_R FILLER_122_112 ();
 DECAPx10_ASAP7_75t_R FILLER_122_134 ();
 DECAPx10_ASAP7_75t_R FILLER_122_156 ();
 DECAPx10_ASAP7_75t_R FILLER_122_178 ();
 DECAPx10_ASAP7_75t_R FILLER_122_200 ();
 DECAPx10_ASAP7_75t_R FILLER_122_222 ();
 DECAPx10_ASAP7_75t_R FILLER_122_244 ();
 DECAPx10_ASAP7_75t_R FILLER_122_266 ();
 DECAPx10_ASAP7_75t_R FILLER_122_288 ();
 DECAPx10_ASAP7_75t_R FILLER_122_310 ();
 DECAPx10_ASAP7_75t_R FILLER_122_332 ();
 DECAPx10_ASAP7_75t_R FILLER_122_354 ();
 DECAPx10_ASAP7_75t_R FILLER_122_376 ();
 DECAPx10_ASAP7_75t_R FILLER_122_398 ();
 DECAPx10_ASAP7_75t_R FILLER_122_420 ();
 DECAPx6_ASAP7_75t_R FILLER_122_442 ();
 DECAPx2_ASAP7_75t_R FILLER_122_456 ();
 DECAPx10_ASAP7_75t_R FILLER_122_464 ();
 DECAPx10_ASAP7_75t_R FILLER_122_486 ();
 DECAPx10_ASAP7_75t_R FILLER_122_508 ();
 DECAPx10_ASAP7_75t_R FILLER_122_530 ();
 DECAPx10_ASAP7_75t_R FILLER_122_552 ();
 DECAPx10_ASAP7_75t_R FILLER_122_574 ();
 DECAPx10_ASAP7_75t_R FILLER_122_596 ();
 DECAPx10_ASAP7_75t_R FILLER_122_618 ();
 DECAPx10_ASAP7_75t_R FILLER_122_640 ();
 DECAPx10_ASAP7_75t_R FILLER_122_662 ();
 DECAPx10_ASAP7_75t_R FILLER_122_684 ();
 DECAPx10_ASAP7_75t_R FILLER_122_706 ();
 DECAPx10_ASAP7_75t_R FILLER_122_728 ();
 DECAPx10_ASAP7_75t_R FILLER_122_750 ();
 DECAPx10_ASAP7_75t_R FILLER_122_772 ();
 DECAPx10_ASAP7_75t_R FILLER_122_794 ();
 DECAPx10_ASAP7_75t_R FILLER_122_816 ();
 DECAPx10_ASAP7_75t_R FILLER_122_838 ();
 FILLER_ASAP7_75t_R FILLER_122_860 ();
 DECAPx6_ASAP7_75t_R FILLER_122_874 ();
 DECAPx2_ASAP7_75t_R FILLER_122_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_894 ();
 DECAPx1_ASAP7_75t_R FILLER_122_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_919 ();
 DECAPx1_ASAP7_75t_R FILLER_122_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_936 ();
 DECAPx1_ASAP7_75t_R FILLER_122_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_944 ();
 DECAPx10_ASAP7_75t_R FILLER_122_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_977 ();
 DECAPx2_ASAP7_75t_R FILLER_122_988 ();
 FILLER_ASAP7_75t_R FILLER_122_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_996 ();
 FILLER_ASAP7_75t_R FILLER_122_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1086 ();
 FILLER_ASAP7_75t_R FILLER_122_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1114 ();
 FILLER_ASAP7_75t_R FILLER_122_1121 ();
 FILLER_ASAP7_75t_R FILLER_122_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1144 ();
 FILLER_ASAP7_75t_R FILLER_122_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1167 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1214 ();
 FILLER_ASAP7_75t_R FILLER_122_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1222 ();
 FILLER_ASAP7_75t_R FILLER_122_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_123_24 ();
 DECAPx10_ASAP7_75t_R FILLER_123_46 ();
 DECAPx10_ASAP7_75t_R FILLER_123_68 ();
 DECAPx10_ASAP7_75t_R FILLER_123_90 ();
 DECAPx10_ASAP7_75t_R FILLER_123_112 ();
 DECAPx10_ASAP7_75t_R FILLER_123_134 ();
 DECAPx10_ASAP7_75t_R FILLER_123_156 ();
 DECAPx10_ASAP7_75t_R FILLER_123_178 ();
 DECAPx10_ASAP7_75t_R FILLER_123_200 ();
 DECAPx10_ASAP7_75t_R FILLER_123_222 ();
 DECAPx10_ASAP7_75t_R FILLER_123_244 ();
 DECAPx10_ASAP7_75t_R FILLER_123_266 ();
 DECAPx10_ASAP7_75t_R FILLER_123_288 ();
 DECAPx10_ASAP7_75t_R FILLER_123_310 ();
 DECAPx10_ASAP7_75t_R FILLER_123_332 ();
 DECAPx10_ASAP7_75t_R FILLER_123_354 ();
 DECAPx10_ASAP7_75t_R FILLER_123_376 ();
 DECAPx10_ASAP7_75t_R FILLER_123_398 ();
 DECAPx10_ASAP7_75t_R FILLER_123_420 ();
 DECAPx6_ASAP7_75t_R FILLER_123_442 ();
 DECAPx2_ASAP7_75t_R FILLER_123_456 ();
 DECAPx10_ASAP7_75t_R FILLER_123_464 ();
 DECAPx10_ASAP7_75t_R FILLER_123_486 ();
 DECAPx10_ASAP7_75t_R FILLER_123_508 ();
 DECAPx10_ASAP7_75t_R FILLER_123_530 ();
 DECAPx10_ASAP7_75t_R FILLER_123_552 ();
 DECAPx10_ASAP7_75t_R FILLER_123_574 ();
 DECAPx10_ASAP7_75t_R FILLER_123_596 ();
 DECAPx10_ASAP7_75t_R FILLER_123_618 ();
 DECAPx10_ASAP7_75t_R FILLER_123_640 ();
 DECAPx10_ASAP7_75t_R FILLER_123_662 ();
 DECAPx10_ASAP7_75t_R FILLER_123_684 ();
 DECAPx10_ASAP7_75t_R FILLER_123_728 ();
 DECAPx10_ASAP7_75t_R FILLER_123_750 ();
 DECAPx10_ASAP7_75t_R FILLER_123_772 ();
 DECAPx10_ASAP7_75t_R FILLER_123_794 ();
 DECAPx10_ASAP7_75t_R FILLER_123_816 ();
 DECAPx10_ASAP7_75t_R FILLER_123_838 ();
 DECAPx10_ASAP7_75t_R FILLER_123_860 ();
 DECAPx10_ASAP7_75t_R FILLER_123_882 ();
 DECAPx6_ASAP7_75t_R FILLER_123_904 ();
 DECAPx2_ASAP7_75t_R FILLER_123_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_953 ();
 DECAPx2_ASAP7_75t_R FILLER_123_975 ();
 FILLER_ASAP7_75t_R FILLER_123_981 ();
 DECAPx4_ASAP7_75t_R FILLER_123_989 ();
 FILLER_ASAP7_75t_R FILLER_123_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_123_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1118 ();
 FILLER_ASAP7_75t_R FILLER_123_1127 ();
 FILLER_ASAP7_75t_R FILLER_123_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1138 ();
 FILLER_ASAP7_75t_R FILLER_123_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1151 ();
 FILLER_ASAP7_75t_R FILLER_123_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1172 ();
 FILLER_ASAP7_75t_R FILLER_123_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1186 ();
 FILLER_ASAP7_75t_R FILLER_123_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1220 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1231 ();
 FILLER_ASAP7_75t_R FILLER_123_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1247 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1255 ();
 FILLER_ASAP7_75t_R FILLER_123_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_124_954 ();
 DECAPx10_ASAP7_75t_R FILLER_124_976 ();
 DECAPx10_ASAP7_75t_R FILLER_124_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1037 ();
 FILLER_ASAP7_75t_R FILLER_124_1051 ();
 FILLER_ASAP7_75t_R FILLER_124_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1113 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1159 ();
 FILLER_ASAP7_75t_R FILLER_124_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_124_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1229 ();
 FILLER_ASAP7_75t_R FILLER_124_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_125_947 ();
 FILLER_ASAP7_75t_R FILLER_125_953 ();
 FILLER_ASAP7_75t_R FILLER_125_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_974 ();
 FILLER_ASAP7_75t_R FILLER_125_981 ();
 DECAPx6_ASAP7_75t_R FILLER_125_995 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1106 ();
 FILLER_ASAP7_75t_R FILLER_125_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_125_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1146 ();
 FILLER_ASAP7_75t_R FILLER_125_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1169 ();
 FILLER_ASAP7_75t_R FILLER_125_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1196 ();
 FILLER_ASAP7_75t_R FILLER_125_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1245 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1277 ();
 FILLER_ASAP7_75t_R FILLER_125_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_126_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_924 ();
 DECAPx2_ASAP7_75t_R FILLER_126_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_961 ();
 DECAPx1_ASAP7_75t_R FILLER_126_983 ();
 DECAPx4_ASAP7_75t_R FILLER_126_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1059 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1070 ();
 FILLER_ASAP7_75t_R FILLER_126_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1101 ();
 FILLER_ASAP7_75t_R FILLER_126_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_126_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1166 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1188 ();
 FILLER_ASAP7_75t_R FILLER_126_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1269 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1281 ();
 FILLER_ASAP7_75t_R FILLER_126_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_127_918 ();
 DECAPx10_ASAP7_75t_R FILLER_127_940 ();
 DECAPx2_ASAP7_75t_R FILLER_127_980 ();
 FILLER_ASAP7_75t_R FILLER_127_986 ();
 DECAPx4_ASAP7_75t_R FILLER_127_998 ();
 FILLER_ASAP7_75t_R FILLER_127_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1017 ();
 FILLER_ASAP7_75t_R FILLER_127_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1107 ();
 FILLER_ASAP7_75t_R FILLER_127_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1168 ();
 FILLER_ASAP7_75t_R FILLER_127_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1198 ();
 FILLER_ASAP7_75t_R FILLER_127_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_128_918 ();
 DECAPx2_ASAP7_75t_R FILLER_128_932 ();
 DECAPx10_ASAP7_75t_R FILLER_128_944 ();
 DECAPx10_ASAP7_75t_R FILLER_128_966 ();
 DECAPx4_ASAP7_75t_R FILLER_128_988 ();
 FILLER_ASAP7_75t_R FILLER_128_998 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1026 ();
 FILLER_ASAP7_75t_R FILLER_128_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_128_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_128_1105 ();
 FILLER_ASAP7_75t_R FILLER_128_1115 ();
 FILLER_ASAP7_75t_R FILLER_128_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1230 ();
 FILLER_ASAP7_75t_R FILLER_128_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1238 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1246 ();
 FILLER_ASAP7_75t_R FILLER_128_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_129_918 ();
 DECAPx1_ASAP7_75t_R FILLER_129_940 ();
 DECAPx4_ASAP7_75t_R FILLER_129_950 ();
 FILLER_ASAP7_75t_R FILLER_129_960 ();
 DECAPx6_ASAP7_75t_R FILLER_129_972 ();
 DECAPx2_ASAP7_75t_R FILLER_129_986 ();
 FILLER_ASAP7_75t_R FILLER_129_1010 ();
 FILLER_ASAP7_75t_R FILLER_129_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1051 ();
 FILLER_ASAP7_75t_R FILLER_129_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1118 ();
 FILLER_ASAP7_75t_R FILLER_129_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1131 ();
 FILLER_ASAP7_75t_R FILLER_129_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1147 ();
 FILLER_ASAP7_75t_R FILLER_129_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1184 ();
 FILLER_ASAP7_75t_R FILLER_129_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1219 ();
 FILLER_ASAP7_75t_R FILLER_129_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1261 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1279 ();
 FILLER_ASAP7_75t_R FILLER_130_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_920 ();
 DECAPx6_ASAP7_75t_R FILLER_130_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_944 ();
 DECAPx2_ASAP7_75t_R FILLER_130_951 ();
 FILLER_ASAP7_75t_R FILLER_130_957 ();
 DECAPx10_ASAP7_75t_R FILLER_130_969 ();
 DECAPx10_ASAP7_75t_R FILLER_130_997 ();
 FILLER_ASAP7_75t_R FILLER_130_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1095 ();
 FILLER_ASAP7_75t_R FILLER_130_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1199 ();
 FILLER_ASAP7_75t_R FILLER_130_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1213 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1220 ();
 FILLER_ASAP7_75t_R FILLER_130_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1247 ();
 FILLER_ASAP7_75t_R FILLER_130_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_131_918 ();
 DECAPx10_ASAP7_75t_R FILLER_131_940 ();
 DECAPx1_ASAP7_75t_R FILLER_131_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_966 ();
 DECAPx4_ASAP7_75t_R FILLER_131_974 ();
 FILLER_ASAP7_75t_R FILLER_131_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1121 ();
 FILLER_ASAP7_75t_R FILLER_131_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1167 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1193 ();
 FILLER_ASAP7_75t_R FILLER_131_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1226 ();
 FILLER_ASAP7_75t_R FILLER_131_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_132_918 ();
 DECAPx10_ASAP7_75t_R FILLER_132_932 ();
 DECAPx2_ASAP7_75t_R FILLER_132_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_960 ();
 DECAPx2_ASAP7_75t_R FILLER_132_994 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1082 ();
 FILLER_ASAP7_75t_R FILLER_132_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1097 ();
 FILLER_ASAP7_75t_R FILLER_132_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1185 ();
 FILLER_ASAP7_75t_R FILLER_132_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1216 ();
 FILLER_ASAP7_75t_R FILLER_132_1222 ();
 FILLER_ASAP7_75t_R FILLER_132_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1271 ();
 DECAPx1_ASAP7_75t_R FILLER_133_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_922 ();
 DECAPx4_ASAP7_75t_R FILLER_133_935 ();
 FILLER_ASAP7_75t_R FILLER_133_945 ();
 DECAPx4_ASAP7_75t_R FILLER_133_950 ();
 FILLER_ASAP7_75t_R FILLER_133_960 ();
 DECAPx1_ASAP7_75t_R FILLER_133_968 ();
 DECAPx4_ASAP7_75t_R FILLER_133_979 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1008 ();
 FILLER_ASAP7_75t_R FILLER_133_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1028 ();
 FILLER_ASAP7_75t_R FILLER_133_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1131 ();
 FILLER_ASAP7_75t_R FILLER_133_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1148 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1195 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1202 ();
 FILLER_ASAP7_75t_R FILLER_133_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1224 ();
 DECAPx6_ASAP7_75t_R FILLER_133_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_134_918 ();
 FILLER_ASAP7_75t_R FILLER_134_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_926 ();
 DECAPx10_ASAP7_75t_R FILLER_134_955 ();
 FILLER_ASAP7_75t_R FILLER_134_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1024 ();
 FILLER_ASAP7_75t_R FILLER_134_1035 ();
 FILLER_ASAP7_75t_R FILLER_134_1051 ();
 FILLER_ASAP7_75t_R FILLER_134_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1236 ();
 FILLER_ASAP7_75t_R FILLER_134_1242 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1265 ();
 FILLER_ASAP7_75t_R FILLER_134_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1281 ();
 FILLER_ASAP7_75t_R FILLER_134_1291 ();
 FILLER_ASAP7_75t_R FILLER_135_918 ();
 DECAPx4_ASAP7_75t_R FILLER_135_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_942 ();
 DECAPx10_ASAP7_75t_R FILLER_135_950 ();
 DECAPx6_ASAP7_75t_R FILLER_135_972 ();
 DECAPx2_ASAP7_75t_R FILLER_135_986 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1046 ();
 FILLER_ASAP7_75t_R FILLER_135_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1077 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1102 ();
 FILLER_ASAP7_75t_R FILLER_135_1133 ();
 FILLER_ASAP7_75t_R FILLER_135_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1188 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1277 ();
 FILLER_ASAP7_75t_R FILLER_135_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_136_918 ();
 FILLER_ASAP7_75t_R FILLER_136_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_934 ();
 DECAPx6_ASAP7_75t_R FILLER_136_940 ();
 DECAPx1_ASAP7_75t_R FILLER_136_954 ();
 DECAPx4_ASAP7_75t_R FILLER_136_964 ();
 DECAPx10_ASAP7_75t_R FILLER_136_980 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1002 ();
 FILLER_ASAP7_75t_R FILLER_136_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1121 ();
 FILLER_ASAP7_75t_R FILLER_136_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_136_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1185 ();
 FILLER_ASAP7_75t_R FILLER_136_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1225 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1260 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_137_918 ();
 DECAPx10_ASAP7_75t_R FILLER_137_943 ();
 DECAPx4_ASAP7_75t_R FILLER_137_965 ();
 FILLER_ASAP7_75t_R FILLER_137_975 ();
 DECAPx10_ASAP7_75t_R FILLER_137_987 ();
 FILLER_ASAP7_75t_R FILLER_137_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1128 ();
 FILLER_ASAP7_75t_R FILLER_137_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1203 ();
 FILLER_ASAP7_75t_R FILLER_137_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_137_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_138_918 ();
 DECAPx10_ASAP7_75t_R FILLER_138_940 ();
 DECAPx10_ASAP7_75t_R FILLER_138_962 ();
 DECAPx6_ASAP7_75t_R FILLER_138_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_998 ();
 FILLER_ASAP7_75t_R FILLER_138_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1041 ();
 FILLER_ASAP7_75t_R FILLER_138_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1054 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1108 ();
 FILLER_ASAP7_75t_R FILLER_138_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_138_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1236 ();
 FILLER_ASAP7_75t_R FILLER_138_1242 ();
 FILLER_ASAP7_75t_R FILLER_138_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_139_918 ();
 DECAPx10_ASAP7_75t_R FILLER_139_940 ();
 DECAPx10_ASAP7_75t_R FILLER_139_962 ();
 DECAPx4_ASAP7_75t_R FILLER_139_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_994 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1015 ();
 FILLER_ASAP7_75t_R FILLER_139_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1061 ();
 FILLER_ASAP7_75t_R FILLER_139_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1076 ();
 FILLER_ASAP7_75t_R FILLER_139_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1109 ();
 FILLER_ASAP7_75t_R FILLER_139_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1117 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1145 ();
 FILLER_ASAP7_75t_R FILLER_139_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_140_918 ();
 DECAPx6_ASAP7_75t_R FILLER_140_940 ();
 FILLER_ASAP7_75t_R FILLER_140_954 ();
 DECAPx10_ASAP7_75t_R FILLER_140_964 ();
 DECAPx10_ASAP7_75t_R FILLER_140_986 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1063 ();
 FILLER_ASAP7_75t_R FILLER_140_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1124 ();
 FILLER_ASAP7_75t_R FILLER_140_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1166 ();
 FILLER_ASAP7_75t_R FILLER_140_1188 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1196 ();
 FILLER_ASAP7_75t_R FILLER_140_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1235 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1246 ();
 FILLER_ASAP7_75t_R FILLER_140_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1292 ();
 FILLER_ASAP7_75t_R FILLER_141_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_920 ();
 DECAPx4_ASAP7_75t_R FILLER_141_943 ();
 FILLER_ASAP7_75t_R FILLER_141_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_955 ();
 FILLER_ASAP7_75t_R FILLER_141_962 ();
 DECAPx6_ASAP7_75t_R FILLER_141_976 ();
 DECAPx10_ASAP7_75t_R FILLER_141_998 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1111 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_141_1142 ();
 FILLER_ASAP7_75t_R FILLER_141_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1232 ();
 FILLER_ASAP7_75t_R FILLER_141_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1240 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1251 ();
 FILLER_ASAP7_75t_R FILLER_141_1261 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_918 ();
 DECAPx2_ASAP7_75t_R FILLER_142_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_946 ();
 DECAPx10_ASAP7_75t_R FILLER_142_953 ();
 DECAPx10_ASAP7_75t_R FILLER_142_975 ();
 DECAPx4_ASAP7_75t_R FILLER_142_997 ();
 FILLER_ASAP7_75t_R FILLER_142_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1028 ();
 FILLER_ASAP7_75t_R FILLER_142_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1082 ();
 FILLER_ASAP7_75t_R FILLER_142_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1144 ();
 FILLER_ASAP7_75t_R FILLER_142_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1232 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1281 ();
 FILLER_ASAP7_75t_R FILLER_142_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_143_918 ();
 DECAPx1_ASAP7_75t_R FILLER_143_945 ();
 DECAPx10_ASAP7_75t_R FILLER_143_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1102 ();
 FILLER_ASAP7_75t_R FILLER_143_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1131 ();
 FILLER_ASAP7_75t_R FILLER_143_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1175 ();
 FILLER_ASAP7_75t_R FILLER_143_1197 ();
 FILLER_ASAP7_75t_R FILLER_143_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1232 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1281 ();
 FILLER_ASAP7_75t_R FILLER_143_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_144_918 ();
 DECAPx6_ASAP7_75t_R FILLER_144_940 ();
 DECAPx1_ASAP7_75t_R FILLER_144_954 ();
 DECAPx6_ASAP7_75t_R FILLER_144_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_978 ();
 DECAPx6_ASAP7_75t_R FILLER_144_992 ();
 FILLER_ASAP7_75t_R FILLER_144_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1070 ();
 FILLER_ASAP7_75t_R FILLER_144_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1089 ();
 FILLER_ASAP7_75t_R FILLER_144_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1235 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1266 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_145_918 ();
 DECAPx6_ASAP7_75t_R FILLER_145_940 ();
 DECAPx6_ASAP7_75t_R FILLER_145_969 ();
 FILLER_ASAP7_75t_R FILLER_145_983 ();
 DECAPx10_ASAP7_75t_R FILLER_145_995 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1017 ();
 FILLER_ASAP7_75t_R FILLER_145_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1142 ();
 FILLER_ASAP7_75t_R FILLER_145_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1156 ();
 FILLER_ASAP7_75t_R FILLER_145_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_145_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1200 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1212 ();
 FILLER_ASAP7_75t_R FILLER_145_1222 ();
 FILLER_ASAP7_75t_R FILLER_145_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1229 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1255 ();
 FILLER_ASAP7_75t_R FILLER_145_1265 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_146_918 ();
 DECAPx10_ASAP7_75t_R FILLER_146_948 ();
 DECAPx2_ASAP7_75t_R FILLER_146_970 ();
 FILLER_ASAP7_75t_R FILLER_146_976 ();
 FILLER_ASAP7_75t_R FILLER_146_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_986 ();
 DECAPx10_ASAP7_75t_R FILLER_146_997 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1084 ();
 FILLER_ASAP7_75t_R FILLER_146_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_146_1103 ();
 FILLER_ASAP7_75t_R FILLER_146_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1150 ();
 FILLER_ASAP7_75t_R FILLER_146_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1201 ();
 FILLER_ASAP7_75t_R FILLER_146_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_147_918 ();
 DECAPx6_ASAP7_75t_R FILLER_147_940 ();
 DECAPx1_ASAP7_75t_R FILLER_147_954 ();
 DECAPx2_ASAP7_75t_R FILLER_147_970 ();
 FILLER_ASAP7_75t_R FILLER_147_976 ();
 DECAPx4_ASAP7_75t_R FILLER_147_994 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1057 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1130 ();
 FILLER_ASAP7_75t_R FILLER_147_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1189 ();
 FILLER_ASAP7_75t_R FILLER_147_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1232 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1280 ();
 FILLER_ASAP7_75t_R FILLER_147_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_148_948 ();
 DECAPx2_ASAP7_75t_R FILLER_148_960 ();
 FILLER_ASAP7_75t_R FILLER_148_978 ();
 DECAPx10_ASAP7_75t_R FILLER_148_988 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1064 ();
 FILLER_ASAP7_75t_R FILLER_148_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_148_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1198 ();
 FILLER_ASAP7_75t_R FILLER_148_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_149_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_928 ();
 DECAPx4_ASAP7_75t_R FILLER_149_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_953 ();
 DECAPx6_ASAP7_75t_R FILLER_149_960 ();
 DECAPx1_ASAP7_75t_R FILLER_149_988 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1008 ();
 FILLER_ASAP7_75t_R FILLER_149_1022 ();
 FILLER_ASAP7_75t_R FILLER_149_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1047 ();
 FILLER_ASAP7_75t_R FILLER_149_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1074 ();
 FILLER_ASAP7_75t_R FILLER_149_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1108 ();
 FILLER_ASAP7_75t_R FILLER_149_1136 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1180 ();
 FILLER_ASAP7_75t_R FILLER_149_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1198 ();
 FILLER_ASAP7_75t_R FILLER_149_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_149_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1252 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1259 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_150_918 ();
 DECAPx10_ASAP7_75t_R FILLER_150_940 ();
 DECAPx10_ASAP7_75t_R FILLER_150_962 ();
 DECAPx6_ASAP7_75t_R FILLER_150_984 ();
 DECAPx2_ASAP7_75t_R FILLER_150_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1051 ();
 FILLER_ASAP7_75t_R FILLER_150_1073 ();
 DECAPx4_ASAP7_75t_R FILLER_150_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1180 ();
 FILLER_ASAP7_75t_R FILLER_150_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1223 ();
 FILLER_ASAP7_75t_R FILLER_150_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_151_918 ();
 DECAPx6_ASAP7_75t_R FILLER_151_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_983 ();
 DECAPx4_ASAP7_75t_R FILLER_151_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1015 ();
 FILLER_ASAP7_75t_R FILLER_151_1025 ();
 FILLER_ASAP7_75t_R FILLER_151_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1061 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1097 ();
 FILLER_ASAP7_75t_R FILLER_151_1110 ();
 FILLER_ASAP7_75t_R FILLER_151_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_152_918 ();
 FILLER_ASAP7_75t_R FILLER_152_928 ();
 FILLER_ASAP7_75t_R FILLER_152_937 ();
 DECAPx6_ASAP7_75t_R FILLER_152_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_960 ();
 DECAPx10_ASAP7_75t_R FILLER_152_981 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1132 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1184 ();
 FILLER_ASAP7_75t_R FILLER_152_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1235 ();
 FILLER_ASAP7_75t_R FILLER_152_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1284 ();
 FILLER_ASAP7_75t_R FILLER_152_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_153_918 ();
 DECAPx2_ASAP7_75t_R FILLER_153_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_946 ();
 DECAPx10_ASAP7_75t_R FILLER_153_953 ();
 DECAPx10_ASAP7_75t_R FILLER_153_975 ();
 DECAPx2_ASAP7_75t_R FILLER_153_997 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_153_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1085 ();
 FILLER_ASAP7_75t_R FILLER_153_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_153_1153 ();
 FILLER_ASAP7_75t_R FILLER_153_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1277 ();
 FILLER_ASAP7_75t_R FILLER_153_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_154_918 ();
 FILLER_ASAP7_75t_R FILLER_154_924 ();
 FILLER_ASAP7_75t_R FILLER_154_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_940 ();
 FILLER_ASAP7_75t_R FILLER_154_944 ();
 DECAPx4_ASAP7_75t_R FILLER_154_969 ();
 FILLER_ASAP7_75t_R FILLER_154_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_981 ();
 DECAPx2_ASAP7_75t_R FILLER_154_988 ();
 FILLER_ASAP7_75t_R FILLER_154_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_996 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1059 ();
 FILLER_ASAP7_75t_R FILLER_154_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1112 ();
 FILLER_ASAP7_75t_R FILLER_154_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1155 ();
 FILLER_ASAP7_75t_R FILLER_154_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1210 ();
 FILLER_ASAP7_75t_R FILLER_154_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1232 ();
 FILLER_ASAP7_75t_R FILLER_154_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1240 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1281 ();
 FILLER_ASAP7_75t_R FILLER_154_1291 ();
 DECAPx4_ASAP7_75t_R FILLER_155_918 ();
 FILLER_ASAP7_75t_R FILLER_155_928 ();
 DECAPx2_ASAP7_75t_R FILLER_155_951 ();
 FILLER_ASAP7_75t_R FILLER_155_957 ();
 DECAPx10_ASAP7_75t_R FILLER_155_966 ();
 DECAPx2_ASAP7_75t_R FILLER_155_988 ();
 FILLER_ASAP7_75t_R FILLER_155_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_996 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1043 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1096 ();
 FILLER_ASAP7_75t_R FILLER_155_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1105 ();
 FILLER_ASAP7_75t_R FILLER_155_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1185 ();
 FILLER_ASAP7_75t_R FILLER_155_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1234 ();
 FILLER_ASAP7_75t_R FILLER_155_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_156_918 ();
 FILLER_ASAP7_75t_R FILLER_156_924 ();
 DECAPx10_ASAP7_75t_R FILLER_156_936 ();
 DECAPx10_ASAP7_75t_R FILLER_156_990 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1012 ();
 FILLER_ASAP7_75t_R FILLER_156_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1080 ();
 FILLER_ASAP7_75t_R FILLER_156_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1096 ();
 FILLER_ASAP7_75t_R FILLER_156_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_157_918 ();
 DECAPx10_ASAP7_75t_R FILLER_157_940 ();
 DECAPx2_ASAP7_75t_R FILLER_157_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_968 ();
 DECAPx10_ASAP7_75t_R FILLER_157_977 ();
 DECAPx10_ASAP7_75t_R FILLER_157_999 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1043 ();
 FILLER_ASAP7_75t_R FILLER_157_1049 ();
 FILLER_ASAP7_75t_R FILLER_157_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1096 ();
 FILLER_ASAP7_75t_R FILLER_157_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1189 ();
 FILLER_ASAP7_75t_R FILLER_157_1196 ();
 FILLER_ASAP7_75t_R FILLER_157_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1228 ();
 FILLER_ASAP7_75t_R FILLER_157_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_158_918 ();
 DECAPx2_ASAP7_75t_R FILLER_158_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_938 ();
 DECAPx10_ASAP7_75t_R FILLER_158_946 ();
 DECAPx10_ASAP7_75t_R FILLER_158_968 ();
 DECAPx4_ASAP7_75t_R FILLER_158_990 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_158_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1155 ();
 FILLER_ASAP7_75t_R FILLER_158_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1189 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1243 ();
 FILLER_ASAP7_75t_R FILLER_158_1270 ();
 DECAPx1_ASAP7_75t_R FILLER_159_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_938 ();
 DECAPx2_ASAP7_75t_R FILLER_159_945 ();
 DECAPx6_ASAP7_75t_R FILLER_159_963 ();
 DECAPx2_ASAP7_75t_R FILLER_159_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_983 ();
 DECAPx6_ASAP7_75t_R FILLER_159_990 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1017 ();
 FILLER_ASAP7_75t_R FILLER_159_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_159_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_159_1113 ();
 FILLER_ASAP7_75t_R FILLER_159_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1224 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1256 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1260 ();
 DECAPx6_ASAP7_75t_R FILLER_159_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_160_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_928 ();
 DECAPx6_ASAP7_75t_R FILLER_160_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_964 ();
 DECAPx1_ASAP7_75t_R FILLER_160_977 ();
 DECAPx10_ASAP7_75t_R FILLER_160_991 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1094 ();
 FILLER_ASAP7_75t_R FILLER_160_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1134 ();
 FILLER_ASAP7_75t_R FILLER_160_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1200 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1222 ();
 FILLER_ASAP7_75t_R FILLER_160_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1283 ();
 DECAPx4_ASAP7_75t_R FILLER_161_918 ();
 FILLER_ASAP7_75t_R FILLER_161_928 ();
 DECAPx10_ASAP7_75t_R FILLER_161_944 ();
 DECAPx10_ASAP7_75t_R FILLER_161_966 ();
 DECAPx10_ASAP7_75t_R FILLER_161_988 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_161_1083 ();
 FILLER_ASAP7_75t_R FILLER_161_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1095 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1118 ();
 FILLER_ASAP7_75t_R FILLER_161_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1231 ();
 FILLER_ASAP7_75t_R FILLER_161_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1267 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_162_918 ();
 DECAPx2_ASAP7_75t_R FILLER_162_940 ();
 DECAPx10_ASAP7_75t_R FILLER_162_956 ();
 DECAPx6_ASAP7_75t_R FILLER_162_978 ();
 FILLER_ASAP7_75t_R FILLER_162_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_994 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1093 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1119 ();
 FILLER_ASAP7_75t_R FILLER_162_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1234 ();
 FILLER_ASAP7_75t_R FILLER_162_1244 ();
 FILLER_ASAP7_75t_R FILLER_162_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1264 ();
 DECAPx4_ASAP7_75t_R FILLER_163_918 ();
 FILLER_ASAP7_75t_R FILLER_163_928 ();
 DECAPx10_ASAP7_75t_R FILLER_163_934 ();
 DECAPx4_ASAP7_75t_R FILLER_163_956 ();
 FILLER_ASAP7_75t_R FILLER_163_966 ();
 DECAPx10_ASAP7_75t_R FILLER_163_974 ();
 DECAPx10_ASAP7_75t_R FILLER_163_996 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1108 ();
 FILLER_ASAP7_75t_R FILLER_163_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1150 ();
 FILLER_ASAP7_75t_R FILLER_163_1157 ();
 FILLER_ASAP7_75t_R FILLER_163_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1285 ();
 FILLER_ASAP7_75t_R FILLER_163_1291 ();
 FILLER_ASAP7_75t_R FILLER_164_918 ();
 DECAPx6_ASAP7_75t_R FILLER_164_951 ();
 DECAPx1_ASAP7_75t_R FILLER_164_965 ();
 DECAPx2_ASAP7_75t_R FILLER_164_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_987 ();
 FILLER_ASAP7_75t_R FILLER_164_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1060 ();
 FILLER_ASAP7_75t_R FILLER_164_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1197 ();
 FILLER_ASAP7_75t_R FILLER_164_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1256 ();
 FILLER_ASAP7_75t_R FILLER_164_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_165_918 ();
 FILLER_ASAP7_75t_R FILLER_165_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_926 ();
 DECAPx1_ASAP7_75t_R FILLER_165_944 ();
 DECAPx10_ASAP7_75t_R FILLER_165_958 ();
 DECAPx10_ASAP7_75t_R FILLER_165_980 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1002 ();
 FILLER_ASAP7_75t_R FILLER_165_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1054 ();
 FILLER_ASAP7_75t_R FILLER_165_1068 ();
 FILLER_ASAP7_75t_R FILLER_165_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1100 ();
 FILLER_ASAP7_75t_R FILLER_165_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1169 ();
 FILLER_ASAP7_75t_R FILLER_165_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1210 ();
 FILLER_ASAP7_75t_R FILLER_165_1216 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1226 ();
 FILLER_ASAP7_75t_R FILLER_165_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_165_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_166_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_928 ();
 DECAPx6_ASAP7_75t_R FILLER_166_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_951 ();
 DECAPx10_ASAP7_75t_R FILLER_166_960 ();
 DECAPx4_ASAP7_75t_R FILLER_166_982 ();
 FILLER_ASAP7_75t_R FILLER_166_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_994 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1005 ();
 FILLER_ASAP7_75t_R FILLER_166_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1044 ();
 FILLER_ASAP7_75t_R FILLER_166_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1200 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1209 ();
 FILLER_ASAP7_75t_R FILLER_166_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1221 ();
 DECAPx6_ASAP7_75t_R FILLER_166_1228 ();
 FILLER_ASAP7_75t_R FILLER_166_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_167_918 ();
 DECAPx10_ASAP7_75t_R FILLER_167_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_962 ();
 DECAPx6_ASAP7_75t_R FILLER_167_982 ();
 FILLER_ASAP7_75t_R FILLER_167_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_998 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_168_918 ();
 DECAPx2_ASAP7_75t_R FILLER_168_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_940 ();
 DECAPx6_ASAP7_75t_R FILLER_168_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_961 ();
 DECAPx4_ASAP7_75t_R FILLER_168_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_999 ();
 FILLER_ASAP7_75t_R FILLER_168_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1176 ();
 FILLER_ASAP7_75t_R FILLER_168_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1230 ();
 FILLER_ASAP7_75t_R FILLER_168_1252 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1281 ();
 FILLER_ASAP7_75t_R FILLER_168_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_169_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_924 ();
 DECAPx2_ASAP7_75t_R FILLER_169_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_970 ();
 DECAPx10_ASAP7_75t_R FILLER_169_978 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1145 ();
 FILLER_ASAP7_75t_R FILLER_169_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1153 ();
 FILLER_ASAP7_75t_R FILLER_169_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1188 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1229 ();
 FILLER_ASAP7_75t_R FILLER_169_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_170_918 ();
 FILLER_ASAP7_75t_R FILLER_170_932 ();
 DECAPx2_ASAP7_75t_R FILLER_170_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_947 ();
 DECAPx4_ASAP7_75t_R FILLER_170_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_971 ();
 FILLER_ASAP7_75t_R FILLER_170_1003 ();
 FILLER_ASAP7_75t_R FILLER_170_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1030 ();
 FILLER_ASAP7_75t_R FILLER_170_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1070 ();
 FILLER_ASAP7_75t_R FILLER_170_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1165 ();
 FILLER_ASAP7_75t_R FILLER_170_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1253 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1281 ();
 FILLER_ASAP7_75t_R FILLER_170_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_918 ();
 DECAPx4_ASAP7_75t_R FILLER_171_929 ();
 DECAPx1_ASAP7_75t_R FILLER_171_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_982 ();
 DECAPx4_ASAP7_75t_R FILLER_171_993 ();
 FILLER_ASAP7_75t_R FILLER_171_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1162 ();
 FILLER_ASAP7_75t_R FILLER_171_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1174 ();
 FILLER_ASAP7_75t_R FILLER_171_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1218 ();
 FILLER_ASAP7_75t_R FILLER_171_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1289 ();
 DECAPx1_ASAP7_75t_R FILLER_172_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_922 ();
 FILLER_ASAP7_75t_R FILLER_172_931 ();
 FILLER_ASAP7_75t_R FILLER_172_943 ();
 FILLER_ASAP7_75t_R FILLER_172_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1040 ();
 FILLER_ASAP7_75t_R FILLER_172_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1100 ();
 FILLER_ASAP7_75t_R FILLER_172_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1141 ();
 FILLER_ASAP7_75t_R FILLER_172_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1167 ();
 FILLER_ASAP7_75t_R FILLER_172_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1175 ();
 FILLER_ASAP7_75t_R FILLER_172_1182 ();
 FILLER_ASAP7_75t_R FILLER_172_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1203 ();
 FILLER_ASAP7_75t_R FILLER_172_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1246 ();
 DECAPx4_ASAP7_75t_R FILLER_172_1253 ();
 FILLER_ASAP7_75t_R FILLER_172_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_173_918 ();
 DECAPx2_ASAP7_75t_R FILLER_173_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_938 ();
 DECAPx2_ASAP7_75t_R FILLER_173_975 ();
 FILLER_ASAP7_75t_R FILLER_173_981 ();
 DECAPx1_ASAP7_75t_R FILLER_173_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1011 ();
 FILLER_ASAP7_75t_R FILLER_173_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1072 ();
 FILLER_ASAP7_75t_R FILLER_173_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1201 ();
 FILLER_ASAP7_75t_R FILLER_173_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_173_1254 ();
 FILLER_ASAP7_75t_R FILLER_173_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1274 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_174_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_922 ();
 DECAPx2_ASAP7_75t_R FILLER_174_944 ();
 FILLER_ASAP7_75t_R FILLER_174_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_952 ();
 DECAPx10_ASAP7_75t_R FILLER_174_968 ();
 FILLER_ASAP7_75t_R FILLER_174_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_992 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1024 ();
 FILLER_ASAP7_75t_R FILLER_174_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1115 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1220 ();
 FILLER_ASAP7_75t_R FILLER_174_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1232 ();
 FILLER_ASAP7_75t_R FILLER_174_1254 ();
 FILLER_ASAP7_75t_R FILLER_174_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_175_918 ();
 FILLER_ASAP7_75t_R FILLER_175_928 ();
 DECAPx10_ASAP7_75t_R FILLER_175_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_964 ();
 DECAPx6_ASAP7_75t_R FILLER_175_968 ();
 DECAPx1_ASAP7_75t_R FILLER_175_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_986 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1026 ();
 FILLER_ASAP7_75t_R FILLER_175_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1070 ();
 FILLER_ASAP7_75t_R FILLER_175_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1263 ();
 FILLER_ASAP7_75t_R FILLER_175_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_176_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_940 ();
 FILLER_ASAP7_75t_R FILLER_176_958 ();
 DECAPx6_ASAP7_75t_R FILLER_176_974 ();
 FILLER_ASAP7_75t_R FILLER_176_988 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1012 ();
 FILLER_ASAP7_75t_R FILLER_176_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1044 ();
 FILLER_ASAP7_75t_R FILLER_176_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1245 ();
 FILLER_ASAP7_75t_R FILLER_176_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_177_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_991 ();
 FILLER_ASAP7_75t_R FILLER_177_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1041 ();
 FILLER_ASAP7_75t_R FILLER_177_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1167 ();
 FILLER_ASAP7_75t_R FILLER_177_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1192 ();
 FILLER_ASAP7_75t_R FILLER_177_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1240 ();
 FILLER_ASAP7_75t_R FILLER_177_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_178_918 ();
 FILLER_ASAP7_75t_R FILLER_178_924 ();
 DECAPx4_ASAP7_75t_R FILLER_178_947 ();
 FILLER_ASAP7_75t_R FILLER_178_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_959 ();
 DECAPx4_ASAP7_75t_R FILLER_178_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_985 ();
 DECAPx6_ASAP7_75t_R FILLER_178_998 ();
 FILLER_ASAP7_75t_R FILLER_178_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1039 ();
 FILLER_ASAP7_75t_R FILLER_178_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1072 ();
 FILLER_ASAP7_75t_R FILLER_178_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1115 ();
 FILLER_ASAP7_75t_R FILLER_178_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1197 ();
 FILLER_ASAP7_75t_R FILLER_178_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1268 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1276 ();
 FILLER_ASAP7_75t_R FILLER_178_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_179_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_942 ();
 DECAPx2_ASAP7_75t_R FILLER_179_951 ();
 DECAPx10_ASAP7_75t_R FILLER_179_967 ();
 DECAPx6_ASAP7_75t_R FILLER_179_989 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1017 ();
 FILLER_ASAP7_75t_R FILLER_179_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1046 ();
 FILLER_ASAP7_75t_R FILLER_179_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1232 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1263 ();
 DECAPx4_ASAP7_75t_R FILLER_179_1280 ();
 FILLER_ASAP7_75t_R FILLER_179_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_180_918 ();
 DECAPx10_ASAP7_75t_R FILLER_180_940 ();
 DECAPx4_ASAP7_75t_R FILLER_180_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_972 ();
 DECAPx2_ASAP7_75t_R FILLER_180_989 ();
 FILLER_ASAP7_75t_R FILLER_180_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_997 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1016 ();
 FILLER_ASAP7_75t_R FILLER_180_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1068 ();
 FILLER_ASAP7_75t_R FILLER_180_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1263 ();
 FILLER_ASAP7_75t_R FILLER_180_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_181_918 ();
 DECAPx4_ASAP7_75t_R FILLER_181_940 ();
 FILLER_ASAP7_75t_R FILLER_181_976 ();
 DECAPx1_ASAP7_75t_R FILLER_181_999 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1110 ();
 FILLER_ASAP7_75t_R FILLER_181_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1159 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_182_918 ();
 DECAPx1_ASAP7_75t_R FILLER_182_940 ();
 FILLER_ASAP7_75t_R FILLER_182_954 ();
 DECAPx1_ASAP7_75t_R FILLER_182_976 ();
 DECAPx4_ASAP7_75t_R FILLER_182_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1040 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1176 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1228 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1265 ();
 FILLER_ASAP7_75t_R FILLER_182_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_183_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_922 ();
 FILLER_ASAP7_75t_R FILLER_183_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_935 ();
 FILLER_ASAP7_75t_R FILLER_183_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_959 ();
 DECAPx4_ASAP7_75t_R FILLER_183_963 ();
 FILLER_ASAP7_75t_R FILLER_183_973 ();
 FILLER_ASAP7_75t_R FILLER_183_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_984 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1056 ();
 FILLER_ASAP7_75t_R FILLER_183_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1134 ();
 FILLER_ASAP7_75t_R FILLER_183_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1151 ();
 FILLER_ASAP7_75t_R FILLER_183_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1173 ();
 FILLER_ASAP7_75t_R FILLER_183_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_184_918 ();
 FILLER_ASAP7_75t_R FILLER_184_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_942 ();
 DECAPx1_ASAP7_75t_R FILLER_184_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_953 ();
 DECAPx4_ASAP7_75t_R FILLER_184_981 ();
 FILLER_ASAP7_75t_R FILLER_184_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_993 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1073 ();
 FILLER_ASAP7_75t_R FILLER_184_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_185_918 ();
 FILLER_ASAP7_75t_R FILLER_185_952 ();
 DECAPx4_ASAP7_75t_R FILLER_185_966 ();
 DECAPx4_ASAP7_75t_R FILLER_185_988 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1057 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1113 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1249 ();
 FILLER_ASAP7_75t_R FILLER_185_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1274 ();
 DECAPx6_ASAP7_75t_R FILLER_186_918 ();
 DECAPx1_ASAP7_75t_R FILLER_186_932 ();
 DECAPx10_ASAP7_75t_R FILLER_186_946 ();
 DECAPx6_ASAP7_75t_R FILLER_186_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_982 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1004 ();
 FILLER_ASAP7_75t_R FILLER_186_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1028 ();
 FILLER_ASAP7_75t_R FILLER_186_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_186_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1077 ();
 FILLER_ASAP7_75t_R FILLER_186_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1107 ();
 FILLER_ASAP7_75t_R FILLER_186_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1142 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1149 ();
 FILLER_ASAP7_75t_R FILLER_186_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1198 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_186_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_187_918 ();
 DECAPx1_ASAP7_75t_R FILLER_187_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_957 ();
 DECAPx10_ASAP7_75t_R FILLER_187_980 ();
 DECAPx1_ASAP7_75t_R FILLER_187_1002 ();
 FILLER_ASAP7_75t_R FILLER_187_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1048 ();
 FILLER_ASAP7_75t_R FILLER_187_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1080 ();
 FILLER_ASAP7_75t_R FILLER_187_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1126 ();
 FILLER_ASAP7_75t_R FILLER_187_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1192 ();
 FILLER_ASAP7_75t_R FILLER_187_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1200 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1208 ();
 FILLER_ASAP7_75t_R FILLER_187_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1259 ();
 FILLER_ASAP7_75t_R FILLER_187_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_188_918 ();
 DECAPx1_ASAP7_75t_R FILLER_188_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_936 ();
 DECAPx1_ASAP7_75t_R FILLER_188_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_948 ();
 DECAPx2_ASAP7_75t_R FILLER_188_962 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1045 ();
 FILLER_ASAP7_75t_R FILLER_188_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1090 ();
 FILLER_ASAP7_75t_R FILLER_188_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1199 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1230 ();
 FILLER_ASAP7_75t_R FILLER_188_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_188_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_188_1277 ();
 FILLER_ASAP7_75t_R FILLER_188_1291 ();
 DECAPx4_ASAP7_75t_R FILLER_189_918 ();
 FILLER_ASAP7_75t_R FILLER_189_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_951 ();
 DECAPx1_ASAP7_75t_R FILLER_189_967 ();
 DECAPx2_ASAP7_75t_R FILLER_189_977 ();
 FILLER_ASAP7_75t_R FILLER_189_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_985 ();
 DECAPx4_ASAP7_75t_R FILLER_189_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1124 ();
 FILLER_ASAP7_75t_R FILLER_189_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1142 ();
 FILLER_ASAP7_75t_R FILLER_189_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1246 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1278 ();
 DECAPx4_ASAP7_75t_R FILLER_190_918 ();
 FILLER_ASAP7_75t_R FILLER_190_928 ();
 FILLER_ASAP7_75t_R FILLER_190_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_992 ();
 DECAPx4_ASAP7_75t_R FILLER_190_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_190_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1096 ();
 FILLER_ASAP7_75t_R FILLER_190_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1171 ();
 FILLER_ASAP7_75t_R FILLER_190_1193 ();
 FILLER_ASAP7_75t_R FILLER_190_1202 ();
 FILLER_ASAP7_75t_R FILLER_190_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_191_918 ();
 DECAPx4_ASAP7_75t_R FILLER_191_940 ();
 FILLER_ASAP7_75t_R FILLER_191_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_952 ();
 DECAPx10_ASAP7_75t_R FILLER_191_956 ();
 DECAPx10_ASAP7_75t_R FILLER_191_978 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_191_1052 ();
 FILLER_ASAP7_75t_R FILLER_191_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1212 ();
 FILLER_ASAP7_75t_R FILLER_191_1226 ();
 FILLER_ASAP7_75t_R FILLER_191_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1292 ();
 FILLER_ASAP7_75t_R FILLER_192_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_942 ();
 FILLER_ASAP7_75t_R FILLER_192_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_958 ();
 DECAPx4_ASAP7_75t_R FILLER_192_962 ();
 FILLER_ASAP7_75t_R FILLER_192_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_981 ();
 FILLER_ASAP7_75t_R FILLER_192_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_990 ();
 DECAPx10_ASAP7_75t_R FILLER_192_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1048 ();
 FILLER_ASAP7_75t_R FILLER_192_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_192_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_192_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1208 ();
 FILLER_ASAP7_75t_R FILLER_192_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1230 ();
 FILLER_ASAP7_75t_R FILLER_192_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_193_918 ();
 FILLER_ASAP7_75t_R FILLER_193_928 ();
 FILLER_ASAP7_75t_R FILLER_193_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_939 ();
 DECAPx4_ASAP7_75t_R FILLER_193_950 ();
 DECAPx2_ASAP7_75t_R FILLER_193_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_987 ();
 DECAPx2_ASAP7_75t_R FILLER_193_994 ();
 FILLER_ASAP7_75t_R FILLER_193_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_193_1034 ();
 FILLER_ASAP7_75t_R FILLER_193_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1072 ();
 FILLER_ASAP7_75t_R FILLER_193_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1241 ();
 FILLER_ASAP7_75t_R FILLER_193_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_194_918 ();
 DECAPx1_ASAP7_75t_R FILLER_194_944 ();
 FILLER_ASAP7_75t_R FILLER_194_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1096 ();
 FILLER_ASAP7_75t_R FILLER_194_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1108 ();
 FILLER_ASAP7_75t_R FILLER_194_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1156 ();
 FILLER_ASAP7_75t_R FILLER_194_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1164 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1193 ();
 FILLER_ASAP7_75t_R FILLER_194_1199 ();
 FILLER_ASAP7_75t_R FILLER_194_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1283 ();
 DECAPx6_ASAP7_75t_R FILLER_195_918 ();
 DECAPx2_ASAP7_75t_R FILLER_195_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_938 ();
 DECAPx1_ASAP7_75t_R FILLER_195_951 ();
 DECAPx6_ASAP7_75t_R FILLER_195_967 ();
 DECAPx2_ASAP7_75t_R FILLER_195_981 ();
 DECAPx2_ASAP7_75t_R FILLER_195_994 ();
 FILLER_ASAP7_75t_R FILLER_195_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1009 ();
 FILLER_ASAP7_75t_R FILLER_195_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1064 ();
 FILLER_ASAP7_75t_R FILLER_195_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1285 ();
 FILLER_ASAP7_75t_R FILLER_195_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_196_918 ();
 FILLER_ASAP7_75t_R FILLER_196_953 ();
 DECAPx2_ASAP7_75t_R FILLER_196_965 ();
 FILLER_ASAP7_75t_R FILLER_196_971 ();
 DECAPx10_ASAP7_75t_R FILLER_196_976 ();
 DECAPx4_ASAP7_75t_R FILLER_196_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1040 ();
 FILLER_ASAP7_75t_R FILLER_196_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1066 ();
 FILLER_ASAP7_75t_R FILLER_196_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1095 ();
 FILLER_ASAP7_75t_R FILLER_196_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1180 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1209 ();
 FILLER_ASAP7_75t_R FILLER_196_1219 ();
 FILLER_ASAP7_75t_R FILLER_196_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_197_918 ();
 DECAPx10_ASAP7_75t_R FILLER_197_940 ();
 DECAPx4_ASAP7_75t_R FILLER_197_965 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1023 ();
 FILLER_ASAP7_75t_R FILLER_197_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1038 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1098 ();
 FILLER_ASAP7_75t_R FILLER_197_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1197 ();
 FILLER_ASAP7_75t_R FILLER_197_1211 ();
 FILLER_ASAP7_75t_R FILLER_197_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1235 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_198_918 ();
 DECAPx2_ASAP7_75t_R FILLER_198_940 ();
 FILLER_ASAP7_75t_R FILLER_198_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_948 ();
 FILLER_ASAP7_75t_R FILLER_198_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_968 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1065 ();
 FILLER_ASAP7_75t_R FILLER_198_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1078 ();
 FILLER_ASAP7_75t_R FILLER_198_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1111 ();
 FILLER_ASAP7_75t_R FILLER_198_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1214 ();
 FILLER_ASAP7_75t_R FILLER_198_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1231 ();
 FILLER_ASAP7_75t_R FILLER_198_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1268 ();
 FILLER_ASAP7_75t_R FILLER_198_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_199_918 ();
 DECAPx1_ASAP7_75t_R FILLER_199_932 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1051 ();
 FILLER_ASAP7_75t_R FILLER_199_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1066 ();
 FILLER_ASAP7_75t_R FILLER_199_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1106 ();
 FILLER_ASAP7_75t_R FILLER_199_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1118 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_200_918 ();
 FILLER_ASAP7_75t_R FILLER_200_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_933 ();
 DECAPx4_ASAP7_75t_R FILLER_200_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_965 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1002 ();
 FILLER_ASAP7_75t_R FILLER_200_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1025 ();
 FILLER_ASAP7_75t_R FILLER_200_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1168 ();
 FILLER_ASAP7_75t_R FILLER_200_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_201_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_932 ();
 DECAPx2_ASAP7_75t_R FILLER_201_945 ();
 FILLER_ASAP7_75t_R FILLER_201_951 ();
 FILLER_ASAP7_75t_R FILLER_201_963 ();
 DECAPx10_ASAP7_75t_R FILLER_201_968 ();
 DECAPx2_ASAP7_75t_R FILLER_201_990 ();
 FILLER_ASAP7_75t_R FILLER_201_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1028 ();
 FILLER_ASAP7_75t_R FILLER_201_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1095 ();
 FILLER_ASAP7_75t_R FILLER_201_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1111 ();
 FILLER_ASAP7_75t_R FILLER_201_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1131 ();
 FILLER_ASAP7_75t_R FILLER_201_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1149 ();
 FILLER_ASAP7_75t_R FILLER_201_1166 ();
 FILLER_ASAP7_75t_R FILLER_201_1175 ();
 FILLER_ASAP7_75t_R FILLER_201_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1284 ();
 FILLER_ASAP7_75t_R FILLER_201_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_202_918 ();
 DECAPx1_ASAP7_75t_R FILLER_202_932 ();
 FILLER_ASAP7_75t_R FILLER_202_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1062 ();
 FILLER_ASAP7_75t_R FILLER_202_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1117 ();
 FILLER_ASAP7_75t_R FILLER_202_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_202_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_203_918 ();
 DECAPx4_ASAP7_75t_R FILLER_203_953 ();
 DECAPx4_ASAP7_75t_R FILLER_203_973 ();
 FILLER_ASAP7_75t_R FILLER_203_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_985 ();
 DECAPx6_ASAP7_75t_R FILLER_203_992 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1010 ();
 FILLER_ASAP7_75t_R FILLER_203_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1058 ();
 FILLER_ASAP7_75t_R FILLER_203_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_203_1109 ();
 FILLER_ASAP7_75t_R FILLER_203_1140 ();
 FILLER_ASAP7_75t_R FILLER_203_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1190 ();
 FILLER_ASAP7_75t_R FILLER_203_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1241 ();
 DECAPx6_ASAP7_75t_R FILLER_203_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_204_918 ();
 DECAPx2_ASAP7_75t_R FILLER_204_940 ();
 FILLER_ASAP7_75t_R FILLER_204_946 ();
 DECAPx2_ASAP7_75t_R FILLER_204_953 ();
 DECAPx2_ASAP7_75t_R FILLER_204_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_986 ();
 DECAPx4_ASAP7_75t_R FILLER_204_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1135 ();
 FILLER_ASAP7_75t_R FILLER_204_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1158 ();
 FILLER_ASAP7_75t_R FILLER_204_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1203 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_205_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_932 ();
 DECAPx1_ASAP7_75t_R FILLER_205_940 ();
 DECAPx1_ASAP7_75t_R FILLER_205_954 ();
 DECAPx6_ASAP7_75t_R FILLER_205_964 ();
 FILLER_ASAP7_75t_R FILLER_205_978 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1165 ();
 FILLER_ASAP7_75t_R FILLER_205_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1213 ();
 DECAPx1_ASAP7_75t_R FILLER_205_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1276 ();
 FILLER_ASAP7_75t_R FILLER_205_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1292 ();
 FILLER_ASAP7_75t_R FILLER_206_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_930 ();
 FILLER_ASAP7_75t_R FILLER_206_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_954 ();
 DECAPx2_ASAP7_75t_R FILLER_206_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_994 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1083 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1105 ();
 FILLER_ASAP7_75t_R FILLER_206_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_207_918 ();
 FILLER_ASAP7_75t_R FILLER_207_932 ();
 DECAPx2_ASAP7_75t_R FILLER_207_948 ();
 FILLER_ASAP7_75t_R FILLER_207_954 ();
 DECAPx2_ASAP7_75t_R FILLER_207_978 ();
 FILLER_ASAP7_75t_R FILLER_207_984 ();
 DECAPx4_ASAP7_75t_R FILLER_207_996 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1023 ();
 FILLER_ASAP7_75t_R FILLER_207_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1031 ();
 FILLER_ASAP7_75t_R FILLER_207_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1066 ();
 FILLER_ASAP7_75t_R FILLER_207_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1104 ();
 FILLER_ASAP7_75t_R FILLER_207_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1144 ();
 FILLER_ASAP7_75t_R FILLER_207_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1194 ();
 FILLER_ASAP7_75t_R FILLER_207_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1210 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_207_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_207_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_208_918 ();
 DECAPx10_ASAP7_75t_R FILLER_208_940 ();
 DECAPx4_ASAP7_75t_R FILLER_208_962 ();
 DECAPx6_ASAP7_75t_R FILLER_208_975 ();
 DECAPx1_ASAP7_75t_R FILLER_208_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1006 ();
 FILLER_ASAP7_75t_R FILLER_208_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1037 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1069 ();
 FILLER_ASAP7_75t_R FILLER_208_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1078 ();
 FILLER_ASAP7_75t_R FILLER_208_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_208_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1191 ();
 FILLER_ASAP7_75t_R FILLER_208_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1203 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1235 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_209_918 ();
 DECAPx10_ASAP7_75t_R FILLER_209_928 ();
 FILLER_ASAP7_75t_R FILLER_209_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_952 ();
 FILLER_ASAP7_75t_R FILLER_209_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_976 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1043 ();
 FILLER_ASAP7_75t_R FILLER_209_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1077 ();
 FILLER_ASAP7_75t_R FILLER_209_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_209_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_210_918 ();
 DECAPx1_ASAP7_75t_R FILLER_210_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_949 ();
 DECAPx2_ASAP7_75t_R FILLER_210_957 ();
 DECAPx1_ASAP7_75t_R FILLER_210_982 ();
 DECAPx4_ASAP7_75t_R FILLER_210_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1057 ();
 FILLER_ASAP7_75t_R FILLER_210_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1090 ();
 FILLER_ASAP7_75t_R FILLER_210_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1156 ();
 FILLER_ASAP7_75t_R FILLER_210_1162 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1212 ();
 FILLER_ASAP7_75t_R FILLER_210_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_210_1242 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_211_918 ();
 FILLER_ASAP7_75t_R FILLER_211_962 ();
 DECAPx10_ASAP7_75t_R FILLER_211_984 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1006 ();
 FILLER_ASAP7_75t_R FILLER_211_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_211_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1143 ();
 FILLER_ASAP7_75t_R FILLER_211_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_1166 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_211_1204 ();
 FILLER_ASAP7_75t_R FILLER_211_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_212_918 ();
 FILLER_ASAP7_75t_R FILLER_212_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_960 ();
 DECAPx6_ASAP7_75t_R FILLER_212_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_994 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_212_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1052 ();
 FILLER_ASAP7_75t_R FILLER_212_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1116 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1152 ();
 FILLER_ASAP7_75t_R FILLER_212_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1219 ();
 FILLER_ASAP7_75t_R FILLER_212_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1276 ();
 FILLER_ASAP7_75t_R FILLER_212_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_213_918 ();
 DECAPx2_ASAP7_75t_R FILLER_213_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_946 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1018 ();
 FILLER_ASAP7_75t_R FILLER_213_1028 ();
 FILLER_ASAP7_75t_R FILLER_213_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1081 ();
 FILLER_ASAP7_75t_R FILLER_213_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1167 ();
 FILLER_ASAP7_75t_R FILLER_213_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1197 ();
 FILLER_ASAP7_75t_R FILLER_213_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1205 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1216 ();
 FILLER_ASAP7_75t_R FILLER_213_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1228 ();
 FILLER_ASAP7_75t_R FILLER_213_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_214_918 ();
 DECAPx1_ASAP7_75t_R FILLER_214_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_936 ();
 DECAPx10_ASAP7_75t_R FILLER_214_989 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_214_1100 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1138 ();
 FILLER_ASAP7_75t_R FILLER_214_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_215_918 ();
 DECAPx2_ASAP7_75t_R FILLER_215_940 ();
 FILLER_ASAP7_75t_R FILLER_215_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_948 ();
 DECAPx1_ASAP7_75t_R FILLER_215_985 ();
 FILLER_ASAP7_75t_R FILLER_215_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_994 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1031 ();
 FILLER_ASAP7_75t_R FILLER_215_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_215_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_215_1161 ();
 FILLER_ASAP7_75t_R FILLER_215_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1269 ();
 FILLER_ASAP7_75t_R FILLER_215_1291 ();
 DECAPx4_ASAP7_75t_R FILLER_216_918 ();
 FILLER_ASAP7_75t_R FILLER_216_928 ();
 DECAPx2_ASAP7_75t_R FILLER_216_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_972 ();
 DECAPx1_ASAP7_75t_R FILLER_216_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1062 ();
 FILLER_ASAP7_75t_R FILLER_216_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_216_1172 ();
 FILLER_ASAP7_75t_R FILLER_216_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1202 ();
 FILLER_ASAP7_75t_R FILLER_216_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_217_918 ();
 FILLER_ASAP7_75t_R FILLER_217_932 ();
 DECAPx6_ASAP7_75t_R FILLER_217_968 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1099 ();
 FILLER_ASAP7_75t_R FILLER_217_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_218_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_924 ();
 DECAPx4_ASAP7_75t_R FILLER_218_939 ();
 FILLER_ASAP7_75t_R FILLER_218_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_951 ();
 DECAPx2_ASAP7_75t_R FILLER_218_970 ();
 DECAPx4_ASAP7_75t_R FILLER_218_988 ();
 FILLER_ASAP7_75t_R FILLER_218_998 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1066 ();
 FILLER_ASAP7_75t_R FILLER_218_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1168 ();
 FILLER_ASAP7_75t_R FILLER_218_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_218_1184 ();
 FILLER_ASAP7_75t_R FILLER_218_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_218_1213 ();
 FILLER_ASAP7_75t_R FILLER_218_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_219_918 ();
 DECAPx2_ASAP7_75t_R FILLER_219_940 ();
 FILLER_ASAP7_75t_R FILLER_219_958 ();
 DECAPx1_ASAP7_75t_R FILLER_219_981 ();
 DECAPx10_ASAP7_75t_R FILLER_219_988 ();
 DECAPx4_ASAP7_75t_R FILLER_219_1010 ();
 FILLER_ASAP7_75t_R FILLER_219_1020 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1176 ();
 FILLER_ASAP7_75t_R FILLER_219_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1243 ();
 DECAPx6_ASAP7_75t_R FILLER_219_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_219_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_220_918 ();
 FILLER_ASAP7_75t_R FILLER_220_959 ();
 DECAPx10_ASAP7_75t_R FILLER_220_994 ();
 FILLER_ASAP7_75t_R FILLER_220_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1065 ();
 FILLER_ASAP7_75t_R FILLER_220_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1134 ();
 FILLER_ASAP7_75t_R FILLER_220_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1174 ();
 FILLER_ASAP7_75t_R FILLER_220_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_220_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_221_918 ();
 DECAPx6_ASAP7_75t_R FILLER_221_940 ();
 FILLER_ASAP7_75t_R FILLER_221_954 ();
 DECAPx10_ASAP7_75t_R FILLER_221_968 ();
 DECAPx6_ASAP7_75t_R FILLER_221_990 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1015 ();
 FILLER_ASAP7_75t_R FILLER_221_1023 ();
 FILLER_ASAP7_75t_R FILLER_221_1042 ();
 FILLER_ASAP7_75t_R FILLER_221_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1067 ();
 FILLER_ASAP7_75t_R FILLER_221_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_221_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_222_918 ();
 DECAPx4_ASAP7_75t_R FILLER_222_940 ();
 FILLER_ASAP7_75t_R FILLER_222_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1024 ();
 FILLER_ASAP7_75t_R FILLER_222_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1082 ();
 FILLER_ASAP7_75t_R FILLER_222_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1133 ();
 FILLER_ASAP7_75t_R FILLER_222_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_222_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1269 ();
 FILLER_ASAP7_75t_R FILLER_222_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_223_918 ();
 DECAPx2_ASAP7_75t_R FILLER_223_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_950 ();
 DECAPx6_ASAP7_75t_R FILLER_223_954 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1004 ();
 DECAPx4_ASAP7_75t_R FILLER_223_1025 ();
 FILLER_ASAP7_75t_R FILLER_223_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_224_918 ();
 DECAPx10_ASAP7_75t_R FILLER_224_981 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1003 ();
 FILLER_ASAP7_75t_R FILLER_224_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1011 ();
 FILLER_ASAP7_75t_R FILLER_224_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_224_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_224_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1166 ();
 FILLER_ASAP7_75t_R FILLER_224_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1269 ();
 FILLER_ASAP7_75t_R FILLER_224_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_225_918 ();
 FILLER_ASAP7_75t_R FILLER_225_932 ();
 DECAPx6_ASAP7_75t_R FILLER_225_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_954 ();
 DECAPx2_ASAP7_75t_R FILLER_225_970 ();
 FILLER_ASAP7_75t_R FILLER_225_976 ();
 DECAPx1_ASAP7_75t_R FILLER_225_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_994 ();
 DECAPx10_ASAP7_75t_R FILLER_225_998 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_225_1072 ();
 FILLER_ASAP7_75t_R FILLER_225_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1190 ();
 FILLER_ASAP7_75t_R FILLER_225_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_226_918 ();
 FILLER_ASAP7_75t_R FILLER_226_928 ();
 DECAPx2_ASAP7_75t_R FILLER_226_951 ();
 DECAPx1_ASAP7_75t_R FILLER_226_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_982 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_226_1112 ();
 FILLER_ASAP7_75t_R FILLER_226_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_226_1194 ();
 FILLER_ASAP7_75t_R FILLER_226_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_226_1212 ();
 FILLER_ASAP7_75t_R FILLER_226_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_227_918 ();
 DECAPx2_ASAP7_75t_R FILLER_227_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_946 ();
 FILLER_ASAP7_75t_R FILLER_227_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_955 ();
 DECAPx2_ASAP7_75t_R FILLER_227_966 ();
 FILLER_ASAP7_75t_R FILLER_227_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_974 ();
 FILLER_ASAP7_75t_R FILLER_227_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1013 ();
 FILLER_ASAP7_75t_R FILLER_227_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1026 ();
 FILLER_ASAP7_75t_R FILLER_227_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_227_1049 ();
 FILLER_ASAP7_75t_R FILLER_227_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_227_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_227_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1190 ();
 FILLER_ASAP7_75t_R FILLER_227_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1287 ();
 DECAPx6_ASAP7_75t_R FILLER_228_918 ();
 FILLER_ASAP7_75t_R FILLER_228_932 ();
 DECAPx2_ASAP7_75t_R FILLER_228_940 ();
 DECAPx2_ASAP7_75t_R FILLER_228_952 ();
 FILLER_ASAP7_75t_R FILLER_228_958 ();
 DECAPx2_ASAP7_75t_R FILLER_228_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_228_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1167 ();
 FILLER_ASAP7_75t_R FILLER_228_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_228_1276 ();
 FILLER_ASAP7_75t_R FILLER_228_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_229_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_928 ();
 DECAPx10_ASAP7_75t_R FILLER_229_977 ();
 DECAPx4_ASAP7_75t_R FILLER_229_999 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1015 ();
 FILLER_ASAP7_75t_R FILLER_229_1021 ();
 FILLER_ASAP7_75t_R FILLER_229_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1057 ();
 FILLER_ASAP7_75t_R FILLER_229_1063 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1121 ();
 FILLER_ASAP7_75t_R FILLER_229_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1133 ();
 FILLER_ASAP7_75t_R FILLER_229_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1179 ();
 FILLER_ASAP7_75t_R FILLER_229_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1289 ();
 DECAPx6_ASAP7_75t_R FILLER_230_918 ();
 FILLER_ASAP7_75t_R FILLER_230_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_934 ();
 DECAPx10_ASAP7_75t_R FILLER_230_962 ();
 FILLER_ASAP7_75t_R FILLER_230_984 ();
 DECAPx1_ASAP7_75t_R FILLER_230_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_995 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1002 ();
 FILLER_ASAP7_75t_R FILLER_230_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1010 ();
 FILLER_ASAP7_75t_R FILLER_230_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1020 ();
 FILLER_ASAP7_75t_R FILLER_230_1074 ();
 FILLER_ASAP7_75t_R FILLER_230_1083 ();
 FILLER_ASAP7_75t_R FILLER_230_1112 ();
 FILLER_ASAP7_75t_R FILLER_230_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1140 ();
 FILLER_ASAP7_75t_R FILLER_230_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1276 ();
 FILLER_ASAP7_75t_R FILLER_230_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_231_918 ();
 DECAPx10_ASAP7_75t_R FILLER_231_940 ();
 DECAPx1_ASAP7_75t_R FILLER_231_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_966 ();
 DECAPx6_ASAP7_75t_R FILLER_231_975 ();
 FILLER_ASAP7_75t_R FILLER_231_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_991 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1026 ();
 FILLER_ASAP7_75t_R FILLER_231_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1036 ();
 FILLER_ASAP7_75t_R FILLER_231_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1088 ();
 FILLER_ASAP7_75t_R FILLER_231_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_231_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1163 ();
 FILLER_ASAP7_75t_R FILLER_231_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_232_918 ();
 DECAPx4_ASAP7_75t_R FILLER_232_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_954 ();
 DECAPx10_ASAP7_75t_R FILLER_232_964 ();
 DECAPx10_ASAP7_75t_R FILLER_232_986 ();
 DECAPx6_ASAP7_75t_R FILLER_232_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1057 ();
 FILLER_ASAP7_75t_R FILLER_232_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1072 ();
 FILLER_ASAP7_75t_R FILLER_232_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_233_918 ();
 FILLER_ASAP7_75t_R FILLER_233_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_930 ();
 DECAPx6_ASAP7_75t_R FILLER_233_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_966 ();
 DECAPx10_ASAP7_75t_R FILLER_233_973 ();
 DECAPx2_ASAP7_75t_R FILLER_233_995 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1090 ();
 FILLER_ASAP7_75t_R FILLER_233_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1098 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1105 ();
 FILLER_ASAP7_75t_R FILLER_233_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1281 ();
 FILLER_ASAP7_75t_R FILLER_233_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_234_918 ();
 DECAPx10_ASAP7_75t_R FILLER_234_940 ();
 DECAPx1_ASAP7_75t_R FILLER_234_962 ();
 DECAPx2_ASAP7_75t_R FILLER_234_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1062 ();
 FILLER_ASAP7_75t_R FILLER_234_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1106 ();
 FILLER_ASAP7_75t_R FILLER_234_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1130 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1152 ();
 FILLER_ASAP7_75t_R FILLER_234_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_235_918 ();
 DECAPx2_ASAP7_75t_R FILLER_235_940 ();
 DECAPx10_ASAP7_75t_R FILLER_235_951 ();
 DECAPx6_ASAP7_75t_R FILLER_235_973 ();
 FILLER_ASAP7_75t_R FILLER_235_987 ();
 DECAPx6_ASAP7_75t_R FILLER_235_996 ();
 FILLER_ASAP7_75t_R FILLER_235_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1134 ();
 FILLER_ASAP7_75t_R FILLER_235_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1164 ();
 FILLER_ASAP7_75t_R FILLER_235_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1276 ();
 FILLER_ASAP7_75t_R FILLER_235_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_236_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_932 ();
 DECAPx2_ASAP7_75t_R FILLER_236_954 ();
 FILLER_ASAP7_75t_R FILLER_236_960 ();
 DECAPx1_ASAP7_75t_R FILLER_236_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_976 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_236_1054 ();
 FILLER_ASAP7_75t_R FILLER_236_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_236_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_236_1276 ();
 FILLER_ASAP7_75t_R FILLER_236_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_237_918 ();
 DECAPx10_ASAP7_75t_R FILLER_237_940 ();
 DECAPx10_ASAP7_75t_R FILLER_237_962 ();
 DECAPx10_ASAP7_75t_R FILLER_237_984 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1056 ();
 FILLER_ASAP7_75t_R FILLER_237_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_237_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1113 ();
 DECAPx6_ASAP7_75t_R FILLER_237_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1281 ();
 FILLER_ASAP7_75t_R FILLER_237_1291 ();
 DECAPx4_ASAP7_75t_R FILLER_238_918 ();
 DECAPx10_ASAP7_75t_R FILLER_238_981 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_238_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_239_918 ();
 DECAPx4_ASAP7_75t_R FILLER_239_952 ();
 DECAPx10_ASAP7_75t_R FILLER_239_992 ();
 FILLER_ASAP7_75t_R FILLER_239_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1113 ();
 FILLER_ASAP7_75t_R FILLER_239_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_239_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_240_918 ();
 FILLER_ASAP7_75t_R FILLER_240_924 ();
 DECAPx2_ASAP7_75t_R FILLER_240_947 ();
 FILLER_ASAP7_75t_R FILLER_240_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_955 ();
 DECAPx2_ASAP7_75t_R FILLER_240_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_995 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_240_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_240_1080 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_240_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_241_918 ();
 DECAPx6_ASAP7_75t_R FILLER_241_940 ();
 DECAPx1_ASAP7_75t_R FILLER_241_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_958 ();
 DECAPx1_ASAP7_75t_R FILLER_241_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_978 ();
 DECAPx2_ASAP7_75t_R FILLER_241_1010 ();
 FILLER_ASAP7_75t_R FILLER_241_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_241_1116 ();
 FILLER_ASAP7_75t_R FILLER_241_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_241_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_242_918 ();
 DECAPx4_ASAP7_75t_R FILLER_242_940 ();
 FILLER_ASAP7_75t_R FILLER_242_950 ();
 DECAPx2_ASAP7_75t_R FILLER_242_984 ();
 FILLER_ASAP7_75t_R FILLER_242_990 ();
 DECAPx10_ASAP7_75t_R FILLER_242_998 ();
 DECAPx4_ASAP7_75t_R FILLER_242_1026 ();
 FILLER_ASAP7_75t_R FILLER_242_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1050 ();
 FILLER_ASAP7_75t_R FILLER_242_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_242_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_243_918 ();
 FILLER_ASAP7_75t_R FILLER_243_932 ();
 DECAPx10_ASAP7_75t_R FILLER_243_950 ();
 DECAPx10_ASAP7_75t_R FILLER_243_976 ();
 DECAPx10_ASAP7_75t_R FILLER_243_998 ();
 DECAPx4_ASAP7_75t_R FILLER_243_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_243_1037 ();
 FILLER_ASAP7_75t_R FILLER_243_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_243_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_244_918 ();
 DECAPx6_ASAP7_75t_R FILLER_244_940 ();
 DECAPx6_ASAP7_75t_R FILLER_244_975 ();
 DECAPx1_ASAP7_75t_R FILLER_244_989 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_244_1052 ();
 FILLER_ASAP7_75t_R FILLER_244_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1258 ();
 DECAPx4_ASAP7_75t_R FILLER_244_1280 ();
 FILLER_ASAP7_75t_R FILLER_244_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_245_918 ();
 DECAPx2_ASAP7_75t_R FILLER_245_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_938 ();
 DECAPx2_ASAP7_75t_R FILLER_245_949 ();
 FILLER_ASAP7_75t_R FILLER_245_955 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1006 ();
 FILLER_ASAP7_75t_R FILLER_245_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_246_918 ();
 DECAPx10_ASAP7_75t_R FILLER_246_967 ();
 DECAPx10_ASAP7_75t_R FILLER_246_989 ();
 FILLER_ASAP7_75t_R FILLER_246_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_246_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_247_918 ();
 DECAPx10_ASAP7_75t_R FILLER_247_940 ();
 DECAPx10_ASAP7_75t_R FILLER_247_962 ();
 DECAPx2_ASAP7_75t_R FILLER_247_984 ();
 FILLER_ASAP7_75t_R FILLER_247_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_992 ();
 DECAPx6_ASAP7_75t_R FILLER_247_997 ();
 DECAPx1_ASAP7_75t_R FILLER_247_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_247_1018 ();
 FILLER_ASAP7_75t_R FILLER_247_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_248_918 ();
 DECAPx1_ASAP7_75t_R FILLER_248_940 ();
 DECAPx6_ASAP7_75t_R FILLER_248_960 ();
 DECAPx2_ASAP7_75t_R FILLER_248_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_980 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_248_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_249_918 ();
 DECAPx4_ASAP7_75t_R FILLER_249_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_961 ();
 DECAPx1_ASAP7_75t_R FILLER_249_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_976 ();
 DECAPx10_ASAP7_75t_R FILLER_249_989 ();
 FILLER_ASAP7_75t_R FILLER_249_1011 ();
 FILLER_ASAP7_75t_R FILLER_249_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1269 ();
 FILLER_ASAP7_75t_R FILLER_249_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_250_918 ();
 DECAPx1_ASAP7_75t_R FILLER_250_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_952 ();
 FILLER_ASAP7_75t_R FILLER_250_963 ();
 DECAPx1_ASAP7_75t_R FILLER_250_980 ();
 DECAPx4_ASAP7_75t_R FILLER_250_996 ();
 FILLER_ASAP7_75t_R FILLER_250_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_250_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_251_918 ();
 DECAPx6_ASAP7_75t_R FILLER_251_935 ();
 FILLER_ASAP7_75t_R FILLER_251_956 ();
 DECAPx6_ASAP7_75t_R FILLER_251_973 ();
 DECAPx2_ASAP7_75t_R FILLER_251_987 ();
 DECAPx6_ASAP7_75t_R FILLER_251_996 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1257 ();
 DECAPx6_ASAP7_75t_R FILLER_251_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_252_918 ();
 DECAPx1_ASAP7_75t_R FILLER_252_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_944 ();
 DECAPx2_ASAP7_75t_R FILLER_252_950 ();
 DECAPx2_ASAP7_75t_R FILLER_252_961 ();
 FILLER_ASAP7_75t_R FILLER_252_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_969 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_252_1276 ();
 FILLER_ASAP7_75t_R FILLER_252_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_253_918 ();
 DECAPx2_ASAP7_75t_R FILLER_253_932 ();
 DECAPx1_ASAP7_75t_R FILLER_253_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_963 ();
 DECAPx10_ASAP7_75t_R FILLER_253_985 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_254_918 ();
 FILLER_ASAP7_75t_R FILLER_254_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_930 ();
 DECAPx10_ASAP7_75t_R FILLER_254_952 ();
 DECAPx10_ASAP7_75t_R FILLER_254_974 ();
 DECAPx10_ASAP7_75t_R FILLER_254_996 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_254_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_255_918 ();
 DECAPx10_ASAP7_75t_R FILLER_255_940 ();
 DECAPx10_ASAP7_75t_R FILLER_255_962 ();
 DECAPx10_ASAP7_75t_R FILLER_255_984 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_256_918 ();
 DECAPx10_ASAP7_75t_R FILLER_256_940 ();
 DECAPx10_ASAP7_75t_R FILLER_256_962 ();
 DECAPx10_ASAP7_75t_R FILLER_256_984 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_257_918 ();
 DECAPx10_ASAP7_75t_R FILLER_257_940 ();
 DECAPx10_ASAP7_75t_R FILLER_257_962 ();
 DECAPx10_ASAP7_75t_R FILLER_257_984 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_258_918 ();
 DECAPx10_ASAP7_75t_R FILLER_258_940 ();
 DECAPx10_ASAP7_75t_R FILLER_258_962 ();
 DECAPx10_ASAP7_75t_R FILLER_258_984 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_259_918 ();
 DECAPx10_ASAP7_75t_R FILLER_259_940 ();
 DECAPx10_ASAP7_75t_R FILLER_259_962 ();
 DECAPx10_ASAP7_75t_R FILLER_259_984 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_260_918 ();
 DECAPx10_ASAP7_75t_R FILLER_260_940 ();
 DECAPx10_ASAP7_75t_R FILLER_260_962 ();
 DECAPx10_ASAP7_75t_R FILLER_260_984 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_261_918 ();
 DECAPx10_ASAP7_75t_R FILLER_261_940 ();
 DECAPx10_ASAP7_75t_R FILLER_261_962 ();
 DECAPx10_ASAP7_75t_R FILLER_261_984 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_262_918 ();
 DECAPx10_ASAP7_75t_R FILLER_262_940 ();
 DECAPx10_ASAP7_75t_R FILLER_262_962 ();
 DECAPx10_ASAP7_75t_R FILLER_262_984 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_263_918 ();
 DECAPx10_ASAP7_75t_R FILLER_263_940 ();
 DECAPx10_ASAP7_75t_R FILLER_263_962 ();
 DECAPx10_ASAP7_75t_R FILLER_263_984 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_264_918 ();
 DECAPx10_ASAP7_75t_R FILLER_264_940 ();
 DECAPx10_ASAP7_75t_R FILLER_264_962 ();
 DECAPx10_ASAP7_75t_R FILLER_264_984 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_265_918 ();
 DECAPx10_ASAP7_75t_R FILLER_265_940 ();
 DECAPx10_ASAP7_75t_R FILLER_265_962 ();
 DECAPx10_ASAP7_75t_R FILLER_265_984 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_266_918 ();
 DECAPx10_ASAP7_75t_R FILLER_266_940 ();
 DECAPx10_ASAP7_75t_R FILLER_266_962 ();
 DECAPx10_ASAP7_75t_R FILLER_266_984 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_267_918 ();
 DECAPx10_ASAP7_75t_R FILLER_267_940 ();
 DECAPx10_ASAP7_75t_R FILLER_267_962 ();
 DECAPx10_ASAP7_75t_R FILLER_267_984 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_268_918 ();
 DECAPx10_ASAP7_75t_R FILLER_268_940 ();
 DECAPx10_ASAP7_75t_R FILLER_268_962 ();
 DECAPx10_ASAP7_75t_R FILLER_268_984 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_269_918 ();
 DECAPx10_ASAP7_75t_R FILLER_269_940 ();
 DECAPx10_ASAP7_75t_R FILLER_269_962 ();
 DECAPx10_ASAP7_75t_R FILLER_269_984 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_270_918 ();
 DECAPx10_ASAP7_75t_R FILLER_270_940 ();
 DECAPx10_ASAP7_75t_R FILLER_270_962 ();
 DECAPx10_ASAP7_75t_R FILLER_270_984 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_271_918 ();
 DECAPx10_ASAP7_75t_R FILLER_271_940 ();
 DECAPx10_ASAP7_75t_R FILLER_271_962 ();
 DECAPx10_ASAP7_75t_R FILLER_271_984 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_272_918 ();
 DECAPx10_ASAP7_75t_R FILLER_272_940 ();
 DECAPx10_ASAP7_75t_R FILLER_272_962 ();
 DECAPx10_ASAP7_75t_R FILLER_272_984 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_273_918 ();
 DECAPx10_ASAP7_75t_R FILLER_273_940 ();
 DECAPx10_ASAP7_75t_R FILLER_273_962 ();
 DECAPx10_ASAP7_75t_R FILLER_273_984 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_274_918 ();
 DECAPx10_ASAP7_75t_R FILLER_274_940 ();
 DECAPx10_ASAP7_75t_R FILLER_274_962 ();
 DECAPx10_ASAP7_75t_R FILLER_274_984 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_275_918 ();
 DECAPx10_ASAP7_75t_R FILLER_275_940 ();
 DECAPx10_ASAP7_75t_R FILLER_275_962 ();
 DECAPx10_ASAP7_75t_R FILLER_275_984 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_275_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_276_918 ();
 DECAPx10_ASAP7_75t_R FILLER_276_940 ();
 DECAPx10_ASAP7_75t_R FILLER_276_962 ();
 DECAPx10_ASAP7_75t_R FILLER_276_984 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_276_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_277_918 ();
 DECAPx10_ASAP7_75t_R FILLER_277_940 ();
 DECAPx10_ASAP7_75t_R FILLER_277_962 ();
 DECAPx10_ASAP7_75t_R FILLER_277_984 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_277_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_278_918 ();
 DECAPx10_ASAP7_75t_R FILLER_278_940 ();
 DECAPx10_ASAP7_75t_R FILLER_278_962 ();
 DECAPx10_ASAP7_75t_R FILLER_278_984 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_278_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_279_918 ();
 DECAPx10_ASAP7_75t_R FILLER_279_940 ();
 DECAPx10_ASAP7_75t_R FILLER_279_962 ();
 DECAPx10_ASAP7_75t_R FILLER_279_984 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_279_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_280_924 ();
 DECAPx10_ASAP7_75t_R FILLER_280_946 ();
 DECAPx10_ASAP7_75t_R FILLER_280_968 ();
 DECAPx10_ASAP7_75t_R FILLER_280_990 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_280_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_280_1276 ();
 FILLER_ASAP7_75t_R FILLER_280_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_281_918 ();
 DECAPx10_ASAP7_75t_R FILLER_281_940 ();
 DECAPx10_ASAP7_75t_R FILLER_281_962 ();
 DECAPx10_ASAP7_75t_R FILLER_281_984 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_281_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_282_918 ();
 DECAPx10_ASAP7_75t_R FILLER_282_940 ();
 DECAPx10_ASAP7_75t_R FILLER_282_962 ();
 DECAPx10_ASAP7_75t_R FILLER_282_984 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_282_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_283_918 ();
 DECAPx10_ASAP7_75t_R FILLER_283_940 ();
 DECAPx10_ASAP7_75t_R FILLER_283_962 ();
 DECAPx10_ASAP7_75t_R FILLER_283_984 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_283_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_284_918 ();
 DECAPx10_ASAP7_75t_R FILLER_284_940 ();
 DECAPx10_ASAP7_75t_R FILLER_284_962 ();
 DECAPx10_ASAP7_75t_R FILLER_284_984 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_284_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_285_918 ();
 DECAPx10_ASAP7_75t_R FILLER_285_940 ();
 DECAPx10_ASAP7_75t_R FILLER_285_962 ();
 DECAPx10_ASAP7_75t_R FILLER_285_984 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_285_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_286_918 ();
 DECAPx10_ASAP7_75t_R FILLER_286_940 ();
 DECAPx10_ASAP7_75t_R FILLER_286_962 ();
 DECAPx10_ASAP7_75t_R FILLER_286_984 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_286_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_287_918 ();
 DECAPx10_ASAP7_75t_R FILLER_287_940 ();
 DECAPx10_ASAP7_75t_R FILLER_287_962 ();
 DECAPx10_ASAP7_75t_R FILLER_287_984 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_287_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_288_918 ();
 DECAPx10_ASAP7_75t_R FILLER_288_940 ();
 DECAPx10_ASAP7_75t_R FILLER_288_962 ();
 DECAPx10_ASAP7_75t_R FILLER_288_984 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_288_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_289_918 ();
 DECAPx10_ASAP7_75t_R FILLER_289_940 ();
 DECAPx10_ASAP7_75t_R FILLER_289_962 ();
 DECAPx10_ASAP7_75t_R FILLER_289_984 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_289_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_290_918 ();
 DECAPx10_ASAP7_75t_R FILLER_290_940 ();
 DECAPx10_ASAP7_75t_R FILLER_290_962 ();
 DECAPx10_ASAP7_75t_R FILLER_290_984 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_290_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_291_918 ();
 DECAPx10_ASAP7_75t_R FILLER_291_940 ();
 DECAPx10_ASAP7_75t_R FILLER_291_962 ();
 DECAPx10_ASAP7_75t_R FILLER_291_984 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_291_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_292_918 ();
 DECAPx10_ASAP7_75t_R FILLER_292_940 ();
 DECAPx10_ASAP7_75t_R FILLER_292_962 ();
 DECAPx10_ASAP7_75t_R FILLER_292_984 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_292_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_293_918 ();
 DECAPx10_ASAP7_75t_R FILLER_293_940 ();
 DECAPx10_ASAP7_75t_R FILLER_293_962 ();
 DECAPx10_ASAP7_75t_R FILLER_293_984 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_293_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_294_918 ();
 DECAPx10_ASAP7_75t_R FILLER_294_940 ();
 DECAPx10_ASAP7_75t_R FILLER_294_962 ();
 DECAPx10_ASAP7_75t_R FILLER_294_984 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_294_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_1292 ();
endmodule
