VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA ibex_if_stage_via2_3_1600_480_1_5_320_320
  VIARULE M1M2_PR ;
  CUTSIZE 0.15 0.15 ;
  LAYERS met1 via met2 ;
  CUTSPACING 0.17 0.17 ;
  ENCLOSURE 0.085 0.165 0.055 0.085 ;
  ROWCOL 1 5 ;
END ibex_if_stage_via2_3_1600_480_1_5_320_320

VIA ibex_if_stage_via3_4_1600_480_1_4_400_400
  VIARULE M2M3_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met2 via2 met3 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.04 0.085 0.065 0.065 ;
  ROWCOL 1 4 ;
END ibex_if_stage_via3_4_1600_480_1_4_400_400

VIA ibex_if_stage_via4_5_1600_480_1_4_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.06 0.1 0.065 ;
  ROWCOL 1 4 ;
END ibex_if_stage_via4_5_1600_480_1_4_400_400

VIA ibex_if_stage_via5_6_1600_1600_1_1_1600_1600
  VIARULE M4M5_PR ;
  CUTSIZE 0.8 0.8 ;
  LAYERS met4 via4 met5 ;
  CUTSPACING 0.8 0.8 ;
  ENCLOSURE 0.4 0.19 0.31 0.4 ;
END ibex_if_stage_via5_6_1600_1600_1_1_1600_1600

MACRO ibex_if_stage
  FOREIGN ibex_if_stage 0 0 ;
  CLASS BLOCK ;
  SIZE 296.22 BY 296.22 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  27.72 273.92 273.58 275.52 ;
        RECT  27.72 246.72 273.58 248.32 ;
        RECT  27.72 219.52 273.58 221.12 ;
        RECT  27.72 192.32 273.58 193.92 ;
        RECT  27.72 165.12 273.58 166.72 ;
        RECT  27.72 137.92 273.58 139.52 ;
        RECT  27.72 110.72 273.58 112.32 ;
        RECT  27.72 83.52 273.58 85.12 ;
        RECT  27.72 56.32 273.58 57.92 ;
        RECT  27.72 29.12 273.58 30.72 ;
      LAYER met4 ;
        RECT  271.98 5.2 273.58 294 ;
        RECT  244.84 5.2 246.44 294 ;
        RECT  217.7 5.2 219.3 294 ;
        RECT  190.56 5.2 192.16 294 ;
        RECT  163.42 5.2 165.02 294 ;
        RECT  136.28 5.2 137.88 294 ;
        RECT  109.14 5.2 110.74 294 ;
        RECT  82 5.2 83.6 294 ;
        RECT  54.86 5.2 56.46 294 ;
        RECT  27.72 5.2 29.32 294 ;
      LAYER met1 ;
        RECT  1.38 293.52 294.86 294 ;
        RECT  1.38 288.08 294.86 288.56 ;
        RECT  1.38 282.64 294.86 283.12 ;
        RECT  1.38 277.2 294.86 277.68 ;
        RECT  1.38 271.76 294.86 272.24 ;
        RECT  1.38 266.32 294.86 266.8 ;
        RECT  1.38 260.88 294.86 261.36 ;
        RECT  1.38 255.44 294.86 255.92 ;
        RECT  1.38 250 294.86 250.48 ;
        RECT  1.38 244.56 294.86 245.04 ;
        RECT  1.38 239.12 294.86 239.6 ;
        RECT  1.38 233.68 294.86 234.16 ;
        RECT  1.38 228.24 294.86 228.72 ;
        RECT  1.38 222.8 294.86 223.28 ;
        RECT  1.38 217.36 294.86 217.84 ;
        RECT  1.38 211.92 294.86 212.4 ;
        RECT  1.38 206.48 294.86 206.96 ;
        RECT  1.38 201.04 294.86 201.52 ;
        RECT  1.38 195.6 294.86 196.08 ;
        RECT  1.38 190.16 294.86 190.64 ;
        RECT  1.38 184.72 294.86 185.2 ;
        RECT  1.38 179.28 294.86 179.76 ;
        RECT  1.38 173.84 294.86 174.32 ;
        RECT  1.38 168.4 294.86 168.88 ;
        RECT  1.38 162.96 294.86 163.44 ;
        RECT  1.38 157.52 294.86 158 ;
        RECT  1.38 152.08 294.86 152.56 ;
        RECT  1.38 146.64 294.86 147.12 ;
        RECT  1.38 141.2 294.86 141.68 ;
        RECT  1.38 135.76 294.86 136.24 ;
        RECT  1.38 130.32 294.86 130.8 ;
        RECT  1.38 124.88 294.86 125.36 ;
        RECT  1.38 119.44 294.86 119.92 ;
        RECT  1.38 114 294.86 114.48 ;
        RECT  1.38 108.56 294.86 109.04 ;
        RECT  1.38 103.12 294.86 103.6 ;
        RECT  1.38 97.68 294.86 98.16 ;
        RECT  1.38 92.24 294.86 92.72 ;
        RECT  1.38 86.8 294.86 87.28 ;
        RECT  1.38 81.36 294.86 81.84 ;
        RECT  1.38 75.92 294.86 76.4 ;
        RECT  1.38 70.48 294.86 70.96 ;
        RECT  1.38 65.04 294.86 65.52 ;
        RECT  1.38 59.6 294.86 60.08 ;
        RECT  1.38 54.16 294.86 54.64 ;
        RECT  1.38 48.72 294.86 49.2 ;
        RECT  1.38 43.28 294.86 43.76 ;
        RECT  1.38 37.84 294.86 38.32 ;
        RECT  1.38 32.4 294.86 32.88 ;
        RECT  1.38 26.96 294.86 27.44 ;
        RECT  1.38 21.52 294.86 22 ;
        RECT  1.38 16.08 294.86 16.56 ;
        RECT  1.38 10.64 294.86 11.12 ;
        RECT  1.38 5.2 294.86 5.68 ;
      VIA 272.78 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 272.78 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.64 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.5 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.36 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 274.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 247.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 220.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 193.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 165.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 138.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 111.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 84.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 57.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 29.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  271.99 293.595 273.57 293.925 ;
      VIA 272.78 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 293.575 273.55 293.945 ;
      VIA 272.78 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 288.155 273.57 288.485 ;
      VIA 272.78 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 288.135 273.55 288.505 ;
      VIA 272.78 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 282.715 273.57 283.045 ;
      VIA 272.78 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 282.695 273.55 283.065 ;
      VIA 272.78 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 277.275 273.57 277.605 ;
      VIA 272.78 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 277.255 273.55 277.625 ;
      VIA 272.78 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 271.835 273.57 272.165 ;
      VIA 272.78 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 271.815 273.55 272.185 ;
      VIA 272.78 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 266.395 273.57 266.725 ;
      VIA 272.78 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 266.375 273.55 266.745 ;
      VIA 272.78 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 260.955 273.57 261.285 ;
      VIA 272.78 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 260.935 273.55 261.305 ;
      VIA 272.78 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 255.515 273.57 255.845 ;
      VIA 272.78 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 255.495 273.55 255.865 ;
      VIA 272.78 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 250.075 273.57 250.405 ;
      VIA 272.78 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 250.055 273.55 250.425 ;
      VIA 272.78 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 244.635 273.57 244.965 ;
      VIA 272.78 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 244.615 273.55 244.985 ;
      VIA 272.78 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 239.195 273.57 239.525 ;
      VIA 272.78 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 239.175 273.55 239.545 ;
      VIA 272.78 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 233.755 273.57 234.085 ;
      VIA 272.78 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 233.735 273.55 234.105 ;
      VIA 272.78 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 228.315 273.57 228.645 ;
      VIA 272.78 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 228.295 273.55 228.665 ;
      VIA 272.78 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 222.875 273.57 223.205 ;
      VIA 272.78 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 222.855 273.55 223.225 ;
      VIA 272.78 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 217.435 273.57 217.765 ;
      VIA 272.78 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 217.415 273.55 217.785 ;
      VIA 272.78 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 211.995 273.57 212.325 ;
      VIA 272.78 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 211.975 273.55 212.345 ;
      VIA 272.78 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 206.555 273.57 206.885 ;
      VIA 272.78 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 206.535 273.55 206.905 ;
      VIA 272.78 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 201.115 273.57 201.445 ;
      VIA 272.78 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 201.095 273.55 201.465 ;
      VIA 272.78 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 195.675 273.57 196.005 ;
      VIA 272.78 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 195.655 273.55 196.025 ;
      VIA 272.78 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 190.235 273.57 190.565 ;
      VIA 272.78 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 190.215 273.55 190.585 ;
      VIA 272.78 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 184.795 273.57 185.125 ;
      VIA 272.78 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 184.775 273.55 185.145 ;
      VIA 272.78 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 179.355 273.57 179.685 ;
      VIA 272.78 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 179.335 273.55 179.705 ;
      VIA 272.78 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 173.915 273.57 174.245 ;
      VIA 272.78 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 173.895 273.55 174.265 ;
      VIA 272.78 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 168.475 273.57 168.805 ;
      VIA 272.78 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 168.455 273.55 168.825 ;
      VIA 272.78 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 163.035 273.57 163.365 ;
      VIA 272.78 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 163.015 273.55 163.385 ;
      VIA 272.78 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 157.595 273.57 157.925 ;
      VIA 272.78 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 157.575 273.55 157.945 ;
      VIA 272.78 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 152.155 273.57 152.485 ;
      VIA 272.78 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 152.135 273.55 152.505 ;
      VIA 272.78 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 146.715 273.57 147.045 ;
      VIA 272.78 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 146.695 273.55 147.065 ;
      VIA 272.78 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 141.275 273.57 141.605 ;
      VIA 272.78 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 141.255 273.55 141.625 ;
      VIA 272.78 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 135.835 273.57 136.165 ;
      VIA 272.78 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 135.815 273.55 136.185 ;
      VIA 272.78 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 130.395 273.57 130.725 ;
      VIA 272.78 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 130.375 273.55 130.745 ;
      VIA 272.78 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 124.955 273.57 125.285 ;
      VIA 272.78 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 124.935 273.55 125.305 ;
      VIA 272.78 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 119.515 273.57 119.845 ;
      VIA 272.78 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 119.495 273.55 119.865 ;
      VIA 272.78 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 114.075 273.57 114.405 ;
      VIA 272.78 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 114.055 273.55 114.425 ;
      VIA 272.78 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 108.635 273.57 108.965 ;
      VIA 272.78 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 108.615 273.55 108.985 ;
      VIA 272.78 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 103.195 273.57 103.525 ;
      VIA 272.78 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 103.175 273.55 103.545 ;
      VIA 272.78 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 97.755 273.57 98.085 ;
      VIA 272.78 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 97.735 273.55 98.105 ;
      VIA 272.78 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 92.315 273.57 92.645 ;
      VIA 272.78 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 92.295 273.55 92.665 ;
      VIA 272.78 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 86.875 273.57 87.205 ;
      VIA 272.78 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 86.855 273.55 87.225 ;
      VIA 272.78 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 81.435 273.57 81.765 ;
      VIA 272.78 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 81.415 273.55 81.785 ;
      VIA 272.78 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 75.995 273.57 76.325 ;
      VIA 272.78 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 75.975 273.55 76.345 ;
      VIA 272.78 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 70.555 273.57 70.885 ;
      VIA 272.78 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 70.535 273.55 70.905 ;
      VIA 272.78 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 65.115 273.57 65.445 ;
      VIA 272.78 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 65.095 273.55 65.465 ;
      VIA 272.78 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 59.675 273.57 60.005 ;
      VIA 272.78 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 59.655 273.55 60.025 ;
      VIA 272.78 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 54.235 273.57 54.565 ;
      VIA 272.78 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 54.215 273.55 54.585 ;
      VIA 272.78 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 48.795 273.57 49.125 ;
      VIA 272.78 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 48.775 273.55 49.145 ;
      VIA 272.78 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 43.355 273.57 43.685 ;
      VIA 272.78 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 43.335 273.55 43.705 ;
      VIA 272.78 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 37.915 273.57 38.245 ;
      VIA 272.78 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 37.895 273.55 38.265 ;
      VIA 272.78 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 32.475 273.57 32.805 ;
      VIA 272.78 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 32.455 273.55 32.825 ;
      VIA 272.78 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 27.035 273.57 27.365 ;
      VIA 272.78 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 27.015 273.55 27.385 ;
      VIA 272.78 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 21.595 273.57 21.925 ;
      VIA 272.78 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 21.575 273.55 21.945 ;
      VIA 272.78 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 16.155 273.57 16.485 ;
      VIA 272.78 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 16.135 273.55 16.505 ;
      VIA 272.78 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 10.715 273.57 11.045 ;
      VIA 272.78 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 10.695 273.55 11.065 ;
      VIA 272.78 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  271.99 5.275 273.57 5.605 ;
      VIA 272.78 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  272.01 5.255 273.55 5.625 ;
      VIA 272.78 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 272.78 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 293.595 246.43 293.925 ;
      VIA 245.64 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 293.575 246.41 293.945 ;
      VIA 245.64 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 288.155 246.43 288.485 ;
      VIA 245.64 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 288.135 246.41 288.505 ;
      VIA 245.64 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 282.715 246.43 283.045 ;
      VIA 245.64 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 282.695 246.41 283.065 ;
      VIA 245.64 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 277.275 246.43 277.605 ;
      VIA 245.64 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 277.255 246.41 277.625 ;
      VIA 245.64 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 271.835 246.43 272.165 ;
      VIA 245.64 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 271.815 246.41 272.185 ;
      VIA 245.64 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 266.395 246.43 266.725 ;
      VIA 245.64 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 266.375 246.41 266.745 ;
      VIA 245.64 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 260.955 246.43 261.285 ;
      VIA 245.64 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 260.935 246.41 261.305 ;
      VIA 245.64 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 255.515 246.43 255.845 ;
      VIA 245.64 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 255.495 246.41 255.865 ;
      VIA 245.64 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 250.075 246.43 250.405 ;
      VIA 245.64 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 250.055 246.41 250.425 ;
      VIA 245.64 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 244.635 246.43 244.965 ;
      VIA 245.64 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 244.615 246.41 244.985 ;
      VIA 245.64 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 239.195 246.43 239.525 ;
      VIA 245.64 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 239.175 246.41 239.545 ;
      VIA 245.64 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 233.755 246.43 234.085 ;
      VIA 245.64 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 233.735 246.41 234.105 ;
      VIA 245.64 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 228.315 246.43 228.645 ;
      VIA 245.64 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 228.295 246.41 228.665 ;
      VIA 245.64 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 222.875 246.43 223.205 ;
      VIA 245.64 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 222.855 246.41 223.225 ;
      VIA 245.64 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 217.435 246.43 217.765 ;
      VIA 245.64 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 217.415 246.41 217.785 ;
      VIA 245.64 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 211.995 246.43 212.325 ;
      VIA 245.64 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 211.975 246.41 212.345 ;
      VIA 245.64 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 206.555 246.43 206.885 ;
      VIA 245.64 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 206.535 246.41 206.905 ;
      VIA 245.64 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 201.115 246.43 201.445 ;
      VIA 245.64 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 201.095 246.41 201.465 ;
      VIA 245.64 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 195.675 246.43 196.005 ;
      VIA 245.64 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 195.655 246.41 196.025 ;
      VIA 245.64 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 190.235 246.43 190.565 ;
      VIA 245.64 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 190.215 246.41 190.585 ;
      VIA 245.64 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 184.795 246.43 185.125 ;
      VIA 245.64 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 184.775 246.41 185.145 ;
      VIA 245.64 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 179.355 246.43 179.685 ;
      VIA 245.64 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 179.335 246.41 179.705 ;
      VIA 245.64 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 173.915 246.43 174.245 ;
      VIA 245.64 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 173.895 246.41 174.265 ;
      VIA 245.64 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 168.475 246.43 168.805 ;
      VIA 245.64 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 168.455 246.41 168.825 ;
      VIA 245.64 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 163.035 246.43 163.365 ;
      VIA 245.64 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 163.015 246.41 163.385 ;
      VIA 245.64 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 157.595 246.43 157.925 ;
      VIA 245.64 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 157.575 246.41 157.945 ;
      VIA 245.64 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 152.155 246.43 152.485 ;
      VIA 245.64 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 152.135 246.41 152.505 ;
      VIA 245.64 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 146.715 246.43 147.045 ;
      VIA 245.64 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 146.695 246.41 147.065 ;
      VIA 245.64 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 141.275 246.43 141.605 ;
      VIA 245.64 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 141.255 246.41 141.625 ;
      VIA 245.64 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 135.835 246.43 136.165 ;
      VIA 245.64 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 135.815 246.41 136.185 ;
      VIA 245.64 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 130.395 246.43 130.725 ;
      VIA 245.64 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 130.375 246.41 130.745 ;
      VIA 245.64 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 124.955 246.43 125.285 ;
      VIA 245.64 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 124.935 246.41 125.305 ;
      VIA 245.64 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 119.515 246.43 119.845 ;
      VIA 245.64 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 119.495 246.41 119.865 ;
      VIA 245.64 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 114.075 246.43 114.405 ;
      VIA 245.64 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 114.055 246.41 114.425 ;
      VIA 245.64 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 108.635 246.43 108.965 ;
      VIA 245.64 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 108.615 246.41 108.985 ;
      VIA 245.64 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 103.195 246.43 103.525 ;
      VIA 245.64 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 103.175 246.41 103.545 ;
      VIA 245.64 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 97.755 246.43 98.085 ;
      VIA 245.64 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 97.735 246.41 98.105 ;
      VIA 245.64 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 92.315 246.43 92.645 ;
      VIA 245.64 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 92.295 246.41 92.665 ;
      VIA 245.64 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 86.875 246.43 87.205 ;
      VIA 245.64 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 86.855 246.41 87.225 ;
      VIA 245.64 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 81.435 246.43 81.765 ;
      VIA 245.64 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 81.415 246.41 81.785 ;
      VIA 245.64 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 75.995 246.43 76.325 ;
      VIA 245.64 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 75.975 246.41 76.345 ;
      VIA 245.64 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 70.555 246.43 70.885 ;
      VIA 245.64 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 70.535 246.41 70.905 ;
      VIA 245.64 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 65.115 246.43 65.445 ;
      VIA 245.64 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 65.095 246.41 65.465 ;
      VIA 245.64 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 59.675 246.43 60.005 ;
      VIA 245.64 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 59.655 246.41 60.025 ;
      VIA 245.64 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 54.235 246.43 54.565 ;
      VIA 245.64 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 54.215 246.41 54.585 ;
      VIA 245.64 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 48.795 246.43 49.125 ;
      VIA 245.64 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 48.775 246.41 49.145 ;
      VIA 245.64 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 43.355 246.43 43.685 ;
      VIA 245.64 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 43.335 246.41 43.705 ;
      VIA 245.64 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 37.915 246.43 38.245 ;
      VIA 245.64 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 37.895 246.41 38.265 ;
      VIA 245.64 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 32.475 246.43 32.805 ;
      VIA 245.64 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 32.455 246.41 32.825 ;
      VIA 245.64 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 27.035 246.43 27.365 ;
      VIA 245.64 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 27.015 246.41 27.385 ;
      VIA 245.64 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 21.595 246.43 21.925 ;
      VIA 245.64 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 21.575 246.41 21.945 ;
      VIA 245.64 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 16.155 246.43 16.485 ;
      VIA 245.64 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 16.135 246.41 16.505 ;
      VIA 245.64 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 10.715 246.43 11.045 ;
      VIA 245.64 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 10.695 246.41 11.065 ;
      VIA 245.64 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.85 5.275 246.43 5.605 ;
      VIA 245.64 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.87 5.255 246.41 5.625 ;
      VIA 245.64 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 245.64 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 293.595 219.29 293.925 ;
      VIA 218.5 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 293.575 219.27 293.945 ;
      VIA 218.5 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 288.155 219.29 288.485 ;
      VIA 218.5 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 288.135 219.27 288.505 ;
      VIA 218.5 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 282.715 219.29 283.045 ;
      VIA 218.5 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 282.695 219.27 283.065 ;
      VIA 218.5 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 277.275 219.29 277.605 ;
      VIA 218.5 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 277.255 219.27 277.625 ;
      VIA 218.5 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 271.835 219.29 272.165 ;
      VIA 218.5 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 271.815 219.27 272.185 ;
      VIA 218.5 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 266.395 219.29 266.725 ;
      VIA 218.5 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 266.375 219.27 266.745 ;
      VIA 218.5 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 260.955 219.29 261.285 ;
      VIA 218.5 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 260.935 219.27 261.305 ;
      VIA 218.5 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 255.515 219.29 255.845 ;
      VIA 218.5 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 255.495 219.27 255.865 ;
      VIA 218.5 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 250.075 219.29 250.405 ;
      VIA 218.5 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 250.055 219.27 250.425 ;
      VIA 218.5 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 244.635 219.29 244.965 ;
      VIA 218.5 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 244.615 219.27 244.985 ;
      VIA 218.5 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 239.195 219.29 239.525 ;
      VIA 218.5 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 239.175 219.27 239.545 ;
      VIA 218.5 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 233.755 219.29 234.085 ;
      VIA 218.5 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 233.735 219.27 234.105 ;
      VIA 218.5 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 228.315 219.29 228.645 ;
      VIA 218.5 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 228.295 219.27 228.665 ;
      VIA 218.5 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 222.875 219.29 223.205 ;
      VIA 218.5 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 222.855 219.27 223.225 ;
      VIA 218.5 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 217.435 219.29 217.765 ;
      VIA 218.5 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 217.415 219.27 217.785 ;
      VIA 218.5 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 211.995 219.29 212.325 ;
      VIA 218.5 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 211.975 219.27 212.345 ;
      VIA 218.5 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 206.555 219.29 206.885 ;
      VIA 218.5 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 206.535 219.27 206.905 ;
      VIA 218.5 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 201.115 219.29 201.445 ;
      VIA 218.5 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 201.095 219.27 201.465 ;
      VIA 218.5 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 195.675 219.29 196.005 ;
      VIA 218.5 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 195.655 219.27 196.025 ;
      VIA 218.5 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 190.235 219.29 190.565 ;
      VIA 218.5 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 190.215 219.27 190.585 ;
      VIA 218.5 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 184.795 219.29 185.125 ;
      VIA 218.5 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 184.775 219.27 185.145 ;
      VIA 218.5 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 179.355 219.29 179.685 ;
      VIA 218.5 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 179.335 219.27 179.705 ;
      VIA 218.5 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 173.915 219.29 174.245 ;
      VIA 218.5 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 173.895 219.27 174.265 ;
      VIA 218.5 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 168.475 219.29 168.805 ;
      VIA 218.5 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 168.455 219.27 168.825 ;
      VIA 218.5 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 163.035 219.29 163.365 ;
      VIA 218.5 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 163.015 219.27 163.385 ;
      VIA 218.5 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 157.595 219.29 157.925 ;
      VIA 218.5 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 157.575 219.27 157.945 ;
      VIA 218.5 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 152.155 219.29 152.485 ;
      VIA 218.5 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 152.135 219.27 152.505 ;
      VIA 218.5 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 146.715 219.29 147.045 ;
      VIA 218.5 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 146.695 219.27 147.065 ;
      VIA 218.5 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 141.275 219.29 141.605 ;
      VIA 218.5 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 141.255 219.27 141.625 ;
      VIA 218.5 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 135.835 219.29 136.165 ;
      VIA 218.5 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 135.815 219.27 136.185 ;
      VIA 218.5 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 130.395 219.29 130.725 ;
      VIA 218.5 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 130.375 219.27 130.745 ;
      VIA 218.5 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 124.955 219.29 125.285 ;
      VIA 218.5 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 124.935 219.27 125.305 ;
      VIA 218.5 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 119.515 219.29 119.845 ;
      VIA 218.5 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 119.495 219.27 119.865 ;
      VIA 218.5 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 114.075 219.29 114.405 ;
      VIA 218.5 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 114.055 219.27 114.425 ;
      VIA 218.5 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 108.635 219.29 108.965 ;
      VIA 218.5 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 108.615 219.27 108.985 ;
      VIA 218.5 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 103.195 219.29 103.525 ;
      VIA 218.5 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 103.175 219.27 103.545 ;
      VIA 218.5 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 97.755 219.29 98.085 ;
      VIA 218.5 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 97.735 219.27 98.105 ;
      VIA 218.5 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 92.315 219.29 92.645 ;
      VIA 218.5 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 92.295 219.27 92.665 ;
      VIA 218.5 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 86.875 219.29 87.205 ;
      VIA 218.5 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 86.855 219.27 87.225 ;
      VIA 218.5 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 81.435 219.29 81.765 ;
      VIA 218.5 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 81.415 219.27 81.785 ;
      VIA 218.5 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 75.995 219.29 76.325 ;
      VIA 218.5 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 75.975 219.27 76.345 ;
      VIA 218.5 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 70.555 219.29 70.885 ;
      VIA 218.5 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 70.535 219.27 70.905 ;
      VIA 218.5 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 65.115 219.29 65.445 ;
      VIA 218.5 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 65.095 219.27 65.465 ;
      VIA 218.5 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 59.675 219.29 60.005 ;
      VIA 218.5 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 59.655 219.27 60.025 ;
      VIA 218.5 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 54.235 219.29 54.565 ;
      VIA 218.5 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 54.215 219.27 54.585 ;
      VIA 218.5 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 48.795 219.29 49.125 ;
      VIA 218.5 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 48.775 219.27 49.145 ;
      VIA 218.5 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 43.355 219.29 43.685 ;
      VIA 218.5 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 43.335 219.27 43.705 ;
      VIA 218.5 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 37.915 219.29 38.245 ;
      VIA 218.5 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 37.895 219.27 38.265 ;
      VIA 218.5 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 32.475 219.29 32.805 ;
      VIA 218.5 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 32.455 219.27 32.825 ;
      VIA 218.5 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 27.035 219.29 27.365 ;
      VIA 218.5 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 27.015 219.27 27.385 ;
      VIA 218.5 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 21.595 219.29 21.925 ;
      VIA 218.5 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 21.575 219.27 21.945 ;
      VIA 218.5 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 16.155 219.29 16.485 ;
      VIA 218.5 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 16.135 219.27 16.505 ;
      VIA 218.5 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 10.715 219.29 11.045 ;
      VIA 218.5 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 10.695 219.27 11.065 ;
      VIA 218.5 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.71 5.275 219.29 5.605 ;
      VIA 218.5 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.73 5.255 219.27 5.625 ;
      VIA 218.5 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 218.5 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 293.595 192.15 293.925 ;
      VIA 191.36 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 293.575 192.13 293.945 ;
      VIA 191.36 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 288.155 192.15 288.485 ;
      VIA 191.36 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 288.135 192.13 288.505 ;
      VIA 191.36 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 282.715 192.15 283.045 ;
      VIA 191.36 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 282.695 192.13 283.065 ;
      VIA 191.36 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 277.275 192.15 277.605 ;
      VIA 191.36 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 277.255 192.13 277.625 ;
      VIA 191.36 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 271.835 192.15 272.165 ;
      VIA 191.36 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 271.815 192.13 272.185 ;
      VIA 191.36 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 266.395 192.15 266.725 ;
      VIA 191.36 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 266.375 192.13 266.745 ;
      VIA 191.36 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 260.955 192.15 261.285 ;
      VIA 191.36 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 260.935 192.13 261.305 ;
      VIA 191.36 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 255.515 192.15 255.845 ;
      VIA 191.36 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 255.495 192.13 255.865 ;
      VIA 191.36 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 250.075 192.15 250.405 ;
      VIA 191.36 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 250.055 192.13 250.425 ;
      VIA 191.36 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 244.635 192.15 244.965 ;
      VIA 191.36 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 244.615 192.13 244.985 ;
      VIA 191.36 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 239.195 192.15 239.525 ;
      VIA 191.36 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 239.175 192.13 239.545 ;
      VIA 191.36 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 233.755 192.15 234.085 ;
      VIA 191.36 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 233.735 192.13 234.105 ;
      VIA 191.36 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 228.315 192.15 228.645 ;
      VIA 191.36 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 228.295 192.13 228.665 ;
      VIA 191.36 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 222.875 192.15 223.205 ;
      VIA 191.36 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 222.855 192.13 223.225 ;
      VIA 191.36 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 217.435 192.15 217.765 ;
      VIA 191.36 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 217.415 192.13 217.785 ;
      VIA 191.36 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 211.995 192.15 212.325 ;
      VIA 191.36 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 211.975 192.13 212.345 ;
      VIA 191.36 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 206.555 192.15 206.885 ;
      VIA 191.36 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 206.535 192.13 206.905 ;
      VIA 191.36 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 201.115 192.15 201.445 ;
      VIA 191.36 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 201.095 192.13 201.465 ;
      VIA 191.36 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 195.675 192.15 196.005 ;
      VIA 191.36 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 195.655 192.13 196.025 ;
      VIA 191.36 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 190.235 192.15 190.565 ;
      VIA 191.36 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 190.215 192.13 190.585 ;
      VIA 191.36 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 184.795 192.15 185.125 ;
      VIA 191.36 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 184.775 192.13 185.145 ;
      VIA 191.36 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 179.355 192.15 179.685 ;
      VIA 191.36 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 179.335 192.13 179.705 ;
      VIA 191.36 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 173.915 192.15 174.245 ;
      VIA 191.36 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 173.895 192.13 174.265 ;
      VIA 191.36 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 168.475 192.15 168.805 ;
      VIA 191.36 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 168.455 192.13 168.825 ;
      VIA 191.36 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 163.035 192.15 163.365 ;
      VIA 191.36 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 163.015 192.13 163.385 ;
      VIA 191.36 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 157.595 192.15 157.925 ;
      VIA 191.36 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 157.575 192.13 157.945 ;
      VIA 191.36 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 152.155 192.15 152.485 ;
      VIA 191.36 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 152.135 192.13 152.505 ;
      VIA 191.36 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 146.715 192.15 147.045 ;
      VIA 191.36 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 146.695 192.13 147.065 ;
      VIA 191.36 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 141.275 192.15 141.605 ;
      VIA 191.36 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 141.255 192.13 141.625 ;
      VIA 191.36 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 135.835 192.15 136.165 ;
      VIA 191.36 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 135.815 192.13 136.185 ;
      VIA 191.36 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 130.395 192.15 130.725 ;
      VIA 191.36 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 130.375 192.13 130.745 ;
      VIA 191.36 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 124.955 192.15 125.285 ;
      VIA 191.36 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 124.935 192.13 125.305 ;
      VIA 191.36 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 119.515 192.15 119.845 ;
      VIA 191.36 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 119.495 192.13 119.865 ;
      VIA 191.36 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 114.075 192.15 114.405 ;
      VIA 191.36 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 114.055 192.13 114.425 ;
      VIA 191.36 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 108.635 192.15 108.965 ;
      VIA 191.36 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 108.615 192.13 108.985 ;
      VIA 191.36 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 103.195 192.15 103.525 ;
      VIA 191.36 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 103.175 192.13 103.545 ;
      VIA 191.36 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 97.755 192.15 98.085 ;
      VIA 191.36 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 97.735 192.13 98.105 ;
      VIA 191.36 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 92.315 192.15 92.645 ;
      VIA 191.36 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 92.295 192.13 92.665 ;
      VIA 191.36 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 86.875 192.15 87.205 ;
      VIA 191.36 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 86.855 192.13 87.225 ;
      VIA 191.36 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 81.435 192.15 81.765 ;
      VIA 191.36 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 81.415 192.13 81.785 ;
      VIA 191.36 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 75.995 192.15 76.325 ;
      VIA 191.36 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 75.975 192.13 76.345 ;
      VIA 191.36 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 70.555 192.15 70.885 ;
      VIA 191.36 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 70.535 192.13 70.905 ;
      VIA 191.36 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 65.115 192.15 65.445 ;
      VIA 191.36 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 65.095 192.13 65.465 ;
      VIA 191.36 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 59.675 192.15 60.005 ;
      VIA 191.36 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 59.655 192.13 60.025 ;
      VIA 191.36 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 54.235 192.15 54.565 ;
      VIA 191.36 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 54.215 192.13 54.585 ;
      VIA 191.36 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 48.795 192.15 49.125 ;
      VIA 191.36 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 48.775 192.13 49.145 ;
      VIA 191.36 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 43.355 192.15 43.685 ;
      VIA 191.36 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 43.335 192.13 43.705 ;
      VIA 191.36 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 37.915 192.15 38.245 ;
      VIA 191.36 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 37.895 192.13 38.265 ;
      VIA 191.36 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 32.475 192.15 32.805 ;
      VIA 191.36 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 32.455 192.13 32.825 ;
      VIA 191.36 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 27.035 192.15 27.365 ;
      VIA 191.36 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 27.015 192.13 27.385 ;
      VIA 191.36 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 21.595 192.15 21.925 ;
      VIA 191.36 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 21.575 192.13 21.945 ;
      VIA 191.36 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 16.155 192.15 16.485 ;
      VIA 191.36 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 16.135 192.13 16.505 ;
      VIA 191.36 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 10.715 192.15 11.045 ;
      VIA 191.36 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 10.695 192.13 11.065 ;
      VIA 191.36 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.57 5.275 192.15 5.605 ;
      VIA 191.36 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.59 5.255 192.13 5.625 ;
      VIA 191.36 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 191.36 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 293.595 165.01 293.925 ;
      VIA 164.22 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 293.575 164.99 293.945 ;
      VIA 164.22 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 288.155 165.01 288.485 ;
      VIA 164.22 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 288.135 164.99 288.505 ;
      VIA 164.22 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 282.715 165.01 283.045 ;
      VIA 164.22 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 282.695 164.99 283.065 ;
      VIA 164.22 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 277.275 165.01 277.605 ;
      VIA 164.22 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 277.255 164.99 277.625 ;
      VIA 164.22 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 271.835 165.01 272.165 ;
      VIA 164.22 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 271.815 164.99 272.185 ;
      VIA 164.22 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 266.395 165.01 266.725 ;
      VIA 164.22 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 266.375 164.99 266.745 ;
      VIA 164.22 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 260.955 165.01 261.285 ;
      VIA 164.22 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 260.935 164.99 261.305 ;
      VIA 164.22 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 255.515 165.01 255.845 ;
      VIA 164.22 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 255.495 164.99 255.865 ;
      VIA 164.22 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 250.075 165.01 250.405 ;
      VIA 164.22 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 250.055 164.99 250.425 ;
      VIA 164.22 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 244.635 165.01 244.965 ;
      VIA 164.22 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 244.615 164.99 244.985 ;
      VIA 164.22 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 239.195 165.01 239.525 ;
      VIA 164.22 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 239.175 164.99 239.545 ;
      VIA 164.22 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 233.755 165.01 234.085 ;
      VIA 164.22 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 233.735 164.99 234.105 ;
      VIA 164.22 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 228.315 165.01 228.645 ;
      VIA 164.22 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 228.295 164.99 228.665 ;
      VIA 164.22 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 222.875 165.01 223.205 ;
      VIA 164.22 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 222.855 164.99 223.225 ;
      VIA 164.22 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 217.435 165.01 217.765 ;
      VIA 164.22 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 217.415 164.99 217.785 ;
      VIA 164.22 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 211.995 165.01 212.325 ;
      VIA 164.22 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 211.975 164.99 212.345 ;
      VIA 164.22 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 206.555 165.01 206.885 ;
      VIA 164.22 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 206.535 164.99 206.905 ;
      VIA 164.22 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 201.115 165.01 201.445 ;
      VIA 164.22 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 201.095 164.99 201.465 ;
      VIA 164.22 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 195.675 165.01 196.005 ;
      VIA 164.22 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 195.655 164.99 196.025 ;
      VIA 164.22 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 190.235 165.01 190.565 ;
      VIA 164.22 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 190.215 164.99 190.585 ;
      VIA 164.22 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 184.795 165.01 185.125 ;
      VIA 164.22 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 184.775 164.99 185.145 ;
      VIA 164.22 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 179.355 165.01 179.685 ;
      VIA 164.22 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 179.335 164.99 179.705 ;
      VIA 164.22 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 173.915 165.01 174.245 ;
      VIA 164.22 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 173.895 164.99 174.265 ;
      VIA 164.22 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 168.475 165.01 168.805 ;
      VIA 164.22 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 168.455 164.99 168.825 ;
      VIA 164.22 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 163.035 165.01 163.365 ;
      VIA 164.22 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 163.015 164.99 163.385 ;
      VIA 164.22 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 157.595 165.01 157.925 ;
      VIA 164.22 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 157.575 164.99 157.945 ;
      VIA 164.22 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 152.155 165.01 152.485 ;
      VIA 164.22 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 152.135 164.99 152.505 ;
      VIA 164.22 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 146.715 165.01 147.045 ;
      VIA 164.22 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 146.695 164.99 147.065 ;
      VIA 164.22 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 141.275 165.01 141.605 ;
      VIA 164.22 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 141.255 164.99 141.625 ;
      VIA 164.22 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 135.835 165.01 136.165 ;
      VIA 164.22 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 135.815 164.99 136.185 ;
      VIA 164.22 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 130.395 165.01 130.725 ;
      VIA 164.22 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 130.375 164.99 130.745 ;
      VIA 164.22 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 124.955 165.01 125.285 ;
      VIA 164.22 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 124.935 164.99 125.305 ;
      VIA 164.22 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 119.515 165.01 119.845 ;
      VIA 164.22 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 119.495 164.99 119.865 ;
      VIA 164.22 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 114.075 165.01 114.405 ;
      VIA 164.22 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 114.055 164.99 114.425 ;
      VIA 164.22 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 108.635 165.01 108.965 ;
      VIA 164.22 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 108.615 164.99 108.985 ;
      VIA 164.22 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 103.195 165.01 103.525 ;
      VIA 164.22 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 103.175 164.99 103.545 ;
      VIA 164.22 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 97.755 165.01 98.085 ;
      VIA 164.22 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 97.735 164.99 98.105 ;
      VIA 164.22 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 92.315 165.01 92.645 ;
      VIA 164.22 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 92.295 164.99 92.665 ;
      VIA 164.22 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 86.875 165.01 87.205 ;
      VIA 164.22 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 86.855 164.99 87.225 ;
      VIA 164.22 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 81.435 165.01 81.765 ;
      VIA 164.22 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 81.415 164.99 81.785 ;
      VIA 164.22 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 75.995 165.01 76.325 ;
      VIA 164.22 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 75.975 164.99 76.345 ;
      VIA 164.22 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 70.555 165.01 70.885 ;
      VIA 164.22 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 70.535 164.99 70.905 ;
      VIA 164.22 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 65.115 165.01 65.445 ;
      VIA 164.22 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 65.095 164.99 65.465 ;
      VIA 164.22 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 59.675 165.01 60.005 ;
      VIA 164.22 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 59.655 164.99 60.025 ;
      VIA 164.22 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 54.235 165.01 54.565 ;
      VIA 164.22 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 54.215 164.99 54.585 ;
      VIA 164.22 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 48.795 165.01 49.125 ;
      VIA 164.22 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 48.775 164.99 49.145 ;
      VIA 164.22 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 43.355 165.01 43.685 ;
      VIA 164.22 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 43.335 164.99 43.705 ;
      VIA 164.22 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 37.915 165.01 38.245 ;
      VIA 164.22 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 37.895 164.99 38.265 ;
      VIA 164.22 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 32.475 165.01 32.805 ;
      VIA 164.22 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 32.455 164.99 32.825 ;
      VIA 164.22 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 27.035 165.01 27.365 ;
      VIA 164.22 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 27.015 164.99 27.385 ;
      VIA 164.22 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 21.595 165.01 21.925 ;
      VIA 164.22 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 21.575 164.99 21.945 ;
      VIA 164.22 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 16.155 165.01 16.485 ;
      VIA 164.22 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 16.135 164.99 16.505 ;
      VIA 164.22 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 10.715 165.01 11.045 ;
      VIA 164.22 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 10.695 164.99 11.065 ;
      VIA 164.22 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 5.275 165.01 5.605 ;
      VIA 164.22 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 5.255 164.99 5.625 ;
      VIA 164.22 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 293.595 137.87 293.925 ;
      VIA 137.08 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 293.575 137.85 293.945 ;
      VIA 137.08 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 288.155 137.87 288.485 ;
      VIA 137.08 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 288.135 137.85 288.505 ;
      VIA 137.08 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 282.715 137.87 283.045 ;
      VIA 137.08 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 282.695 137.85 283.065 ;
      VIA 137.08 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 277.275 137.87 277.605 ;
      VIA 137.08 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 277.255 137.85 277.625 ;
      VIA 137.08 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 271.835 137.87 272.165 ;
      VIA 137.08 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 271.815 137.85 272.185 ;
      VIA 137.08 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 266.395 137.87 266.725 ;
      VIA 137.08 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 266.375 137.85 266.745 ;
      VIA 137.08 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 260.955 137.87 261.285 ;
      VIA 137.08 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 260.935 137.85 261.305 ;
      VIA 137.08 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 255.515 137.87 255.845 ;
      VIA 137.08 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 255.495 137.85 255.865 ;
      VIA 137.08 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 250.075 137.87 250.405 ;
      VIA 137.08 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 250.055 137.85 250.425 ;
      VIA 137.08 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 244.635 137.87 244.965 ;
      VIA 137.08 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 244.615 137.85 244.985 ;
      VIA 137.08 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 239.195 137.87 239.525 ;
      VIA 137.08 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 239.175 137.85 239.545 ;
      VIA 137.08 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 233.755 137.87 234.085 ;
      VIA 137.08 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 233.735 137.85 234.105 ;
      VIA 137.08 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 228.315 137.87 228.645 ;
      VIA 137.08 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 228.295 137.85 228.665 ;
      VIA 137.08 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 222.875 137.87 223.205 ;
      VIA 137.08 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 222.855 137.85 223.225 ;
      VIA 137.08 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 217.435 137.87 217.765 ;
      VIA 137.08 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 217.415 137.85 217.785 ;
      VIA 137.08 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 211.995 137.87 212.325 ;
      VIA 137.08 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 211.975 137.85 212.345 ;
      VIA 137.08 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 206.555 137.87 206.885 ;
      VIA 137.08 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 206.535 137.85 206.905 ;
      VIA 137.08 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 201.115 137.87 201.445 ;
      VIA 137.08 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 201.095 137.85 201.465 ;
      VIA 137.08 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 195.675 137.87 196.005 ;
      VIA 137.08 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 195.655 137.85 196.025 ;
      VIA 137.08 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 190.235 137.87 190.565 ;
      VIA 137.08 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 190.215 137.85 190.585 ;
      VIA 137.08 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 184.795 137.87 185.125 ;
      VIA 137.08 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 184.775 137.85 185.145 ;
      VIA 137.08 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 179.355 137.87 179.685 ;
      VIA 137.08 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 179.335 137.85 179.705 ;
      VIA 137.08 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 173.915 137.87 174.245 ;
      VIA 137.08 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 173.895 137.85 174.265 ;
      VIA 137.08 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 168.475 137.87 168.805 ;
      VIA 137.08 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 168.455 137.85 168.825 ;
      VIA 137.08 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 163.035 137.87 163.365 ;
      VIA 137.08 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 163.015 137.85 163.385 ;
      VIA 137.08 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 157.595 137.87 157.925 ;
      VIA 137.08 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 157.575 137.85 157.945 ;
      VIA 137.08 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 152.155 137.87 152.485 ;
      VIA 137.08 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 152.135 137.85 152.505 ;
      VIA 137.08 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 146.715 137.87 147.045 ;
      VIA 137.08 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 146.695 137.85 147.065 ;
      VIA 137.08 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 141.275 137.87 141.605 ;
      VIA 137.08 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 141.255 137.85 141.625 ;
      VIA 137.08 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 135.835 137.87 136.165 ;
      VIA 137.08 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 135.815 137.85 136.185 ;
      VIA 137.08 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 130.395 137.87 130.725 ;
      VIA 137.08 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 130.375 137.85 130.745 ;
      VIA 137.08 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 124.955 137.87 125.285 ;
      VIA 137.08 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 124.935 137.85 125.305 ;
      VIA 137.08 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 119.515 137.87 119.845 ;
      VIA 137.08 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 119.495 137.85 119.865 ;
      VIA 137.08 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 114.075 137.87 114.405 ;
      VIA 137.08 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 114.055 137.85 114.425 ;
      VIA 137.08 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 108.635 137.87 108.965 ;
      VIA 137.08 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 108.615 137.85 108.985 ;
      VIA 137.08 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 103.195 137.87 103.525 ;
      VIA 137.08 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 103.175 137.85 103.545 ;
      VIA 137.08 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 97.755 137.87 98.085 ;
      VIA 137.08 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 97.735 137.85 98.105 ;
      VIA 137.08 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 92.315 137.87 92.645 ;
      VIA 137.08 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 92.295 137.85 92.665 ;
      VIA 137.08 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 86.875 137.87 87.205 ;
      VIA 137.08 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 86.855 137.85 87.225 ;
      VIA 137.08 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 81.435 137.87 81.765 ;
      VIA 137.08 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 81.415 137.85 81.785 ;
      VIA 137.08 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 75.995 137.87 76.325 ;
      VIA 137.08 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 75.975 137.85 76.345 ;
      VIA 137.08 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 70.555 137.87 70.885 ;
      VIA 137.08 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 70.535 137.85 70.905 ;
      VIA 137.08 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 65.115 137.87 65.445 ;
      VIA 137.08 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 65.095 137.85 65.465 ;
      VIA 137.08 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 59.675 137.87 60.005 ;
      VIA 137.08 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 59.655 137.85 60.025 ;
      VIA 137.08 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 54.235 137.87 54.565 ;
      VIA 137.08 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 54.215 137.85 54.585 ;
      VIA 137.08 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 48.795 137.87 49.125 ;
      VIA 137.08 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 48.775 137.85 49.145 ;
      VIA 137.08 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 43.355 137.87 43.685 ;
      VIA 137.08 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 43.335 137.85 43.705 ;
      VIA 137.08 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 37.915 137.87 38.245 ;
      VIA 137.08 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 37.895 137.85 38.265 ;
      VIA 137.08 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 32.475 137.87 32.805 ;
      VIA 137.08 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 32.455 137.85 32.825 ;
      VIA 137.08 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 27.035 137.87 27.365 ;
      VIA 137.08 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 27.015 137.85 27.385 ;
      VIA 137.08 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 21.595 137.87 21.925 ;
      VIA 137.08 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 21.575 137.85 21.945 ;
      VIA 137.08 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 16.155 137.87 16.485 ;
      VIA 137.08 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 16.135 137.85 16.505 ;
      VIA 137.08 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 10.715 137.87 11.045 ;
      VIA 137.08 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 10.695 137.85 11.065 ;
      VIA 137.08 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 5.275 137.87 5.605 ;
      VIA 137.08 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 5.255 137.85 5.625 ;
      VIA 137.08 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 293.595 110.73 293.925 ;
      VIA 109.94 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 293.575 110.71 293.945 ;
      VIA 109.94 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 288.155 110.73 288.485 ;
      VIA 109.94 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 288.135 110.71 288.505 ;
      VIA 109.94 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 282.715 110.73 283.045 ;
      VIA 109.94 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 282.695 110.71 283.065 ;
      VIA 109.94 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 277.275 110.73 277.605 ;
      VIA 109.94 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 277.255 110.71 277.625 ;
      VIA 109.94 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 271.835 110.73 272.165 ;
      VIA 109.94 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 271.815 110.71 272.185 ;
      VIA 109.94 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 266.395 110.73 266.725 ;
      VIA 109.94 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 266.375 110.71 266.745 ;
      VIA 109.94 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 260.955 110.73 261.285 ;
      VIA 109.94 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 260.935 110.71 261.305 ;
      VIA 109.94 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 255.515 110.73 255.845 ;
      VIA 109.94 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 255.495 110.71 255.865 ;
      VIA 109.94 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 250.075 110.73 250.405 ;
      VIA 109.94 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 250.055 110.71 250.425 ;
      VIA 109.94 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 244.635 110.73 244.965 ;
      VIA 109.94 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 244.615 110.71 244.985 ;
      VIA 109.94 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 239.195 110.73 239.525 ;
      VIA 109.94 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 239.175 110.71 239.545 ;
      VIA 109.94 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 233.755 110.73 234.085 ;
      VIA 109.94 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 233.735 110.71 234.105 ;
      VIA 109.94 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 228.315 110.73 228.645 ;
      VIA 109.94 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 228.295 110.71 228.665 ;
      VIA 109.94 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 222.875 110.73 223.205 ;
      VIA 109.94 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 222.855 110.71 223.225 ;
      VIA 109.94 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 217.435 110.73 217.765 ;
      VIA 109.94 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 217.415 110.71 217.785 ;
      VIA 109.94 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 211.995 110.73 212.325 ;
      VIA 109.94 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 211.975 110.71 212.345 ;
      VIA 109.94 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 206.555 110.73 206.885 ;
      VIA 109.94 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 206.535 110.71 206.905 ;
      VIA 109.94 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 201.115 110.73 201.445 ;
      VIA 109.94 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 201.095 110.71 201.465 ;
      VIA 109.94 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 195.675 110.73 196.005 ;
      VIA 109.94 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 195.655 110.71 196.025 ;
      VIA 109.94 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 190.235 110.73 190.565 ;
      VIA 109.94 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 190.215 110.71 190.585 ;
      VIA 109.94 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 184.795 110.73 185.125 ;
      VIA 109.94 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 184.775 110.71 185.145 ;
      VIA 109.94 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 179.355 110.73 179.685 ;
      VIA 109.94 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 179.335 110.71 179.705 ;
      VIA 109.94 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 173.915 110.73 174.245 ;
      VIA 109.94 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 173.895 110.71 174.265 ;
      VIA 109.94 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 168.475 110.73 168.805 ;
      VIA 109.94 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 168.455 110.71 168.825 ;
      VIA 109.94 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 163.035 110.73 163.365 ;
      VIA 109.94 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 163.015 110.71 163.385 ;
      VIA 109.94 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 157.595 110.73 157.925 ;
      VIA 109.94 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 157.575 110.71 157.945 ;
      VIA 109.94 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 152.155 110.73 152.485 ;
      VIA 109.94 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 152.135 110.71 152.505 ;
      VIA 109.94 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 146.715 110.73 147.045 ;
      VIA 109.94 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 146.695 110.71 147.065 ;
      VIA 109.94 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 141.275 110.73 141.605 ;
      VIA 109.94 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 141.255 110.71 141.625 ;
      VIA 109.94 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 135.835 110.73 136.165 ;
      VIA 109.94 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 135.815 110.71 136.185 ;
      VIA 109.94 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 130.395 110.73 130.725 ;
      VIA 109.94 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 130.375 110.71 130.745 ;
      VIA 109.94 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 124.955 110.73 125.285 ;
      VIA 109.94 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 124.935 110.71 125.305 ;
      VIA 109.94 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 119.515 110.73 119.845 ;
      VIA 109.94 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 119.495 110.71 119.865 ;
      VIA 109.94 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 114.075 110.73 114.405 ;
      VIA 109.94 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 114.055 110.71 114.425 ;
      VIA 109.94 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 108.635 110.73 108.965 ;
      VIA 109.94 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 108.615 110.71 108.985 ;
      VIA 109.94 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 103.195 110.73 103.525 ;
      VIA 109.94 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 103.175 110.71 103.545 ;
      VIA 109.94 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 97.755 110.73 98.085 ;
      VIA 109.94 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 97.735 110.71 98.105 ;
      VIA 109.94 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 92.315 110.73 92.645 ;
      VIA 109.94 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 92.295 110.71 92.665 ;
      VIA 109.94 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 86.875 110.73 87.205 ;
      VIA 109.94 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 86.855 110.71 87.225 ;
      VIA 109.94 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 81.435 110.73 81.765 ;
      VIA 109.94 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 81.415 110.71 81.785 ;
      VIA 109.94 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 75.995 110.73 76.325 ;
      VIA 109.94 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 75.975 110.71 76.345 ;
      VIA 109.94 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 70.555 110.73 70.885 ;
      VIA 109.94 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 70.535 110.71 70.905 ;
      VIA 109.94 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 65.115 110.73 65.445 ;
      VIA 109.94 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 65.095 110.71 65.465 ;
      VIA 109.94 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 59.675 110.73 60.005 ;
      VIA 109.94 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 59.655 110.71 60.025 ;
      VIA 109.94 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 54.235 110.73 54.565 ;
      VIA 109.94 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 54.215 110.71 54.585 ;
      VIA 109.94 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 48.795 110.73 49.125 ;
      VIA 109.94 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 48.775 110.71 49.145 ;
      VIA 109.94 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 43.355 110.73 43.685 ;
      VIA 109.94 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 43.335 110.71 43.705 ;
      VIA 109.94 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 37.915 110.73 38.245 ;
      VIA 109.94 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 37.895 110.71 38.265 ;
      VIA 109.94 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 32.475 110.73 32.805 ;
      VIA 109.94 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 32.455 110.71 32.825 ;
      VIA 109.94 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 27.035 110.73 27.365 ;
      VIA 109.94 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 27.015 110.71 27.385 ;
      VIA 109.94 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 21.595 110.73 21.925 ;
      VIA 109.94 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 21.575 110.71 21.945 ;
      VIA 109.94 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 16.155 110.73 16.485 ;
      VIA 109.94 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 16.135 110.71 16.505 ;
      VIA 109.94 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 10.715 110.73 11.045 ;
      VIA 109.94 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 10.695 110.71 11.065 ;
      VIA 109.94 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 5.275 110.73 5.605 ;
      VIA 109.94 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 5.255 110.71 5.625 ;
      VIA 109.94 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 293.595 83.59 293.925 ;
      VIA 82.8 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 293.575 83.57 293.945 ;
      VIA 82.8 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 288.155 83.59 288.485 ;
      VIA 82.8 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 288.135 83.57 288.505 ;
      VIA 82.8 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 282.715 83.59 283.045 ;
      VIA 82.8 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 282.695 83.57 283.065 ;
      VIA 82.8 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 277.275 83.59 277.605 ;
      VIA 82.8 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 277.255 83.57 277.625 ;
      VIA 82.8 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 271.835 83.59 272.165 ;
      VIA 82.8 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 271.815 83.57 272.185 ;
      VIA 82.8 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 266.395 83.59 266.725 ;
      VIA 82.8 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 266.375 83.57 266.745 ;
      VIA 82.8 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 260.955 83.59 261.285 ;
      VIA 82.8 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 260.935 83.57 261.305 ;
      VIA 82.8 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 255.515 83.59 255.845 ;
      VIA 82.8 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 255.495 83.57 255.865 ;
      VIA 82.8 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 250.075 83.59 250.405 ;
      VIA 82.8 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 250.055 83.57 250.425 ;
      VIA 82.8 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 244.635 83.59 244.965 ;
      VIA 82.8 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 244.615 83.57 244.985 ;
      VIA 82.8 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 239.195 83.59 239.525 ;
      VIA 82.8 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 239.175 83.57 239.545 ;
      VIA 82.8 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 233.755 83.59 234.085 ;
      VIA 82.8 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 233.735 83.57 234.105 ;
      VIA 82.8 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 228.315 83.59 228.645 ;
      VIA 82.8 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 228.295 83.57 228.665 ;
      VIA 82.8 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 222.875 83.59 223.205 ;
      VIA 82.8 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 222.855 83.57 223.225 ;
      VIA 82.8 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 217.435 83.59 217.765 ;
      VIA 82.8 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 217.415 83.57 217.785 ;
      VIA 82.8 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 211.995 83.59 212.325 ;
      VIA 82.8 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 211.975 83.57 212.345 ;
      VIA 82.8 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 206.555 83.59 206.885 ;
      VIA 82.8 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 206.535 83.57 206.905 ;
      VIA 82.8 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 201.115 83.59 201.445 ;
      VIA 82.8 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 201.095 83.57 201.465 ;
      VIA 82.8 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 195.675 83.59 196.005 ;
      VIA 82.8 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 195.655 83.57 196.025 ;
      VIA 82.8 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 190.235 83.59 190.565 ;
      VIA 82.8 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 190.215 83.57 190.585 ;
      VIA 82.8 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 184.795 83.59 185.125 ;
      VIA 82.8 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 184.775 83.57 185.145 ;
      VIA 82.8 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 179.355 83.59 179.685 ;
      VIA 82.8 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 179.335 83.57 179.705 ;
      VIA 82.8 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 173.915 83.59 174.245 ;
      VIA 82.8 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 173.895 83.57 174.265 ;
      VIA 82.8 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 168.475 83.59 168.805 ;
      VIA 82.8 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 168.455 83.57 168.825 ;
      VIA 82.8 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 163.035 83.59 163.365 ;
      VIA 82.8 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 163.015 83.57 163.385 ;
      VIA 82.8 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 157.595 83.59 157.925 ;
      VIA 82.8 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 157.575 83.57 157.945 ;
      VIA 82.8 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 152.155 83.59 152.485 ;
      VIA 82.8 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 152.135 83.57 152.505 ;
      VIA 82.8 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 146.715 83.59 147.045 ;
      VIA 82.8 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 146.695 83.57 147.065 ;
      VIA 82.8 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 141.275 83.59 141.605 ;
      VIA 82.8 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 141.255 83.57 141.625 ;
      VIA 82.8 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 135.835 83.59 136.165 ;
      VIA 82.8 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 135.815 83.57 136.185 ;
      VIA 82.8 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 130.395 83.59 130.725 ;
      VIA 82.8 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 130.375 83.57 130.745 ;
      VIA 82.8 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 124.955 83.59 125.285 ;
      VIA 82.8 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 124.935 83.57 125.305 ;
      VIA 82.8 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 119.515 83.59 119.845 ;
      VIA 82.8 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 119.495 83.57 119.865 ;
      VIA 82.8 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 114.075 83.59 114.405 ;
      VIA 82.8 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 114.055 83.57 114.425 ;
      VIA 82.8 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 108.635 83.59 108.965 ;
      VIA 82.8 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 108.615 83.57 108.985 ;
      VIA 82.8 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 103.195 83.59 103.525 ;
      VIA 82.8 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 103.175 83.57 103.545 ;
      VIA 82.8 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 97.755 83.59 98.085 ;
      VIA 82.8 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 97.735 83.57 98.105 ;
      VIA 82.8 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 92.315 83.59 92.645 ;
      VIA 82.8 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 92.295 83.57 92.665 ;
      VIA 82.8 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 86.875 83.59 87.205 ;
      VIA 82.8 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 86.855 83.57 87.225 ;
      VIA 82.8 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 81.435 83.59 81.765 ;
      VIA 82.8 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 81.415 83.57 81.785 ;
      VIA 82.8 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 75.995 83.59 76.325 ;
      VIA 82.8 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 75.975 83.57 76.345 ;
      VIA 82.8 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 70.555 83.59 70.885 ;
      VIA 82.8 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 70.535 83.57 70.905 ;
      VIA 82.8 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 65.115 83.59 65.445 ;
      VIA 82.8 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 65.095 83.57 65.465 ;
      VIA 82.8 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 59.675 83.59 60.005 ;
      VIA 82.8 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 59.655 83.57 60.025 ;
      VIA 82.8 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 54.235 83.59 54.565 ;
      VIA 82.8 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 54.215 83.57 54.585 ;
      VIA 82.8 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 48.795 83.59 49.125 ;
      VIA 82.8 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 48.775 83.57 49.145 ;
      VIA 82.8 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 43.355 83.59 43.685 ;
      VIA 82.8 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 43.335 83.57 43.705 ;
      VIA 82.8 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 37.915 83.59 38.245 ;
      VIA 82.8 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 37.895 83.57 38.265 ;
      VIA 82.8 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 32.475 83.59 32.805 ;
      VIA 82.8 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 32.455 83.57 32.825 ;
      VIA 82.8 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 27.035 83.59 27.365 ;
      VIA 82.8 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 27.015 83.57 27.385 ;
      VIA 82.8 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 21.595 83.59 21.925 ;
      VIA 82.8 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 21.575 83.57 21.945 ;
      VIA 82.8 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 16.155 83.59 16.485 ;
      VIA 82.8 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 16.135 83.57 16.505 ;
      VIA 82.8 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 10.715 83.59 11.045 ;
      VIA 82.8 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 10.695 83.57 11.065 ;
      VIA 82.8 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 5.275 83.59 5.605 ;
      VIA 82.8 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 5.255 83.57 5.625 ;
      VIA 82.8 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 293.595 56.45 293.925 ;
      VIA 55.66 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 293.575 56.43 293.945 ;
      VIA 55.66 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 288.155 56.45 288.485 ;
      VIA 55.66 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 288.135 56.43 288.505 ;
      VIA 55.66 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 282.715 56.45 283.045 ;
      VIA 55.66 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 282.695 56.43 283.065 ;
      VIA 55.66 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 277.275 56.45 277.605 ;
      VIA 55.66 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 277.255 56.43 277.625 ;
      VIA 55.66 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 271.835 56.45 272.165 ;
      VIA 55.66 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 271.815 56.43 272.185 ;
      VIA 55.66 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 266.395 56.45 266.725 ;
      VIA 55.66 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 266.375 56.43 266.745 ;
      VIA 55.66 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 260.955 56.45 261.285 ;
      VIA 55.66 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 260.935 56.43 261.305 ;
      VIA 55.66 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 255.515 56.45 255.845 ;
      VIA 55.66 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 255.495 56.43 255.865 ;
      VIA 55.66 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 250.075 56.45 250.405 ;
      VIA 55.66 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 250.055 56.43 250.425 ;
      VIA 55.66 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 244.635 56.45 244.965 ;
      VIA 55.66 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 244.615 56.43 244.985 ;
      VIA 55.66 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 239.195 56.45 239.525 ;
      VIA 55.66 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 239.175 56.43 239.545 ;
      VIA 55.66 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 233.755 56.45 234.085 ;
      VIA 55.66 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 233.735 56.43 234.105 ;
      VIA 55.66 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 228.315 56.45 228.645 ;
      VIA 55.66 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 228.295 56.43 228.665 ;
      VIA 55.66 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 222.875 56.45 223.205 ;
      VIA 55.66 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 222.855 56.43 223.225 ;
      VIA 55.66 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 217.435 56.45 217.765 ;
      VIA 55.66 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 217.415 56.43 217.785 ;
      VIA 55.66 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 211.995 56.45 212.325 ;
      VIA 55.66 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 211.975 56.43 212.345 ;
      VIA 55.66 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 206.555 56.45 206.885 ;
      VIA 55.66 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 206.535 56.43 206.905 ;
      VIA 55.66 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 201.115 56.45 201.445 ;
      VIA 55.66 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 201.095 56.43 201.465 ;
      VIA 55.66 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 195.675 56.45 196.005 ;
      VIA 55.66 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 195.655 56.43 196.025 ;
      VIA 55.66 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 190.235 56.45 190.565 ;
      VIA 55.66 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 190.215 56.43 190.585 ;
      VIA 55.66 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 184.795 56.45 185.125 ;
      VIA 55.66 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 184.775 56.43 185.145 ;
      VIA 55.66 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 179.355 56.45 179.685 ;
      VIA 55.66 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 179.335 56.43 179.705 ;
      VIA 55.66 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 173.915 56.45 174.245 ;
      VIA 55.66 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 173.895 56.43 174.265 ;
      VIA 55.66 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 168.475 56.45 168.805 ;
      VIA 55.66 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 168.455 56.43 168.825 ;
      VIA 55.66 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 163.035 56.45 163.365 ;
      VIA 55.66 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 163.015 56.43 163.385 ;
      VIA 55.66 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 157.595 56.45 157.925 ;
      VIA 55.66 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 157.575 56.43 157.945 ;
      VIA 55.66 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 152.155 56.45 152.485 ;
      VIA 55.66 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 152.135 56.43 152.505 ;
      VIA 55.66 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 146.715 56.45 147.045 ;
      VIA 55.66 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 146.695 56.43 147.065 ;
      VIA 55.66 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 141.275 56.45 141.605 ;
      VIA 55.66 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 141.255 56.43 141.625 ;
      VIA 55.66 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 135.835 56.45 136.165 ;
      VIA 55.66 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 135.815 56.43 136.185 ;
      VIA 55.66 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 130.395 56.45 130.725 ;
      VIA 55.66 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 130.375 56.43 130.745 ;
      VIA 55.66 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 124.955 56.45 125.285 ;
      VIA 55.66 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 124.935 56.43 125.305 ;
      VIA 55.66 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 119.515 56.45 119.845 ;
      VIA 55.66 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 119.495 56.43 119.865 ;
      VIA 55.66 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 114.075 56.45 114.405 ;
      VIA 55.66 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 114.055 56.43 114.425 ;
      VIA 55.66 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 108.635 56.45 108.965 ;
      VIA 55.66 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 108.615 56.43 108.985 ;
      VIA 55.66 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 103.195 56.45 103.525 ;
      VIA 55.66 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 103.175 56.43 103.545 ;
      VIA 55.66 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 97.755 56.45 98.085 ;
      VIA 55.66 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 97.735 56.43 98.105 ;
      VIA 55.66 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 92.315 56.45 92.645 ;
      VIA 55.66 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 92.295 56.43 92.665 ;
      VIA 55.66 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 86.875 56.45 87.205 ;
      VIA 55.66 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 86.855 56.43 87.225 ;
      VIA 55.66 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 81.435 56.45 81.765 ;
      VIA 55.66 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 81.415 56.43 81.785 ;
      VIA 55.66 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 75.995 56.45 76.325 ;
      VIA 55.66 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 75.975 56.43 76.345 ;
      VIA 55.66 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 70.555 56.45 70.885 ;
      VIA 55.66 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 70.535 56.43 70.905 ;
      VIA 55.66 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 65.115 56.45 65.445 ;
      VIA 55.66 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 65.095 56.43 65.465 ;
      VIA 55.66 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 59.675 56.45 60.005 ;
      VIA 55.66 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 59.655 56.43 60.025 ;
      VIA 55.66 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 54.235 56.45 54.565 ;
      VIA 55.66 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 54.215 56.43 54.585 ;
      VIA 55.66 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 48.795 56.45 49.125 ;
      VIA 55.66 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 48.775 56.43 49.145 ;
      VIA 55.66 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 43.355 56.45 43.685 ;
      VIA 55.66 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 43.335 56.43 43.705 ;
      VIA 55.66 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 37.915 56.45 38.245 ;
      VIA 55.66 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 37.895 56.43 38.265 ;
      VIA 55.66 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 32.475 56.45 32.805 ;
      VIA 55.66 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 32.455 56.43 32.825 ;
      VIA 55.66 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 27.035 56.45 27.365 ;
      VIA 55.66 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 27.015 56.43 27.385 ;
      VIA 55.66 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 21.595 56.45 21.925 ;
      VIA 55.66 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 21.575 56.43 21.945 ;
      VIA 55.66 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 16.155 56.45 16.485 ;
      VIA 55.66 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 16.135 56.43 16.505 ;
      VIA 55.66 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 10.715 56.45 11.045 ;
      VIA 55.66 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 10.695 56.43 11.065 ;
      VIA 55.66 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 5.275 56.45 5.605 ;
      VIA 55.66 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 5.255 56.43 5.625 ;
      VIA 55.66 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 293.595 29.31 293.925 ;
      VIA 28.52 293.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 293.575 29.29 293.945 ;
      VIA 28.52 293.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 293.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 288.155 29.31 288.485 ;
      VIA 28.52 288.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 288.135 29.29 288.505 ;
      VIA 28.52 288.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 288.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 282.715 29.31 283.045 ;
      VIA 28.52 282.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 282.695 29.29 283.065 ;
      VIA 28.52 282.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 282.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 277.275 29.31 277.605 ;
      VIA 28.52 277.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 277.255 29.29 277.625 ;
      VIA 28.52 277.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 277.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 271.835 29.31 272.165 ;
      VIA 28.52 272 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 271.815 29.29 272.185 ;
      VIA 28.52 272 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 272 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 266.395 29.31 266.725 ;
      VIA 28.52 266.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 266.375 29.29 266.745 ;
      VIA 28.52 266.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 266.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 260.955 29.31 261.285 ;
      VIA 28.52 261.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 260.935 29.29 261.305 ;
      VIA 28.52 261.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 261.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 255.515 29.31 255.845 ;
      VIA 28.52 255.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 255.495 29.29 255.865 ;
      VIA 28.52 255.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 255.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 250.075 29.31 250.405 ;
      VIA 28.52 250.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 250.055 29.29 250.425 ;
      VIA 28.52 250.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 250.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 244.635 29.31 244.965 ;
      VIA 28.52 244.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 244.615 29.29 244.985 ;
      VIA 28.52 244.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 244.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 239.195 29.31 239.525 ;
      VIA 28.52 239.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 239.175 29.29 239.545 ;
      VIA 28.52 239.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 239.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 233.755 29.31 234.085 ;
      VIA 28.52 233.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 233.735 29.29 234.105 ;
      VIA 28.52 233.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 233.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 228.315 29.31 228.645 ;
      VIA 28.52 228.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 228.295 29.29 228.665 ;
      VIA 28.52 228.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 228.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 222.875 29.31 223.205 ;
      VIA 28.52 223.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 222.855 29.29 223.225 ;
      VIA 28.52 223.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 223.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 217.435 29.31 217.765 ;
      VIA 28.52 217.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 217.415 29.29 217.785 ;
      VIA 28.52 217.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 217.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 211.995 29.31 212.325 ;
      VIA 28.52 212.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 211.975 29.29 212.345 ;
      VIA 28.52 212.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 212.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 206.555 29.31 206.885 ;
      VIA 28.52 206.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 206.535 29.29 206.905 ;
      VIA 28.52 206.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 206.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 201.115 29.31 201.445 ;
      VIA 28.52 201.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 201.095 29.29 201.465 ;
      VIA 28.52 201.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 201.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 195.675 29.31 196.005 ;
      VIA 28.52 195.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 195.655 29.29 196.025 ;
      VIA 28.52 195.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 195.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 190.235 29.31 190.565 ;
      VIA 28.52 190.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 190.215 29.29 190.585 ;
      VIA 28.52 190.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 190.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 184.795 29.31 185.125 ;
      VIA 28.52 184.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 184.775 29.29 185.145 ;
      VIA 28.52 184.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 184.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 179.355 29.31 179.685 ;
      VIA 28.52 179.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 179.335 29.29 179.705 ;
      VIA 28.52 179.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 179.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 173.915 29.31 174.245 ;
      VIA 28.52 174.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 173.895 29.29 174.265 ;
      VIA 28.52 174.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 174.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 168.475 29.31 168.805 ;
      VIA 28.52 168.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 168.455 29.29 168.825 ;
      VIA 28.52 168.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 168.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 163.035 29.31 163.365 ;
      VIA 28.52 163.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 163.015 29.29 163.385 ;
      VIA 28.52 163.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 163.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 157.595 29.31 157.925 ;
      VIA 28.52 157.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 157.575 29.29 157.945 ;
      VIA 28.52 157.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 157.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 152.155 29.31 152.485 ;
      VIA 28.52 152.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 152.135 29.29 152.505 ;
      VIA 28.52 152.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 152.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 146.715 29.31 147.045 ;
      VIA 28.52 146.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 146.695 29.29 147.065 ;
      VIA 28.52 146.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 146.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 141.275 29.31 141.605 ;
      VIA 28.52 141.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 141.255 29.29 141.625 ;
      VIA 28.52 141.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 141.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 135.835 29.31 136.165 ;
      VIA 28.52 136 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 135.815 29.29 136.185 ;
      VIA 28.52 136 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 136 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 130.395 29.31 130.725 ;
      VIA 28.52 130.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 130.375 29.29 130.745 ;
      VIA 28.52 130.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 130.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 124.955 29.31 125.285 ;
      VIA 28.52 125.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 124.935 29.29 125.305 ;
      VIA 28.52 125.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 125.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 119.515 29.31 119.845 ;
      VIA 28.52 119.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 119.495 29.29 119.865 ;
      VIA 28.52 119.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 119.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 114.075 29.31 114.405 ;
      VIA 28.52 114.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 114.055 29.29 114.425 ;
      VIA 28.52 114.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 114.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 108.635 29.31 108.965 ;
      VIA 28.52 108.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 108.615 29.29 108.985 ;
      VIA 28.52 108.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 108.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 103.195 29.31 103.525 ;
      VIA 28.52 103.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 103.175 29.29 103.545 ;
      VIA 28.52 103.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 103.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 97.755 29.31 98.085 ;
      VIA 28.52 97.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 97.735 29.29 98.105 ;
      VIA 28.52 97.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 97.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 92.315 29.31 92.645 ;
      VIA 28.52 92.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 92.295 29.29 92.665 ;
      VIA 28.52 92.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 92.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 86.875 29.31 87.205 ;
      VIA 28.52 87.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 86.855 29.29 87.225 ;
      VIA 28.52 87.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 87.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 81.435 29.31 81.765 ;
      VIA 28.52 81.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 81.415 29.29 81.785 ;
      VIA 28.52 81.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 81.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 75.995 29.31 76.325 ;
      VIA 28.52 76.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 75.975 29.29 76.345 ;
      VIA 28.52 76.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 76.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 70.555 29.31 70.885 ;
      VIA 28.52 70.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 70.535 29.29 70.905 ;
      VIA 28.52 70.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 70.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 65.115 29.31 65.445 ;
      VIA 28.52 65.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 65.095 29.29 65.465 ;
      VIA 28.52 65.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 65.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 59.675 29.31 60.005 ;
      VIA 28.52 59.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 59.655 29.29 60.025 ;
      VIA 28.52 59.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 59.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 54.235 29.31 54.565 ;
      VIA 28.52 54.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 54.215 29.29 54.585 ;
      VIA 28.52 54.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 54.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 48.795 29.31 49.125 ;
      VIA 28.52 48.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 48.775 29.29 49.145 ;
      VIA 28.52 48.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 48.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 43.355 29.31 43.685 ;
      VIA 28.52 43.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 43.335 29.29 43.705 ;
      VIA 28.52 43.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 43.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 37.915 29.31 38.245 ;
      VIA 28.52 38.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 37.895 29.29 38.265 ;
      VIA 28.52 38.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 38.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 32.475 29.31 32.805 ;
      VIA 28.52 32.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 32.455 29.29 32.825 ;
      VIA 28.52 32.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 32.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 27.035 29.31 27.365 ;
      VIA 28.52 27.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 27.015 29.29 27.385 ;
      VIA 28.52 27.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 27.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 21.595 29.31 21.925 ;
      VIA 28.52 21.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 21.575 29.29 21.945 ;
      VIA 28.52 21.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 21.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 16.155 29.31 16.485 ;
      VIA 28.52 16.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 16.135 29.29 16.505 ;
      VIA 28.52 16.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 16.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 10.715 29.31 11.045 ;
      VIA 28.52 10.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 10.695 29.29 11.065 ;
      VIA 28.52 10.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 10.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 5.275 29.31 5.605 ;
      VIA 28.52 5.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 5.255 29.29 5.625 ;
      VIA 28.52 5.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 5.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  14.15 287.52 287.15 289.12 ;
        RECT  14.15 260.32 287.15 261.92 ;
        RECT  14.15 233.12 287.15 234.72 ;
        RECT  14.15 205.92 287.15 207.52 ;
        RECT  14.15 178.72 287.15 180.32 ;
        RECT  14.15 151.52 287.15 153.12 ;
        RECT  14.15 124.32 287.15 125.92 ;
        RECT  14.15 97.12 287.15 98.72 ;
        RECT  14.15 69.92 287.15 71.52 ;
        RECT  14.15 42.72 287.15 44.32 ;
        RECT  14.15 15.52 287.15 17.12 ;
      LAYER met4 ;
        RECT  285.55 2.48 287.15 291.28 ;
        RECT  258.41 2.48 260.01 291.28 ;
        RECT  231.27 2.48 232.87 291.28 ;
        RECT  204.13 2.48 205.73 291.28 ;
        RECT  176.99 2.48 178.59 291.28 ;
        RECT  149.85 2.48 151.45 291.28 ;
        RECT  122.71 2.48 124.31 291.28 ;
        RECT  95.57 2.48 97.17 291.28 ;
        RECT  68.43 2.48 70.03 291.28 ;
        RECT  41.29 2.48 42.89 291.28 ;
        RECT  14.15 2.48 15.75 291.28 ;
      LAYER met1 ;
        RECT  1.38 290.8 294.86 291.28 ;
        RECT  1.38 285.36 294.86 285.84 ;
        RECT  1.38 279.92 294.86 280.4 ;
        RECT  1.38 274.48 294.86 274.96 ;
        RECT  1.38 269.04 294.86 269.52 ;
        RECT  1.38 263.6 294.86 264.08 ;
        RECT  1.38 258.16 294.86 258.64 ;
        RECT  1.38 252.72 294.86 253.2 ;
        RECT  1.38 247.28 294.86 247.76 ;
        RECT  1.38 241.84 294.86 242.32 ;
        RECT  1.38 236.4 294.86 236.88 ;
        RECT  1.38 230.96 294.86 231.44 ;
        RECT  1.38 225.52 294.86 226 ;
        RECT  1.38 220.08 294.86 220.56 ;
        RECT  1.38 214.64 294.86 215.12 ;
        RECT  1.38 209.2 294.86 209.68 ;
        RECT  1.38 203.76 294.86 204.24 ;
        RECT  1.38 198.32 294.86 198.8 ;
        RECT  1.38 192.88 294.86 193.36 ;
        RECT  1.38 187.44 294.86 187.92 ;
        RECT  1.38 182 294.86 182.48 ;
        RECT  1.38 176.56 294.86 177.04 ;
        RECT  1.38 171.12 294.86 171.6 ;
        RECT  1.38 165.68 294.86 166.16 ;
        RECT  1.38 160.24 294.86 160.72 ;
        RECT  1.38 154.8 294.86 155.28 ;
        RECT  1.38 149.36 294.86 149.84 ;
        RECT  1.38 143.92 294.86 144.4 ;
        RECT  1.38 138.48 294.86 138.96 ;
        RECT  1.38 133.04 294.86 133.52 ;
        RECT  1.38 127.6 294.86 128.08 ;
        RECT  1.38 122.16 294.86 122.64 ;
        RECT  1.38 116.72 294.86 117.2 ;
        RECT  1.38 111.28 294.86 111.76 ;
        RECT  1.38 105.84 294.86 106.32 ;
        RECT  1.38 100.4 294.86 100.88 ;
        RECT  1.38 94.96 294.86 95.44 ;
        RECT  1.38 89.52 294.86 90 ;
        RECT  1.38 84.08 294.86 84.56 ;
        RECT  1.38 78.64 294.86 79.12 ;
        RECT  1.38 73.2 294.86 73.68 ;
        RECT  1.38 67.76 294.86 68.24 ;
        RECT  1.38 62.32 294.86 62.8 ;
        RECT  1.38 56.88 294.86 57.36 ;
        RECT  1.38 51.44 294.86 51.92 ;
        RECT  1.38 46 294.86 46.48 ;
        RECT  1.38 40.56 294.86 41.04 ;
        RECT  1.38 35.12 294.86 35.6 ;
        RECT  1.38 29.68 294.86 30.16 ;
        RECT  1.38 24.24 294.86 24.72 ;
        RECT  1.38 18.8 294.86 19.28 ;
        RECT  1.38 13.36 294.86 13.84 ;
        RECT  1.38 7.92 294.86 8.4 ;
        RECT  1.38 2.48 294.86 2.96 ;
      VIA 286.35 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 286.35 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.21 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.07 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.93 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.79 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 288.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 261.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 233.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 206.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 179.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 152.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 125.12 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 97.92 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 70.72 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 43.52 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 16.32 ibex_if_stage_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  285.56 290.875 287.14 291.205 ;
      VIA 286.35 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 290.855 287.12 291.225 ;
      VIA 286.35 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 285.435 287.14 285.765 ;
      VIA 286.35 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 285.415 287.12 285.785 ;
      VIA 286.35 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 279.995 287.14 280.325 ;
      VIA 286.35 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 279.975 287.12 280.345 ;
      VIA 286.35 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 274.555 287.14 274.885 ;
      VIA 286.35 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 274.535 287.12 274.905 ;
      VIA 286.35 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 269.115 287.14 269.445 ;
      VIA 286.35 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 269.095 287.12 269.465 ;
      VIA 286.35 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 263.675 287.14 264.005 ;
      VIA 286.35 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 263.655 287.12 264.025 ;
      VIA 286.35 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 258.235 287.14 258.565 ;
      VIA 286.35 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 258.215 287.12 258.585 ;
      VIA 286.35 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 252.795 287.14 253.125 ;
      VIA 286.35 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 252.775 287.12 253.145 ;
      VIA 286.35 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 247.355 287.14 247.685 ;
      VIA 286.35 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 247.335 287.12 247.705 ;
      VIA 286.35 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 241.915 287.14 242.245 ;
      VIA 286.35 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 241.895 287.12 242.265 ;
      VIA 286.35 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 236.475 287.14 236.805 ;
      VIA 286.35 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 236.455 287.12 236.825 ;
      VIA 286.35 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 231.035 287.14 231.365 ;
      VIA 286.35 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 231.015 287.12 231.385 ;
      VIA 286.35 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 225.595 287.14 225.925 ;
      VIA 286.35 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 225.575 287.12 225.945 ;
      VIA 286.35 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 220.155 287.14 220.485 ;
      VIA 286.35 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 220.135 287.12 220.505 ;
      VIA 286.35 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 214.715 287.14 215.045 ;
      VIA 286.35 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 214.695 287.12 215.065 ;
      VIA 286.35 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 209.275 287.14 209.605 ;
      VIA 286.35 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 209.255 287.12 209.625 ;
      VIA 286.35 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 203.835 287.14 204.165 ;
      VIA 286.35 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 203.815 287.12 204.185 ;
      VIA 286.35 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 198.395 287.14 198.725 ;
      VIA 286.35 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 198.375 287.12 198.745 ;
      VIA 286.35 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 192.955 287.14 193.285 ;
      VIA 286.35 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 192.935 287.12 193.305 ;
      VIA 286.35 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 187.515 287.14 187.845 ;
      VIA 286.35 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 187.495 287.12 187.865 ;
      VIA 286.35 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 182.075 287.14 182.405 ;
      VIA 286.35 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 182.055 287.12 182.425 ;
      VIA 286.35 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 176.635 287.14 176.965 ;
      VIA 286.35 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 176.615 287.12 176.985 ;
      VIA 286.35 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 171.195 287.14 171.525 ;
      VIA 286.35 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 171.175 287.12 171.545 ;
      VIA 286.35 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 165.755 287.14 166.085 ;
      VIA 286.35 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 165.735 287.12 166.105 ;
      VIA 286.35 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 160.315 287.14 160.645 ;
      VIA 286.35 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 160.295 287.12 160.665 ;
      VIA 286.35 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 154.875 287.14 155.205 ;
      VIA 286.35 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 154.855 287.12 155.225 ;
      VIA 286.35 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 149.435 287.14 149.765 ;
      VIA 286.35 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 149.415 287.12 149.785 ;
      VIA 286.35 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 143.995 287.14 144.325 ;
      VIA 286.35 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 143.975 287.12 144.345 ;
      VIA 286.35 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 138.555 287.14 138.885 ;
      VIA 286.35 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 138.535 287.12 138.905 ;
      VIA 286.35 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 133.115 287.14 133.445 ;
      VIA 286.35 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 133.095 287.12 133.465 ;
      VIA 286.35 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 127.675 287.14 128.005 ;
      VIA 286.35 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 127.655 287.12 128.025 ;
      VIA 286.35 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 122.235 287.14 122.565 ;
      VIA 286.35 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 122.215 287.12 122.585 ;
      VIA 286.35 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 116.795 287.14 117.125 ;
      VIA 286.35 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 116.775 287.12 117.145 ;
      VIA 286.35 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 111.355 287.14 111.685 ;
      VIA 286.35 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 111.335 287.12 111.705 ;
      VIA 286.35 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 105.915 287.14 106.245 ;
      VIA 286.35 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 105.895 287.12 106.265 ;
      VIA 286.35 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 100.475 287.14 100.805 ;
      VIA 286.35 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 100.455 287.12 100.825 ;
      VIA 286.35 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 95.035 287.14 95.365 ;
      VIA 286.35 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 95.015 287.12 95.385 ;
      VIA 286.35 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 89.595 287.14 89.925 ;
      VIA 286.35 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 89.575 287.12 89.945 ;
      VIA 286.35 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 84.155 287.14 84.485 ;
      VIA 286.35 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 84.135 287.12 84.505 ;
      VIA 286.35 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 78.715 287.14 79.045 ;
      VIA 286.35 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 78.695 287.12 79.065 ;
      VIA 286.35 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 73.275 287.14 73.605 ;
      VIA 286.35 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 73.255 287.12 73.625 ;
      VIA 286.35 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 67.835 287.14 68.165 ;
      VIA 286.35 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 67.815 287.12 68.185 ;
      VIA 286.35 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 62.395 287.14 62.725 ;
      VIA 286.35 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 62.375 287.12 62.745 ;
      VIA 286.35 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 56.955 287.14 57.285 ;
      VIA 286.35 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 56.935 287.12 57.305 ;
      VIA 286.35 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 51.515 287.14 51.845 ;
      VIA 286.35 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 51.495 287.12 51.865 ;
      VIA 286.35 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 46.075 287.14 46.405 ;
      VIA 286.35 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 46.055 287.12 46.425 ;
      VIA 286.35 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 40.635 287.14 40.965 ;
      VIA 286.35 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 40.615 287.12 40.985 ;
      VIA 286.35 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 35.195 287.14 35.525 ;
      VIA 286.35 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 35.175 287.12 35.545 ;
      VIA 286.35 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 29.755 287.14 30.085 ;
      VIA 286.35 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 29.735 287.12 30.105 ;
      VIA 286.35 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 24.315 287.14 24.645 ;
      VIA 286.35 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 24.295 287.12 24.665 ;
      VIA 286.35 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 18.875 287.14 19.205 ;
      VIA 286.35 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 18.855 287.12 19.225 ;
      VIA 286.35 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 13.435 287.14 13.765 ;
      VIA 286.35 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 13.415 287.12 13.785 ;
      VIA 286.35 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 7.995 287.14 8.325 ;
      VIA 286.35 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 7.975 287.12 8.345 ;
      VIA 286.35 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  285.56 2.555 287.14 2.885 ;
      VIA 286.35 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  285.58 2.535 287.12 2.905 ;
      VIA 286.35 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 286.35 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 290.875 260 291.205 ;
      VIA 259.21 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 290.855 259.98 291.225 ;
      VIA 259.21 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 285.435 260 285.765 ;
      VIA 259.21 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 285.415 259.98 285.785 ;
      VIA 259.21 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 279.995 260 280.325 ;
      VIA 259.21 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 279.975 259.98 280.345 ;
      VIA 259.21 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 274.555 260 274.885 ;
      VIA 259.21 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 274.535 259.98 274.905 ;
      VIA 259.21 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 269.115 260 269.445 ;
      VIA 259.21 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 269.095 259.98 269.465 ;
      VIA 259.21 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 263.675 260 264.005 ;
      VIA 259.21 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 263.655 259.98 264.025 ;
      VIA 259.21 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 258.235 260 258.565 ;
      VIA 259.21 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 258.215 259.98 258.585 ;
      VIA 259.21 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 252.795 260 253.125 ;
      VIA 259.21 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 252.775 259.98 253.145 ;
      VIA 259.21 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 247.355 260 247.685 ;
      VIA 259.21 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 247.335 259.98 247.705 ;
      VIA 259.21 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 241.915 260 242.245 ;
      VIA 259.21 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 241.895 259.98 242.265 ;
      VIA 259.21 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 236.475 260 236.805 ;
      VIA 259.21 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 236.455 259.98 236.825 ;
      VIA 259.21 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 231.035 260 231.365 ;
      VIA 259.21 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 231.015 259.98 231.385 ;
      VIA 259.21 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 225.595 260 225.925 ;
      VIA 259.21 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 225.575 259.98 225.945 ;
      VIA 259.21 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 220.155 260 220.485 ;
      VIA 259.21 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 220.135 259.98 220.505 ;
      VIA 259.21 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 214.715 260 215.045 ;
      VIA 259.21 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 214.695 259.98 215.065 ;
      VIA 259.21 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 209.275 260 209.605 ;
      VIA 259.21 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 209.255 259.98 209.625 ;
      VIA 259.21 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 203.835 260 204.165 ;
      VIA 259.21 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 203.815 259.98 204.185 ;
      VIA 259.21 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 198.395 260 198.725 ;
      VIA 259.21 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 198.375 259.98 198.745 ;
      VIA 259.21 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 192.955 260 193.285 ;
      VIA 259.21 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 192.935 259.98 193.305 ;
      VIA 259.21 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 187.515 260 187.845 ;
      VIA 259.21 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 187.495 259.98 187.865 ;
      VIA 259.21 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 182.075 260 182.405 ;
      VIA 259.21 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 182.055 259.98 182.425 ;
      VIA 259.21 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 176.635 260 176.965 ;
      VIA 259.21 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 176.615 259.98 176.985 ;
      VIA 259.21 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 171.195 260 171.525 ;
      VIA 259.21 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 171.175 259.98 171.545 ;
      VIA 259.21 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 165.755 260 166.085 ;
      VIA 259.21 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 165.735 259.98 166.105 ;
      VIA 259.21 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 160.315 260 160.645 ;
      VIA 259.21 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 160.295 259.98 160.665 ;
      VIA 259.21 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 154.875 260 155.205 ;
      VIA 259.21 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 154.855 259.98 155.225 ;
      VIA 259.21 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 149.435 260 149.765 ;
      VIA 259.21 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 149.415 259.98 149.785 ;
      VIA 259.21 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 143.995 260 144.325 ;
      VIA 259.21 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 143.975 259.98 144.345 ;
      VIA 259.21 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 138.555 260 138.885 ;
      VIA 259.21 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 138.535 259.98 138.905 ;
      VIA 259.21 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 133.115 260 133.445 ;
      VIA 259.21 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 133.095 259.98 133.465 ;
      VIA 259.21 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 127.675 260 128.005 ;
      VIA 259.21 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 127.655 259.98 128.025 ;
      VIA 259.21 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 122.235 260 122.565 ;
      VIA 259.21 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 122.215 259.98 122.585 ;
      VIA 259.21 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 116.795 260 117.125 ;
      VIA 259.21 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 116.775 259.98 117.145 ;
      VIA 259.21 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 111.355 260 111.685 ;
      VIA 259.21 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 111.335 259.98 111.705 ;
      VIA 259.21 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 105.915 260 106.245 ;
      VIA 259.21 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 105.895 259.98 106.265 ;
      VIA 259.21 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 100.475 260 100.805 ;
      VIA 259.21 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 100.455 259.98 100.825 ;
      VIA 259.21 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 95.035 260 95.365 ;
      VIA 259.21 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 95.015 259.98 95.385 ;
      VIA 259.21 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 89.595 260 89.925 ;
      VIA 259.21 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 89.575 259.98 89.945 ;
      VIA 259.21 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 84.155 260 84.485 ;
      VIA 259.21 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 84.135 259.98 84.505 ;
      VIA 259.21 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 78.715 260 79.045 ;
      VIA 259.21 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 78.695 259.98 79.065 ;
      VIA 259.21 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 73.275 260 73.605 ;
      VIA 259.21 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 73.255 259.98 73.625 ;
      VIA 259.21 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 67.835 260 68.165 ;
      VIA 259.21 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 67.815 259.98 68.185 ;
      VIA 259.21 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 62.395 260 62.725 ;
      VIA 259.21 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 62.375 259.98 62.745 ;
      VIA 259.21 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 56.955 260 57.285 ;
      VIA 259.21 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 56.935 259.98 57.305 ;
      VIA 259.21 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 51.515 260 51.845 ;
      VIA 259.21 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 51.495 259.98 51.865 ;
      VIA 259.21 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 46.075 260 46.405 ;
      VIA 259.21 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 46.055 259.98 46.425 ;
      VIA 259.21 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 40.635 260 40.965 ;
      VIA 259.21 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 40.615 259.98 40.985 ;
      VIA 259.21 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 35.195 260 35.525 ;
      VIA 259.21 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 35.175 259.98 35.545 ;
      VIA 259.21 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 29.755 260 30.085 ;
      VIA 259.21 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 29.735 259.98 30.105 ;
      VIA 259.21 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 24.315 260 24.645 ;
      VIA 259.21 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 24.295 259.98 24.665 ;
      VIA 259.21 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 18.875 260 19.205 ;
      VIA 259.21 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 18.855 259.98 19.225 ;
      VIA 259.21 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 13.435 260 13.765 ;
      VIA 259.21 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 13.415 259.98 13.785 ;
      VIA 259.21 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 7.995 260 8.325 ;
      VIA 259.21 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 7.975 259.98 8.345 ;
      VIA 259.21 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.42 2.555 260 2.885 ;
      VIA 259.21 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.44 2.535 259.98 2.905 ;
      VIA 259.21 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 259.21 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 290.875 232.86 291.205 ;
      VIA 232.07 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 290.855 232.84 291.225 ;
      VIA 232.07 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 285.435 232.86 285.765 ;
      VIA 232.07 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 285.415 232.84 285.785 ;
      VIA 232.07 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 279.995 232.86 280.325 ;
      VIA 232.07 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 279.975 232.84 280.345 ;
      VIA 232.07 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 274.555 232.86 274.885 ;
      VIA 232.07 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 274.535 232.84 274.905 ;
      VIA 232.07 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 269.115 232.86 269.445 ;
      VIA 232.07 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 269.095 232.84 269.465 ;
      VIA 232.07 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 263.675 232.86 264.005 ;
      VIA 232.07 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 263.655 232.84 264.025 ;
      VIA 232.07 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 258.235 232.86 258.565 ;
      VIA 232.07 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 258.215 232.84 258.585 ;
      VIA 232.07 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 252.795 232.86 253.125 ;
      VIA 232.07 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 252.775 232.84 253.145 ;
      VIA 232.07 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 247.355 232.86 247.685 ;
      VIA 232.07 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 247.335 232.84 247.705 ;
      VIA 232.07 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 241.915 232.86 242.245 ;
      VIA 232.07 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 241.895 232.84 242.265 ;
      VIA 232.07 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 236.475 232.86 236.805 ;
      VIA 232.07 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 236.455 232.84 236.825 ;
      VIA 232.07 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 231.035 232.86 231.365 ;
      VIA 232.07 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 231.015 232.84 231.385 ;
      VIA 232.07 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 225.595 232.86 225.925 ;
      VIA 232.07 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 225.575 232.84 225.945 ;
      VIA 232.07 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 220.155 232.86 220.485 ;
      VIA 232.07 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 220.135 232.84 220.505 ;
      VIA 232.07 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 214.715 232.86 215.045 ;
      VIA 232.07 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 214.695 232.84 215.065 ;
      VIA 232.07 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 209.275 232.86 209.605 ;
      VIA 232.07 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 209.255 232.84 209.625 ;
      VIA 232.07 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 203.835 232.86 204.165 ;
      VIA 232.07 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 203.815 232.84 204.185 ;
      VIA 232.07 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 198.395 232.86 198.725 ;
      VIA 232.07 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 198.375 232.84 198.745 ;
      VIA 232.07 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 192.955 232.86 193.285 ;
      VIA 232.07 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 192.935 232.84 193.305 ;
      VIA 232.07 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 187.515 232.86 187.845 ;
      VIA 232.07 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 187.495 232.84 187.865 ;
      VIA 232.07 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 182.075 232.86 182.405 ;
      VIA 232.07 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 182.055 232.84 182.425 ;
      VIA 232.07 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 176.635 232.86 176.965 ;
      VIA 232.07 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 176.615 232.84 176.985 ;
      VIA 232.07 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 171.195 232.86 171.525 ;
      VIA 232.07 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 171.175 232.84 171.545 ;
      VIA 232.07 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 165.755 232.86 166.085 ;
      VIA 232.07 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 165.735 232.84 166.105 ;
      VIA 232.07 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 160.315 232.86 160.645 ;
      VIA 232.07 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 160.295 232.84 160.665 ;
      VIA 232.07 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 154.875 232.86 155.205 ;
      VIA 232.07 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 154.855 232.84 155.225 ;
      VIA 232.07 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 149.435 232.86 149.765 ;
      VIA 232.07 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 149.415 232.84 149.785 ;
      VIA 232.07 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 143.995 232.86 144.325 ;
      VIA 232.07 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 143.975 232.84 144.345 ;
      VIA 232.07 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 138.555 232.86 138.885 ;
      VIA 232.07 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 138.535 232.84 138.905 ;
      VIA 232.07 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 133.115 232.86 133.445 ;
      VIA 232.07 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 133.095 232.84 133.465 ;
      VIA 232.07 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 127.675 232.86 128.005 ;
      VIA 232.07 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 127.655 232.84 128.025 ;
      VIA 232.07 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 122.235 232.86 122.565 ;
      VIA 232.07 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 122.215 232.84 122.585 ;
      VIA 232.07 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 116.795 232.86 117.125 ;
      VIA 232.07 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 116.775 232.84 117.145 ;
      VIA 232.07 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 111.355 232.86 111.685 ;
      VIA 232.07 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 111.335 232.84 111.705 ;
      VIA 232.07 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 105.915 232.86 106.245 ;
      VIA 232.07 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 105.895 232.84 106.265 ;
      VIA 232.07 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 100.475 232.86 100.805 ;
      VIA 232.07 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 100.455 232.84 100.825 ;
      VIA 232.07 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 95.035 232.86 95.365 ;
      VIA 232.07 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 95.015 232.84 95.385 ;
      VIA 232.07 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 89.595 232.86 89.925 ;
      VIA 232.07 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 89.575 232.84 89.945 ;
      VIA 232.07 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 84.155 232.86 84.485 ;
      VIA 232.07 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 84.135 232.84 84.505 ;
      VIA 232.07 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 78.715 232.86 79.045 ;
      VIA 232.07 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 78.695 232.84 79.065 ;
      VIA 232.07 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 73.275 232.86 73.605 ;
      VIA 232.07 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 73.255 232.84 73.625 ;
      VIA 232.07 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 67.835 232.86 68.165 ;
      VIA 232.07 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 67.815 232.84 68.185 ;
      VIA 232.07 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 62.395 232.86 62.725 ;
      VIA 232.07 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 62.375 232.84 62.745 ;
      VIA 232.07 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 56.955 232.86 57.285 ;
      VIA 232.07 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 56.935 232.84 57.305 ;
      VIA 232.07 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 51.515 232.86 51.845 ;
      VIA 232.07 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 51.495 232.84 51.865 ;
      VIA 232.07 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 46.075 232.86 46.405 ;
      VIA 232.07 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 46.055 232.84 46.425 ;
      VIA 232.07 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 40.635 232.86 40.965 ;
      VIA 232.07 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 40.615 232.84 40.985 ;
      VIA 232.07 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 35.195 232.86 35.525 ;
      VIA 232.07 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 35.175 232.84 35.545 ;
      VIA 232.07 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 29.755 232.86 30.085 ;
      VIA 232.07 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 29.735 232.84 30.105 ;
      VIA 232.07 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 24.315 232.86 24.645 ;
      VIA 232.07 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 24.295 232.84 24.665 ;
      VIA 232.07 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 18.875 232.86 19.205 ;
      VIA 232.07 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 18.855 232.84 19.225 ;
      VIA 232.07 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 13.435 232.86 13.765 ;
      VIA 232.07 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 13.415 232.84 13.785 ;
      VIA 232.07 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 7.995 232.86 8.325 ;
      VIA 232.07 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 7.975 232.84 8.345 ;
      VIA 232.07 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.28 2.555 232.86 2.885 ;
      VIA 232.07 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.3 2.535 232.84 2.905 ;
      VIA 232.07 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 232.07 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 290.875 205.72 291.205 ;
      VIA 204.93 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 290.855 205.7 291.225 ;
      VIA 204.93 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 285.435 205.72 285.765 ;
      VIA 204.93 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 285.415 205.7 285.785 ;
      VIA 204.93 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 279.995 205.72 280.325 ;
      VIA 204.93 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 279.975 205.7 280.345 ;
      VIA 204.93 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 274.555 205.72 274.885 ;
      VIA 204.93 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 274.535 205.7 274.905 ;
      VIA 204.93 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 269.115 205.72 269.445 ;
      VIA 204.93 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 269.095 205.7 269.465 ;
      VIA 204.93 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 263.675 205.72 264.005 ;
      VIA 204.93 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 263.655 205.7 264.025 ;
      VIA 204.93 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 258.235 205.72 258.565 ;
      VIA 204.93 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 258.215 205.7 258.585 ;
      VIA 204.93 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 252.795 205.72 253.125 ;
      VIA 204.93 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 252.775 205.7 253.145 ;
      VIA 204.93 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 247.355 205.72 247.685 ;
      VIA 204.93 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 247.335 205.7 247.705 ;
      VIA 204.93 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 241.915 205.72 242.245 ;
      VIA 204.93 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 241.895 205.7 242.265 ;
      VIA 204.93 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 236.475 205.72 236.805 ;
      VIA 204.93 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 236.455 205.7 236.825 ;
      VIA 204.93 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 231.035 205.72 231.365 ;
      VIA 204.93 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 231.015 205.7 231.385 ;
      VIA 204.93 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 225.595 205.72 225.925 ;
      VIA 204.93 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 225.575 205.7 225.945 ;
      VIA 204.93 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 220.155 205.72 220.485 ;
      VIA 204.93 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 220.135 205.7 220.505 ;
      VIA 204.93 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 214.715 205.72 215.045 ;
      VIA 204.93 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 214.695 205.7 215.065 ;
      VIA 204.93 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 209.275 205.72 209.605 ;
      VIA 204.93 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 209.255 205.7 209.625 ;
      VIA 204.93 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 203.835 205.72 204.165 ;
      VIA 204.93 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 203.815 205.7 204.185 ;
      VIA 204.93 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 198.395 205.72 198.725 ;
      VIA 204.93 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 198.375 205.7 198.745 ;
      VIA 204.93 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 192.955 205.72 193.285 ;
      VIA 204.93 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 192.935 205.7 193.305 ;
      VIA 204.93 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 187.515 205.72 187.845 ;
      VIA 204.93 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 187.495 205.7 187.865 ;
      VIA 204.93 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 182.075 205.72 182.405 ;
      VIA 204.93 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 182.055 205.7 182.425 ;
      VIA 204.93 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 176.635 205.72 176.965 ;
      VIA 204.93 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 176.615 205.7 176.985 ;
      VIA 204.93 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 171.195 205.72 171.525 ;
      VIA 204.93 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 171.175 205.7 171.545 ;
      VIA 204.93 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 165.755 205.72 166.085 ;
      VIA 204.93 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 165.735 205.7 166.105 ;
      VIA 204.93 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 160.315 205.72 160.645 ;
      VIA 204.93 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 160.295 205.7 160.665 ;
      VIA 204.93 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 154.875 205.72 155.205 ;
      VIA 204.93 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 154.855 205.7 155.225 ;
      VIA 204.93 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 149.435 205.72 149.765 ;
      VIA 204.93 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 149.415 205.7 149.785 ;
      VIA 204.93 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 143.995 205.72 144.325 ;
      VIA 204.93 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 143.975 205.7 144.345 ;
      VIA 204.93 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 138.555 205.72 138.885 ;
      VIA 204.93 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 138.535 205.7 138.905 ;
      VIA 204.93 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 133.115 205.72 133.445 ;
      VIA 204.93 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 133.095 205.7 133.465 ;
      VIA 204.93 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 127.675 205.72 128.005 ;
      VIA 204.93 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 127.655 205.7 128.025 ;
      VIA 204.93 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 122.235 205.72 122.565 ;
      VIA 204.93 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 122.215 205.7 122.585 ;
      VIA 204.93 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 116.795 205.72 117.125 ;
      VIA 204.93 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 116.775 205.7 117.145 ;
      VIA 204.93 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 111.355 205.72 111.685 ;
      VIA 204.93 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 111.335 205.7 111.705 ;
      VIA 204.93 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 105.915 205.72 106.245 ;
      VIA 204.93 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 105.895 205.7 106.265 ;
      VIA 204.93 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 100.475 205.72 100.805 ;
      VIA 204.93 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 100.455 205.7 100.825 ;
      VIA 204.93 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 95.035 205.72 95.365 ;
      VIA 204.93 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 95.015 205.7 95.385 ;
      VIA 204.93 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 89.595 205.72 89.925 ;
      VIA 204.93 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 89.575 205.7 89.945 ;
      VIA 204.93 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 84.155 205.72 84.485 ;
      VIA 204.93 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 84.135 205.7 84.505 ;
      VIA 204.93 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 78.715 205.72 79.045 ;
      VIA 204.93 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 78.695 205.7 79.065 ;
      VIA 204.93 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 73.275 205.72 73.605 ;
      VIA 204.93 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 73.255 205.7 73.625 ;
      VIA 204.93 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 67.835 205.72 68.165 ;
      VIA 204.93 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 67.815 205.7 68.185 ;
      VIA 204.93 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 62.395 205.72 62.725 ;
      VIA 204.93 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 62.375 205.7 62.745 ;
      VIA 204.93 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 56.955 205.72 57.285 ;
      VIA 204.93 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 56.935 205.7 57.305 ;
      VIA 204.93 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 51.515 205.72 51.845 ;
      VIA 204.93 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 51.495 205.7 51.865 ;
      VIA 204.93 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 46.075 205.72 46.405 ;
      VIA 204.93 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 46.055 205.7 46.425 ;
      VIA 204.93 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 40.635 205.72 40.965 ;
      VIA 204.93 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 40.615 205.7 40.985 ;
      VIA 204.93 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 35.195 205.72 35.525 ;
      VIA 204.93 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 35.175 205.7 35.545 ;
      VIA 204.93 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 29.755 205.72 30.085 ;
      VIA 204.93 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 29.735 205.7 30.105 ;
      VIA 204.93 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 24.315 205.72 24.645 ;
      VIA 204.93 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 24.295 205.7 24.665 ;
      VIA 204.93 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 18.875 205.72 19.205 ;
      VIA 204.93 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 18.855 205.7 19.225 ;
      VIA 204.93 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 13.435 205.72 13.765 ;
      VIA 204.93 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 13.415 205.7 13.785 ;
      VIA 204.93 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 7.995 205.72 8.325 ;
      VIA 204.93 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 7.975 205.7 8.345 ;
      VIA 204.93 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.14 2.555 205.72 2.885 ;
      VIA 204.93 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.16 2.535 205.7 2.905 ;
      VIA 204.93 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 204.93 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 290.875 178.58 291.205 ;
      VIA 177.79 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 290.855 178.56 291.225 ;
      VIA 177.79 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 285.435 178.58 285.765 ;
      VIA 177.79 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 285.415 178.56 285.785 ;
      VIA 177.79 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 279.995 178.58 280.325 ;
      VIA 177.79 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 279.975 178.56 280.345 ;
      VIA 177.79 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 274.555 178.58 274.885 ;
      VIA 177.79 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 274.535 178.56 274.905 ;
      VIA 177.79 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 269.115 178.58 269.445 ;
      VIA 177.79 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 269.095 178.56 269.465 ;
      VIA 177.79 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 263.675 178.58 264.005 ;
      VIA 177.79 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 263.655 178.56 264.025 ;
      VIA 177.79 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 258.235 178.58 258.565 ;
      VIA 177.79 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 258.215 178.56 258.585 ;
      VIA 177.79 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 252.795 178.58 253.125 ;
      VIA 177.79 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 252.775 178.56 253.145 ;
      VIA 177.79 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 247.355 178.58 247.685 ;
      VIA 177.79 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 247.335 178.56 247.705 ;
      VIA 177.79 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 241.915 178.58 242.245 ;
      VIA 177.79 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 241.895 178.56 242.265 ;
      VIA 177.79 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 236.475 178.58 236.805 ;
      VIA 177.79 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 236.455 178.56 236.825 ;
      VIA 177.79 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 231.035 178.58 231.365 ;
      VIA 177.79 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 231.015 178.56 231.385 ;
      VIA 177.79 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 225.595 178.58 225.925 ;
      VIA 177.79 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 225.575 178.56 225.945 ;
      VIA 177.79 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 220.155 178.58 220.485 ;
      VIA 177.79 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 220.135 178.56 220.505 ;
      VIA 177.79 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 214.715 178.58 215.045 ;
      VIA 177.79 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 214.695 178.56 215.065 ;
      VIA 177.79 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 209.275 178.58 209.605 ;
      VIA 177.79 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 209.255 178.56 209.625 ;
      VIA 177.79 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 203.835 178.58 204.165 ;
      VIA 177.79 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 203.815 178.56 204.185 ;
      VIA 177.79 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 198.395 178.58 198.725 ;
      VIA 177.79 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 198.375 178.56 198.745 ;
      VIA 177.79 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 192.955 178.58 193.285 ;
      VIA 177.79 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 192.935 178.56 193.305 ;
      VIA 177.79 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 187.515 178.58 187.845 ;
      VIA 177.79 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 187.495 178.56 187.865 ;
      VIA 177.79 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 182.075 178.58 182.405 ;
      VIA 177.79 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 182.055 178.56 182.425 ;
      VIA 177.79 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 176.635 178.58 176.965 ;
      VIA 177.79 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 176.615 178.56 176.985 ;
      VIA 177.79 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 171.195 178.58 171.525 ;
      VIA 177.79 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 171.175 178.56 171.545 ;
      VIA 177.79 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 165.755 178.58 166.085 ;
      VIA 177.79 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 165.735 178.56 166.105 ;
      VIA 177.79 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 160.315 178.58 160.645 ;
      VIA 177.79 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 160.295 178.56 160.665 ;
      VIA 177.79 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 154.875 178.58 155.205 ;
      VIA 177.79 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 154.855 178.56 155.225 ;
      VIA 177.79 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 149.435 178.58 149.765 ;
      VIA 177.79 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 149.415 178.56 149.785 ;
      VIA 177.79 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 143.995 178.58 144.325 ;
      VIA 177.79 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 143.975 178.56 144.345 ;
      VIA 177.79 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 138.555 178.58 138.885 ;
      VIA 177.79 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 138.535 178.56 138.905 ;
      VIA 177.79 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 133.115 178.58 133.445 ;
      VIA 177.79 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 133.095 178.56 133.465 ;
      VIA 177.79 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 127.675 178.58 128.005 ;
      VIA 177.79 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 127.655 178.56 128.025 ;
      VIA 177.79 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 122.235 178.58 122.565 ;
      VIA 177.79 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 122.215 178.56 122.585 ;
      VIA 177.79 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 116.795 178.58 117.125 ;
      VIA 177.79 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 116.775 178.56 117.145 ;
      VIA 177.79 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 111.355 178.58 111.685 ;
      VIA 177.79 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 111.335 178.56 111.705 ;
      VIA 177.79 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 105.915 178.58 106.245 ;
      VIA 177.79 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 105.895 178.56 106.265 ;
      VIA 177.79 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 100.475 178.58 100.805 ;
      VIA 177.79 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 100.455 178.56 100.825 ;
      VIA 177.79 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 95.035 178.58 95.365 ;
      VIA 177.79 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 95.015 178.56 95.385 ;
      VIA 177.79 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 89.595 178.58 89.925 ;
      VIA 177.79 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 89.575 178.56 89.945 ;
      VIA 177.79 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 84.155 178.58 84.485 ;
      VIA 177.79 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 84.135 178.56 84.505 ;
      VIA 177.79 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 78.715 178.58 79.045 ;
      VIA 177.79 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 78.695 178.56 79.065 ;
      VIA 177.79 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 73.275 178.58 73.605 ;
      VIA 177.79 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 73.255 178.56 73.625 ;
      VIA 177.79 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 67.835 178.58 68.165 ;
      VIA 177.79 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 67.815 178.56 68.185 ;
      VIA 177.79 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 62.395 178.58 62.725 ;
      VIA 177.79 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 62.375 178.56 62.745 ;
      VIA 177.79 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 56.955 178.58 57.285 ;
      VIA 177.79 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 56.935 178.56 57.305 ;
      VIA 177.79 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 51.515 178.58 51.845 ;
      VIA 177.79 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 51.495 178.56 51.865 ;
      VIA 177.79 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 46.075 178.58 46.405 ;
      VIA 177.79 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 46.055 178.56 46.425 ;
      VIA 177.79 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 40.635 178.58 40.965 ;
      VIA 177.79 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 40.615 178.56 40.985 ;
      VIA 177.79 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 35.195 178.58 35.525 ;
      VIA 177.79 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 35.175 178.56 35.545 ;
      VIA 177.79 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 29.755 178.58 30.085 ;
      VIA 177.79 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 29.735 178.56 30.105 ;
      VIA 177.79 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 24.315 178.58 24.645 ;
      VIA 177.79 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 24.295 178.56 24.665 ;
      VIA 177.79 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 18.875 178.58 19.205 ;
      VIA 177.79 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 18.855 178.56 19.225 ;
      VIA 177.79 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 13.435 178.58 13.765 ;
      VIA 177.79 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 13.415 178.56 13.785 ;
      VIA 177.79 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 7.995 178.58 8.325 ;
      VIA 177.79 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 7.975 178.56 8.345 ;
      VIA 177.79 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177 2.555 178.58 2.885 ;
      VIA 177.79 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.02 2.535 178.56 2.905 ;
      VIA 177.79 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 177.79 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 290.875 151.44 291.205 ;
      VIA 150.65 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 290.855 151.42 291.225 ;
      VIA 150.65 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 285.435 151.44 285.765 ;
      VIA 150.65 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 285.415 151.42 285.785 ;
      VIA 150.65 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 279.995 151.44 280.325 ;
      VIA 150.65 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 279.975 151.42 280.345 ;
      VIA 150.65 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 274.555 151.44 274.885 ;
      VIA 150.65 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 274.535 151.42 274.905 ;
      VIA 150.65 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 269.115 151.44 269.445 ;
      VIA 150.65 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 269.095 151.42 269.465 ;
      VIA 150.65 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 263.675 151.44 264.005 ;
      VIA 150.65 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 263.655 151.42 264.025 ;
      VIA 150.65 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 258.235 151.44 258.565 ;
      VIA 150.65 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 258.215 151.42 258.585 ;
      VIA 150.65 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 252.795 151.44 253.125 ;
      VIA 150.65 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 252.775 151.42 253.145 ;
      VIA 150.65 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 247.355 151.44 247.685 ;
      VIA 150.65 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 247.335 151.42 247.705 ;
      VIA 150.65 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 241.915 151.44 242.245 ;
      VIA 150.65 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 241.895 151.42 242.265 ;
      VIA 150.65 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 236.475 151.44 236.805 ;
      VIA 150.65 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 236.455 151.42 236.825 ;
      VIA 150.65 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 231.035 151.44 231.365 ;
      VIA 150.65 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 231.015 151.42 231.385 ;
      VIA 150.65 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 225.595 151.44 225.925 ;
      VIA 150.65 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 225.575 151.42 225.945 ;
      VIA 150.65 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 220.155 151.44 220.485 ;
      VIA 150.65 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 220.135 151.42 220.505 ;
      VIA 150.65 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 214.715 151.44 215.045 ;
      VIA 150.65 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 214.695 151.42 215.065 ;
      VIA 150.65 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 209.275 151.44 209.605 ;
      VIA 150.65 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 209.255 151.42 209.625 ;
      VIA 150.65 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 203.835 151.44 204.165 ;
      VIA 150.65 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 203.815 151.42 204.185 ;
      VIA 150.65 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 198.395 151.44 198.725 ;
      VIA 150.65 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 198.375 151.42 198.745 ;
      VIA 150.65 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 192.955 151.44 193.285 ;
      VIA 150.65 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 192.935 151.42 193.305 ;
      VIA 150.65 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 187.515 151.44 187.845 ;
      VIA 150.65 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 187.495 151.42 187.865 ;
      VIA 150.65 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 182.075 151.44 182.405 ;
      VIA 150.65 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 182.055 151.42 182.425 ;
      VIA 150.65 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 176.635 151.44 176.965 ;
      VIA 150.65 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 176.615 151.42 176.985 ;
      VIA 150.65 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 171.195 151.44 171.525 ;
      VIA 150.65 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 171.175 151.42 171.545 ;
      VIA 150.65 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 165.755 151.44 166.085 ;
      VIA 150.65 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 165.735 151.42 166.105 ;
      VIA 150.65 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 160.315 151.44 160.645 ;
      VIA 150.65 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 160.295 151.42 160.665 ;
      VIA 150.65 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 154.875 151.44 155.205 ;
      VIA 150.65 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 154.855 151.42 155.225 ;
      VIA 150.65 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 149.435 151.44 149.765 ;
      VIA 150.65 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 149.415 151.42 149.785 ;
      VIA 150.65 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 143.995 151.44 144.325 ;
      VIA 150.65 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 143.975 151.42 144.345 ;
      VIA 150.65 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 138.555 151.44 138.885 ;
      VIA 150.65 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 138.535 151.42 138.905 ;
      VIA 150.65 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 133.115 151.44 133.445 ;
      VIA 150.65 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 133.095 151.42 133.465 ;
      VIA 150.65 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 127.675 151.44 128.005 ;
      VIA 150.65 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 127.655 151.42 128.025 ;
      VIA 150.65 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 122.235 151.44 122.565 ;
      VIA 150.65 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 122.215 151.42 122.585 ;
      VIA 150.65 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 116.795 151.44 117.125 ;
      VIA 150.65 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 116.775 151.42 117.145 ;
      VIA 150.65 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 111.355 151.44 111.685 ;
      VIA 150.65 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 111.335 151.42 111.705 ;
      VIA 150.65 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 105.915 151.44 106.245 ;
      VIA 150.65 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 105.895 151.42 106.265 ;
      VIA 150.65 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 100.475 151.44 100.805 ;
      VIA 150.65 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 100.455 151.42 100.825 ;
      VIA 150.65 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 95.035 151.44 95.365 ;
      VIA 150.65 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 95.015 151.42 95.385 ;
      VIA 150.65 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 89.595 151.44 89.925 ;
      VIA 150.65 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 89.575 151.42 89.945 ;
      VIA 150.65 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 84.155 151.44 84.485 ;
      VIA 150.65 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 84.135 151.42 84.505 ;
      VIA 150.65 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 78.715 151.44 79.045 ;
      VIA 150.65 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 78.695 151.42 79.065 ;
      VIA 150.65 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 73.275 151.44 73.605 ;
      VIA 150.65 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 73.255 151.42 73.625 ;
      VIA 150.65 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 67.835 151.44 68.165 ;
      VIA 150.65 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 67.815 151.42 68.185 ;
      VIA 150.65 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 62.395 151.44 62.725 ;
      VIA 150.65 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 62.375 151.42 62.745 ;
      VIA 150.65 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 56.955 151.44 57.285 ;
      VIA 150.65 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 56.935 151.42 57.305 ;
      VIA 150.65 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 51.515 151.44 51.845 ;
      VIA 150.65 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 51.495 151.42 51.865 ;
      VIA 150.65 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 46.075 151.44 46.405 ;
      VIA 150.65 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 46.055 151.42 46.425 ;
      VIA 150.65 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 40.635 151.44 40.965 ;
      VIA 150.65 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 40.615 151.42 40.985 ;
      VIA 150.65 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 35.195 151.44 35.525 ;
      VIA 150.65 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 35.175 151.42 35.545 ;
      VIA 150.65 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 29.755 151.44 30.085 ;
      VIA 150.65 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 29.735 151.42 30.105 ;
      VIA 150.65 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 24.315 151.44 24.645 ;
      VIA 150.65 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 24.295 151.42 24.665 ;
      VIA 150.65 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 18.875 151.44 19.205 ;
      VIA 150.65 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 18.855 151.42 19.225 ;
      VIA 150.65 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 13.435 151.44 13.765 ;
      VIA 150.65 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 13.415 151.42 13.785 ;
      VIA 150.65 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 7.995 151.44 8.325 ;
      VIA 150.65 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 7.975 151.42 8.345 ;
      VIA 150.65 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 2.555 151.44 2.885 ;
      VIA 150.65 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 2.535 151.42 2.905 ;
      VIA 150.65 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 290.875 124.3 291.205 ;
      VIA 123.51 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 290.855 124.28 291.225 ;
      VIA 123.51 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 285.435 124.3 285.765 ;
      VIA 123.51 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 285.415 124.28 285.785 ;
      VIA 123.51 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 279.995 124.3 280.325 ;
      VIA 123.51 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 279.975 124.28 280.345 ;
      VIA 123.51 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 274.555 124.3 274.885 ;
      VIA 123.51 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 274.535 124.28 274.905 ;
      VIA 123.51 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 269.115 124.3 269.445 ;
      VIA 123.51 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 269.095 124.28 269.465 ;
      VIA 123.51 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 263.675 124.3 264.005 ;
      VIA 123.51 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 263.655 124.28 264.025 ;
      VIA 123.51 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 258.235 124.3 258.565 ;
      VIA 123.51 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 258.215 124.28 258.585 ;
      VIA 123.51 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 252.795 124.3 253.125 ;
      VIA 123.51 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 252.775 124.28 253.145 ;
      VIA 123.51 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 247.355 124.3 247.685 ;
      VIA 123.51 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 247.335 124.28 247.705 ;
      VIA 123.51 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 241.915 124.3 242.245 ;
      VIA 123.51 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 241.895 124.28 242.265 ;
      VIA 123.51 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 236.475 124.3 236.805 ;
      VIA 123.51 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 236.455 124.28 236.825 ;
      VIA 123.51 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 231.035 124.3 231.365 ;
      VIA 123.51 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 231.015 124.28 231.385 ;
      VIA 123.51 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 225.595 124.3 225.925 ;
      VIA 123.51 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 225.575 124.28 225.945 ;
      VIA 123.51 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 220.155 124.3 220.485 ;
      VIA 123.51 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 220.135 124.28 220.505 ;
      VIA 123.51 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 214.715 124.3 215.045 ;
      VIA 123.51 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 214.695 124.28 215.065 ;
      VIA 123.51 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 209.275 124.3 209.605 ;
      VIA 123.51 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 209.255 124.28 209.625 ;
      VIA 123.51 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 203.835 124.3 204.165 ;
      VIA 123.51 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 203.815 124.28 204.185 ;
      VIA 123.51 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 198.395 124.3 198.725 ;
      VIA 123.51 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 198.375 124.28 198.745 ;
      VIA 123.51 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 192.955 124.3 193.285 ;
      VIA 123.51 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 192.935 124.28 193.305 ;
      VIA 123.51 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 187.515 124.3 187.845 ;
      VIA 123.51 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 187.495 124.28 187.865 ;
      VIA 123.51 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 182.075 124.3 182.405 ;
      VIA 123.51 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 182.055 124.28 182.425 ;
      VIA 123.51 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 176.635 124.3 176.965 ;
      VIA 123.51 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 176.615 124.28 176.985 ;
      VIA 123.51 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 171.195 124.3 171.525 ;
      VIA 123.51 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 171.175 124.28 171.545 ;
      VIA 123.51 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 165.755 124.3 166.085 ;
      VIA 123.51 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 165.735 124.28 166.105 ;
      VIA 123.51 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 160.315 124.3 160.645 ;
      VIA 123.51 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 160.295 124.28 160.665 ;
      VIA 123.51 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 154.875 124.3 155.205 ;
      VIA 123.51 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 154.855 124.28 155.225 ;
      VIA 123.51 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 149.435 124.3 149.765 ;
      VIA 123.51 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 149.415 124.28 149.785 ;
      VIA 123.51 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 143.995 124.3 144.325 ;
      VIA 123.51 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 143.975 124.28 144.345 ;
      VIA 123.51 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 138.555 124.3 138.885 ;
      VIA 123.51 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 138.535 124.28 138.905 ;
      VIA 123.51 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 133.115 124.3 133.445 ;
      VIA 123.51 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 133.095 124.28 133.465 ;
      VIA 123.51 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 127.675 124.3 128.005 ;
      VIA 123.51 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 127.655 124.28 128.025 ;
      VIA 123.51 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 122.235 124.3 122.565 ;
      VIA 123.51 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 122.215 124.28 122.585 ;
      VIA 123.51 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 116.795 124.3 117.125 ;
      VIA 123.51 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 116.775 124.28 117.145 ;
      VIA 123.51 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 111.355 124.3 111.685 ;
      VIA 123.51 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 111.335 124.28 111.705 ;
      VIA 123.51 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 105.915 124.3 106.245 ;
      VIA 123.51 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 105.895 124.28 106.265 ;
      VIA 123.51 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 100.475 124.3 100.805 ;
      VIA 123.51 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 100.455 124.28 100.825 ;
      VIA 123.51 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 95.035 124.3 95.365 ;
      VIA 123.51 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 95.015 124.28 95.385 ;
      VIA 123.51 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 89.595 124.3 89.925 ;
      VIA 123.51 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 89.575 124.28 89.945 ;
      VIA 123.51 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 84.155 124.3 84.485 ;
      VIA 123.51 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 84.135 124.28 84.505 ;
      VIA 123.51 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 78.715 124.3 79.045 ;
      VIA 123.51 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 78.695 124.28 79.065 ;
      VIA 123.51 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 73.275 124.3 73.605 ;
      VIA 123.51 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 73.255 124.28 73.625 ;
      VIA 123.51 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 67.835 124.3 68.165 ;
      VIA 123.51 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 67.815 124.28 68.185 ;
      VIA 123.51 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 62.395 124.3 62.725 ;
      VIA 123.51 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 62.375 124.28 62.745 ;
      VIA 123.51 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 56.955 124.3 57.285 ;
      VIA 123.51 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 56.935 124.28 57.305 ;
      VIA 123.51 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 51.515 124.3 51.845 ;
      VIA 123.51 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 51.495 124.28 51.865 ;
      VIA 123.51 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 46.075 124.3 46.405 ;
      VIA 123.51 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 46.055 124.28 46.425 ;
      VIA 123.51 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 40.635 124.3 40.965 ;
      VIA 123.51 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 40.615 124.28 40.985 ;
      VIA 123.51 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 35.195 124.3 35.525 ;
      VIA 123.51 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 35.175 124.28 35.545 ;
      VIA 123.51 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 29.755 124.3 30.085 ;
      VIA 123.51 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 29.735 124.28 30.105 ;
      VIA 123.51 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 24.315 124.3 24.645 ;
      VIA 123.51 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 24.295 124.28 24.665 ;
      VIA 123.51 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 18.875 124.3 19.205 ;
      VIA 123.51 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 18.855 124.28 19.225 ;
      VIA 123.51 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 13.435 124.3 13.765 ;
      VIA 123.51 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 13.415 124.28 13.785 ;
      VIA 123.51 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 7.995 124.3 8.325 ;
      VIA 123.51 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 7.975 124.28 8.345 ;
      VIA 123.51 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 2.555 124.3 2.885 ;
      VIA 123.51 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 2.535 124.28 2.905 ;
      VIA 123.51 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 290.875 97.16 291.205 ;
      VIA 96.37 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 290.855 97.14 291.225 ;
      VIA 96.37 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 285.435 97.16 285.765 ;
      VIA 96.37 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 285.415 97.14 285.785 ;
      VIA 96.37 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 279.995 97.16 280.325 ;
      VIA 96.37 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 279.975 97.14 280.345 ;
      VIA 96.37 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 274.555 97.16 274.885 ;
      VIA 96.37 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 274.535 97.14 274.905 ;
      VIA 96.37 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 269.115 97.16 269.445 ;
      VIA 96.37 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 269.095 97.14 269.465 ;
      VIA 96.37 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 263.675 97.16 264.005 ;
      VIA 96.37 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 263.655 97.14 264.025 ;
      VIA 96.37 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 258.235 97.16 258.565 ;
      VIA 96.37 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 258.215 97.14 258.585 ;
      VIA 96.37 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 252.795 97.16 253.125 ;
      VIA 96.37 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 252.775 97.14 253.145 ;
      VIA 96.37 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 247.355 97.16 247.685 ;
      VIA 96.37 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 247.335 97.14 247.705 ;
      VIA 96.37 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 241.915 97.16 242.245 ;
      VIA 96.37 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 241.895 97.14 242.265 ;
      VIA 96.37 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 236.475 97.16 236.805 ;
      VIA 96.37 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 236.455 97.14 236.825 ;
      VIA 96.37 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 231.035 97.16 231.365 ;
      VIA 96.37 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 231.015 97.14 231.385 ;
      VIA 96.37 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 225.595 97.16 225.925 ;
      VIA 96.37 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 225.575 97.14 225.945 ;
      VIA 96.37 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 220.155 97.16 220.485 ;
      VIA 96.37 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 220.135 97.14 220.505 ;
      VIA 96.37 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 214.715 97.16 215.045 ;
      VIA 96.37 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 214.695 97.14 215.065 ;
      VIA 96.37 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 209.275 97.16 209.605 ;
      VIA 96.37 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 209.255 97.14 209.625 ;
      VIA 96.37 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 203.835 97.16 204.165 ;
      VIA 96.37 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 203.815 97.14 204.185 ;
      VIA 96.37 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 198.395 97.16 198.725 ;
      VIA 96.37 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 198.375 97.14 198.745 ;
      VIA 96.37 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 192.955 97.16 193.285 ;
      VIA 96.37 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 192.935 97.14 193.305 ;
      VIA 96.37 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 187.515 97.16 187.845 ;
      VIA 96.37 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 187.495 97.14 187.865 ;
      VIA 96.37 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 182.075 97.16 182.405 ;
      VIA 96.37 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 182.055 97.14 182.425 ;
      VIA 96.37 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 176.635 97.16 176.965 ;
      VIA 96.37 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 176.615 97.14 176.985 ;
      VIA 96.37 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 171.195 97.16 171.525 ;
      VIA 96.37 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 171.175 97.14 171.545 ;
      VIA 96.37 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 165.755 97.16 166.085 ;
      VIA 96.37 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 165.735 97.14 166.105 ;
      VIA 96.37 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 160.315 97.16 160.645 ;
      VIA 96.37 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 160.295 97.14 160.665 ;
      VIA 96.37 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 154.875 97.16 155.205 ;
      VIA 96.37 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 154.855 97.14 155.225 ;
      VIA 96.37 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 149.435 97.16 149.765 ;
      VIA 96.37 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 149.415 97.14 149.785 ;
      VIA 96.37 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 143.995 97.16 144.325 ;
      VIA 96.37 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 143.975 97.14 144.345 ;
      VIA 96.37 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 138.555 97.16 138.885 ;
      VIA 96.37 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 138.535 97.14 138.905 ;
      VIA 96.37 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 133.115 97.16 133.445 ;
      VIA 96.37 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 133.095 97.14 133.465 ;
      VIA 96.37 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 127.675 97.16 128.005 ;
      VIA 96.37 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 127.655 97.14 128.025 ;
      VIA 96.37 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 122.235 97.16 122.565 ;
      VIA 96.37 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 122.215 97.14 122.585 ;
      VIA 96.37 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 116.795 97.16 117.125 ;
      VIA 96.37 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 116.775 97.14 117.145 ;
      VIA 96.37 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 111.355 97.16 111.685 ;
      VIA 96.37 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 111.335 97.14 111.705 ;
      VIA 96.37 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 105.915 97.16 106.245 ;
      VIA 96.37 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 105.895 97.14 106.265 ;
      VIA 96.37 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 100.475 97.16 100.805 ;
      VIA 96.37 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 100.455 97.14 100.825 ;
      VIA 96.37 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 95.035 97.16 95.365 ;
      VIA 96.37 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 95.015 97.14 95.385 ;
      VIA 96.37 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 89.595 97.16 89.925 ;
      VIA 96.37 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 89.575 97.14 89.945 ;
      VIA 96.37 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 84.155 97.16 84.485 ;
      VIA 96.37 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 84.135 97.14 84.505 ;
      VIA 96.37 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 78.715 97.16 79.045 ;
      VIA 96.37 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 78.695 97.14 79.065 ;
      VIA 96.37 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 73.275 97.16 73.605 ;
      VIA 96.37 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 73.255 97.14 73.625 ;
      VIA 96.37 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 67.835 97.16 68.165 ;
      VIA 96.37 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 67.815 97.14 68.185 ;
      VIA 96.37 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 62.395 97.16 62.725 ;
      VIA 96.37 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 62.375 97.14 62.745 ;
      VIA 96.37 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 56.955 97.16 57.285 ;
      VIA 96.37 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 56.935 97.14 57.305 ;
      VIA 96.37 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 51.515 97.16 51.845 ;
      VIA 96.37 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 51.495 97.14 51.865 ;
      VIA 96.37 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 46.075 97.16 46.405 ;
      VIA 96.37 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 46.055 97.14 46.425 ;
      VIA 96.37 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 40.635 97.16 40.965 ;
      VIA 96.37 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 40.615 97.14 40.985 ;
      VIA 96.37 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 35.195 97.16 35.525 ;
      VIA 96.37 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 35.175 97.14 35.545 ;
      VIA 96.37 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 29.755 97.16 30.085 ;
      VIA 96.37 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 29.735 97.14 30.105 ;
      VIA 96.37 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 24.315 97.16 24.645 ;
      VIA 96.37 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 24.295 97.14 24.665 ;
      VIA 96.37 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 18.875 97.16 19.205 ;
      VIA 96.37 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 18.855 97.14 19.225 ;
      VIA 96.37 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 13.435 97.16 13.765 ;
      VIA 96.37 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 13.415 97.14 13.785 ;
      VIA 96.37 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 7.995 97.16 8.325 ;
      VIA 96.37 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 7.975 97.14 8.345 ;
      VIA 96.37 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 2.555 97.16 2.885 ;
      VIA 96.37 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 2.535 97.14 2.905 ;
      VIA 96.37 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 290.875 70.02 291.205 ;
      VIA 69.23 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 290.855 70 291.225 ;
      VIA 69.23 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 285.435 70.02 285.765 ;
      VIA 69.23 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 285.415 70 285.785 ;
      VIA 69.23 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 279.995 70.02 280.325 ;
      VIA 69.23 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 279.975 70 280.345 ;
      VIA 69.23 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 274.555 70.02 274.885 ;
      VIA 69.23 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 274.535 70 274.905 ;
      VIA 69.23 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 269.115 70.02 269.445 ;
      VIA 69.23 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 269.095 70 269.465 ;
      VIA 69.23 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 263.675 70.02 264.005 ;
      VIA 69.23 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 263.655 70 264.025 ;
      VIA 69.23 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 258.235 70.02 258.565 ;
      VIA 69.23 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 258.215 70 258.585 ;
      VIA 69.23 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 252.795 70.02 253.125 ;
      VIA 69.23 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 252.775 70 253.145 ;
      VIA 69.23 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 247.355 70.02 247.685 ;
      VIA 69.23 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 247.335 70 247.705 ;
      VIA 69.23 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 241.915 70.02 242.245 ;
      VIA 69.23 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 241.895 70 242.265 ;
      VIA 69.23 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 236.475 70.02 236.805 ;
      VIA 69.23 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 236.455 70 236.825 ;
      VIA 69.23 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 231.035 70.02 231.365 ;
      VIA 69.23 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 231.015 70 231.385 ;
      VIA 69.23 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 225.595 70.02 225.925 ;
      VIA 69.23 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 225.575 70 225.945 ;
      VIA 69.23 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 220.155 70.02 220.485 ;
      VIA 69.23 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 220.135 70 220.505 ;
      VIA 69.23 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 214.715 70.02 215.045 ;
      VIA 69.23 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 214.695 70 215.065 ;
      VIA 69.23 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 209.275 70.02 209.605 ;
      VIA 69.23 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 209.255 70 209.625 ;
      VIA 69.23 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 203.835 70.02 204.165 ;
      VIA 69.23 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 203.815 70 204.185 ;
      VIA 69.23 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 198.395 70.02 198.725 ;
      VIA 69.23 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 198.375 70 198.745 ;
      VIA 69.23 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 192.955 70.02 193.285 ;
      VIA 69.23 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 192.935 70 193.305 ;
      VIA 69.23 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 187.515 70.02 187.845 ;
      VIA 69.23 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 187.495 70 187.865 ;
      VIA 69.23 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 182.075 70.02 182.405 ;
      VIA 69.23 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 182.055 70 182.425 ;
      VIA 69.23 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 176.635 70.02 176.965 ;
      VIA 69.23 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 176.615 70 176.985 ;
      VIA 69.23 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 171.195 70.02 171.525 ;
      VIA 69.23 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 171.175 70 171.545 ;
      VIA 69.23 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 165.755 70.02 166.085 ;
      VIA 69.23 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 165.735 70 166.105 ;
      VIA 69.23 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 160.315 70.02 160.645 ;
      VIA 69.23 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 160.295 70 160.665 ;
      VIA 69.23 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 154.875 70.02 155.205 ;
      VIA 69.23 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 154.855 70 155.225 ;
      VIA 69.23 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 149.435 70.02 149.765 ;
      VIA 69.23 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 149.415 70 149.785 ;
      VIA 69.23 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 143.995 70.02 144.325 ;
      VIA 69.23 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 143.975 70 144.345 ;
      VIA 69.23 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 138.555 70.02 138.885 ;
      VIA 69.23 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 138.535 70 138.905 ;
      VIA 69.23 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 133.115 70.02 133.445 ;
      VIA 69.23 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 133.095 70 133.465 ;
      VIA 69.23 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 127.675 70.02 128.005 ;
      VIA 69.23 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 127.655 70 128.025 ;
      VIA 69.23 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 122.235 70.02 122.565 ;
      VIA 69.23 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 122.215 70 122.585 ;
      VIA 69.23 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 116.795 70.02 117.125 ;
      VIA 69.23 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 116.775 70 117.145 ;
      VIA 69.23 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 111.355 70.02 111.685 ;
      VIA 69.23 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 111.335 70 111.705 ;
      VIA 69.23 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 105.915 70.02 106.245 ;
      VIA 69.23 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 105.895 70 106.265 ;
      VIA 69.23 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 100.475 70.02 100.805 ;
      VIA 69.23 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 100.455 70 100.825 ;
      VIA 69.23 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 95.035 70.02 95.365 ;
      VIA 69.23 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 95.015 70 95.385 ;
      VIA 69.23 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 89.595 70.02 89.925 ;
      VIA 69.23 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 89.575 70 89.945 ;
      VIA 69.23 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 84.155 70.02 84.485 ;
      VIA 69.23 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 84.135 70 84.505 ;
      VIA 69.23 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 78.715 70.02 79.045 ;
      VIA 69.23 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 78.695 70 79.065 ;
      VIA 69.23 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 73.275 70.02 73.605 ;
      VIA 69.23 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 73.255 70 73.625 ;
      VIA 69.23 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 67.835 70.02 68.165 ;
      VIA 69.23 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 67.815 70 68.185 ;
      VIA 69.23 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 62.395 70.02 62.725 ;
      VIA 69.23 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 62.375 70 62.745 ;
      VIA 69.23 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 56.955 70.02 57.285 ;
      VIA 69.23 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 56.935 70 57.305 ;
      VIA 69.23 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 51.515 70.02 51.845 ;
      VIA 69.23 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 51.495 70 51.865 ;
      VIA 69.23 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 46.075 70.02 46.405 ;
      VIA 69.23 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 46.055 70 46.425 ;
      VIA 69.23 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 40.635 70.02 40.965 ;
      VIA 69.23 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 40.615 70 40.985 ;
      VIA 69.23 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 35.195 70.02 35.525 ;
      VIA 69.23 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 35.175 70 35.545 ;
      VIA 69.23 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 29.755 70.02 30.085 ;
      VIA 69.23 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 29.735 70 30.105 ;
      VIA 69.23 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 24.315 70.02 24.645 ;
      VIA 69.23 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 24.295 70 24.665 ;
      VIA 69.23 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 18.875 70.02 19.205 ;
      VIA 69.23 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 18.855 70 19.225 ;
      VIA 69.23 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 13.435 70.02 13.765 ;
      VIA 69.23 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 13.415 70 13.785 ;
      VIA 69.23 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 7.995 70.02 8.325 ;
      VIA 69.23 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 7.975 70 8.345 ;
      VIA 69.23 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 2.555 70.02 2.885 ;
      VIA 69.23 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 2.535 70 2.905 ;
      VIA 69.23 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 290.875 42.88 291.205 ;
      VIA 42.09 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 290.855 42.86 291.225 ;
      VIA 42.09 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 285.435 42.88 285.765 ;
      VIA 42.09 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 285.415 42.86 285.785 ;
      VIA 42.09 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 279.995 42.88 280.325 ;
      VIA 42.09 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 279.975 42.86 280.345 ;
      VIA 42.09 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 274.555 42.88 274.885 ;
      VIA 42.09 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 274.535 42.86 274.905 ;
      VIA 42.09 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 269.115 42.88 269.445 ;
      VIA 42.09 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 269.095 42.86 269.465 ;
      VIA 42.09 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 263.675 42.88 264.005 ;
      VIA 42.09 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 263.655 42.86 264.025 ;
      VIA 42.09 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 258.235 42.88 258.565 ;
      VIA 42.09 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 258.215 42.86 258.585 ;
      VIA 42.09 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 252.795 42.88 253.125 ;
      VIA 42.09 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 252.775 42.86 253.145 ;
      VIA 42.09 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 247.355 42.88 247.685 ;
      VIA 42.09 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 247.335 42.86 247.705 ;
      VIA 42.09 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 241.915 42.88 242.245 ;
      VIA 42.09 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 241.895 42.86 242.265 ;
      VIA 42.09 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 236.475 42.88 236.805 ;
      VIA 42.09 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 236.455 42.86 236.825 ;
      VIA 42.09 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 231.035 42.88 231.365 ;
      VIA 42.09 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 231.015 42.86 231.385 ;
      VIA 42.09 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 225.595 42.88 225.925 ;
      VIA 42.09 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 225.575 42.86 225.945 ;
      VIA 42.09 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 220.155 42.88 220.485 ;
      VIA 42.09 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 220.135 42.86 220.505 ;
      VIA 42.09 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 214.715 42.88 215.045 ;
      VIA 42.09 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 214.695 42.86 215.065 ;
      VIA 42.09 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 209.275 42.88 209.605 ;
      VIA 42.09 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 209.255 42.86 209.625 ;
      VIA 42.09 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 203.835 42.88 204.165 ;
      VIA 42.09 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 203.815 42.86 204.185 ;
      VIA 42.09 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 198.395 42.88 198.725 ;
      VIA 42.09 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 198.375 42.86 198.745 ;
      VIA 42.09 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 192.955 42.88 193.285 ;
      VIA 42.09 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 192.935 42.86 193.305 ;
      VIA 42.09 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 187.515 42.88 187.845 ;
      VIA 42.09 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 187.495 42.86 187.865 ;
      VIA 42.09 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 182.075 42.88 182.405 ;
      VIA 42.09 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 182.055 42.86 182.425 ;
      VIA 42.09 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 176.635 42.88 176.965 ;
      VIA 42.09 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 176.615 42.86 176.985 ;
      VIA 42.09 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 171.195 42.88 171.525 ;
      VIA 42.09 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 171.175 42.86 171.545 ;
      VIA 42.09 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 165.755 42.88 166.085 ;
      VIA 42.09 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 165.735 42.86 166.105 ;
      VIA 42.09 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 160.315 42.88 160.645 ;
      VIA 42.09 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 160.295 42.86 160.665 ;
      VIA 42.09 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 154.875 42.88 155.205 ;
      VIA 42.09 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 154.855 42.86 155.225 ;
      VIA 42.09 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 149.435 42.88 149.765 ;
      VIA 42.09 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 149.415 42.86 149.785 ;
      VIA 42.09 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 143.995 42.88 144.325 ;
      VIA 42.09 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 143.975 42.86 144.345 ;
      VIA 42.09 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 138.555 42.88 138.885 ;
      VIA 42.09 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 138.535 42.86 138.905 ;
      VIA 42.09 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 133.115 42.88 133.445 ;
      VIA 42.09 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 133.095 42.86 133.465 ;
      VIA 42.09 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 127.675 42.88 128.005 ;
      VIA 42.09 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 127.655 42.86 128.025 ;
      VIA 42.09 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 122.235 42.88 122.565 ;
      VIA 42.09 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 122.215 42.86 122.585 ;
      VIA 42.09 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 116.795 42.88 117.125 ;
      VIA 42.09 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 116.775 42.86 117.145 ;
      VIA 42.09 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 111.355 42.88 111.685 ;
      VIA 42.09 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 111.335 42.86 111.705 ;
      VIA 42.09 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 105.915 42.88 106.245 ;
      VIA 42.09 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 105.895 42.86 106.265 ;
      VIA 42.09 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 100.475 42.88 100.805 ;
      VIA 42.09 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 100.455 42.86 100.825 ;
      VIA 42.09 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 95.035 42.88 95.365 ;
      VIA 42.09 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 95.015 42.86 95.385 ;
      VIA 42.09 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 89.595 42.88 89.925 ;
      VIA 42.09 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 89.575 42.86 89.945 ;
      VIA 42.09 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 84.155 42.88 84.485 ;
      VIA 42.09 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 84.135 42.86 84.505 ;
      VIA 42.09 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 78.715 42.88 79.045 ;
      VIA 42.09 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 78.695 42.86 79.065 ;
      VIA 42.09 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 73.275 42.88 73.605 ;
      VIA 42.09 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 73.255 42.86 73.625 ;
      VIA 42.09 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 67.835 42.88 68.165 ;
      VIA 42.09 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 67.815 42.86 68.185 ;
      VIA 42.09 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 62.395 42.88 62.725 ;
      VIA 42.09 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 62.375 42.86 62.745 ;
      VIA 42.09 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 56.955 42.88 57.285 ;
      VIA 42.09 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 56.935 42.86 57.305 ;
      VIA 42.09 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 51.515 42.88 51.845 ;
      VIA 42.09 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 51.495 42.86 51.865 ;
      VIA 42.09 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 46.075 42.88 46.405 ;
      VIA 42.09 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 46.055 42.86 46.425 ;
      VIA 42.09 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 40.635 42.88 40.965 ;
      VIA 42.09 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 40.615 42.86 40.985 ;
      VIA 42.09 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 35.195 42.88 35.525 ;
      VIA 42.09 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 35.175 42.86 35.545 ;
      VIA 42.09 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 29.755 42.88 30.085 ;
      VIA 42.09 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 29.735 42.86 30.105 ;
      VIA 42.09 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 24.315 42.88 24.645 ;
      VIA 42.09 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 24.295 42.86 24.665 ;
      VIA 42.09 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 18.875 42.88 19.205 ;
      VIA 42.09 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 18.855 42.86 19.225 ;
      VIA 42.09 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 13.435 42.88 13.765 ;
      VIA 42.09 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 13.415 42.86 13.785 ;
      VIA 42.09 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 7.995 42.88 8.325 ;
      VIA 42.09 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 7.975 42.86 8.345 ;
      VIA 42.09 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 2.555 42.88 2.885 ;
      VIA 42.09 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 2.535 42.86 2.905 ;
      VIA 42.09 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 290.875 15.74 291.205 ;
      VIA 14.95 291.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 290.855 15.72 291.225 ;
      VIA 14.95 291.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 291.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 285.435 15.74 285.765 ;
      VIA 14.95 285.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 285.415 15.72 285.785 ;
      VIA 14.95 285.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 285.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 279.995 15.74 280.325 ;
      VIA 14.95 280.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 279.975 15.72 280.345 ;
      VIA 14.95 280.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 280.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 274.555 15.74 274.885 ;
      VIA 14.95 274.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 274.535 15.72 274.905 ;
      VIA 14.95 274.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 274.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 269.115 15.74 269.445 ;
      VIA 14.95 269.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 269.095 15.72 269.465 ;
      VIA 14.95 269.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 269.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 263.675 15.74 264.005 ;
      VIA 14.95 263.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 263.655 15.72 264.025 ;
      VIA 14.95 263.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 263.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 258.235 15.74 258.565 ;
      VIA 14.95 258.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 258.215 15.72 258.585 ;
      VIA 14.95 258.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 258.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 252.795 15.74 253.125 ;
      VIA 14.95 252.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 252.775 15.72 253.145 ;
      VIA 14.95 252.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 252.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 247.355 15.74 247.685 ;
      VIA 14.95 247.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 247.335 15.72 247.705 ;
      VIA 14.95 247.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 247.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 241.915 15.74 242.245 ;
      VIA 14.95 242.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 241.895 15.72 242.265 ;
      VIA 14.95 242.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 242.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 236.475 15.74 236.805 ;
      VIA 14.95 236.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 236.455 15.72 236.825 ;
      VIA 14.95 236.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 236.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 231.035 15.74 231.365 ;
      VIA 14.95 231.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 231.015 15.72 231.385 ;
      VIA 14.95 231.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 231.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 225.595 15.74 225.925 ;
      VIA 14.95 225.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 225.575 15.72 225.945 ;
      VIA 14.95 225.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 225.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 220.155 15.74 220.485 ;
      VIA 14.95 220.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 220.135 15.72 220.505 ;
      VIA 14.95 220.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 220.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 214.715 15.74 215.045 ;
      VIA 14.95 214.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 214.695 15.72 215.065 ;
      VIA 14.95 214.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 214.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 209.275 15.74 209.605 ;
      VIA 14.95 209.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 209.255 15.72 209.625 ;
      VIA 14.95 209.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 209.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 203.835 15.74 204.165 ;
      VIA 14.95 204 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 203.815 15.72 204.185 ;
      VIA 14.95 204 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 204 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 198.395 15.74 198.725 ;
      VIA 14.95 198.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 198.375 15.72 198.745 ;
      VIA 14.95 198.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 198.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 192.955 15.74 193.285 ;
      VIA 14.95 193.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 192.935 15.72 193.305 ;
      VIA 14.95 193.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 193.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 187.515 15.74 187.845 ;
      VIA 14.95 187.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 187.495 15.72 187.865 ;
      VIA 14.95 187.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 187.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 182.075 15.74 182.405 ;
      VIA 14.95 182.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 182.055 15.72 182.425 ;
      VIA 14.95 182.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 182.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 176.635 15.74 176.965 ;
      VIA 14.95 176.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 176.615 15.72 176.985 ;
      VIA 14.95 176.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 176.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 171.195 15.74 171.525 ;
      VIA 14.95 171.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 171.175 15.72 171.545 ;
      VIA 14.95 171.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 171.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 165.755 15.74 166.085 ;
      VIA 14.95 165.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 165.735 15.72 166.105 ;
      VIA 14.95 165.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 165.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 160.315 15.74 160.645 ;
      VIA 14.95 160.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 160.295 15.72 160.665 ;
      VIA 14.95 160.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 160.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 154.875 15.74 155.205 ;
      VIA 14.95 155.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 154.855 15.72 155.225 ;
      VIA 14.95 155.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 155.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 149.435 15.74 149.765 ;
      VIA 14.95 149.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 149.415 15.72 149.785 ;
      VIA 14.95 149.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 149.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 143.995 15.74 144.325 ;
      VIA 14.95 144.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 143.975 15.72 144.345 ;
      VIA 14.95 144.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 144.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 138.555 15.74 138.885 ;
      VIA 14.95 138.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 138.535 15.72 138.905 ;
      VIA 14.95 138.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 138.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 133.115 15.74 133.445 ;
      VIA 14.95 133.28 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 133.095 15.72 133.465 ;
      VIA 14.95 133.28 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 133.28 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 127.675 15.74 128.005 ;
      VIA 14.95 127.84 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 127.655 15.72 128.025 ;
      VIA 14.95 127.84 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 127.84 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 122.235 15.74 122.565 ;
      VIA 14.95 122.4 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 122.215 15.72 122.585 ;
      VIA 14.95 122.4 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 122.4 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 116.795 15.74 117.125 ;
      VIA 14.95 116.96 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 116.775 15.72 117.145 ;
      VIA 14.95 116.96 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 116.96 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 111.355 15.74 111.685 ;
      VIA 14.95 111.52 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 111.335 15.72 111.705 ;
      VIA 14.95 111.52 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 111.52 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 105.915 15.74 106.245 ;
      VIA 14.95 106.08 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 105.895 15.72 106.265 ;
      VIA 14.95 106.08 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 106.08 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 100.475 15.74 100.805 ;
      VIA 14.95 100.64 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 100.455 15.72 100.825 ;
      VIA 14.95 100.64 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 100.64 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 95.035 15.74 95.365 ;
      VIA 14.95 95.2 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 95.015 15.72 95.385 ;
      VIA 14.95 95.2 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 95.2 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 89.595 15.74 89.925 ;
      VIA 14.95 89.76 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 89.575 15.72 89.945 ;
      VIA 14.95 89.76 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 89.76 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 84.155 15.74 84.485 ;
      VIA 14.95 84.32 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 84.135 15.72 84.505 ;
      VIA 14.95 84.32 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 84.32 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 78.715 15.74 79.045 ;
      VIA 14.95 78.88 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 78.695 15.72 79.065 ;
      VIA 14.95 78.88 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 78.88 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 73.275 15.74 73.605 ;
      VIA 14.95 73.44 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 73.255 15.72 73.625 ;
      VIA 14.95 73.44 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 73.44 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 67.835 15.74 68.165 ;
      VIA 14.95 68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 67.815 15.72 68.185 ;
      VIA 14.95 68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 62.395 15.74 62.725 ;
      VIA 14.95 62.56 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 62.375 15.72 62.745 ;
      VIA 14.95 62.56 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 62.56 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 56.955 15.74 57.285 ;
      VIA 14.95 57.12 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 56.935 15.72 57.305 ;
      VIA 14.95 57.12 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 57.12 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 51.515 15.74 51.845 ;
      VIA 14.95 51.68 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 51.495 15.72 51.865 ;
      VIA 14.95 51.68 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 51.68 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 46.075 15.74 46.405 ;
      VIA 14.95 46.24 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 46.055 15.72 46.425 ;
      VIA 14.95 46.24 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 46.24 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 40.635 15.74 40.965 ;
      VIA 14.95 40.8 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 40.615 15.72 40.985 ;
      VIA 14.95 40.8 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 40.8 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 35.195 15.74 35.525 ;
      VIA 14.95 35.36 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 35.175 15.72 35.545 ;
      VIA 14.95 35.36 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 35.36 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 29.755 15.74 30.085 ;
      VIA 14.95 29.92 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 29.735 15.72 30.105 ;
      VIA 14.95 29.92 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 29.92 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 24.315 15.74 24.645 ;
      VIA 14.95 24.48 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 24.295 15.72 24.665 ;
      VIA 14.95 24.48 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 24.48 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 18.875 15.74 19.205 ;
      VIA 14.95 19.04 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 18.855 15.72 19.225 ;
      VIA 14.95 19.04 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 19.04 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 13.435 15.74 13.765 ;
      VIA 14.95 13.6 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 13.415 15.72 13.785 ;
      VIA 14.95 13.6 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 13.6 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 7.995 15.74 8.325 ;
      VIA 14.95 8.16 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 7.975 15.72 8.345 ;
      VIA 14.95 8.16 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 8.16 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 2.555 15.74 2.885 ;
      VIA 14.95 2.72 ibex_if_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 2.535 15.72 2.905 ;
      VIA 14.95 2.72 ibex_if_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 2.72 ibex_if_stage_via2_3_1600_480_1_5_320_320 ;
    END
  END VSS
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.26 0 16.4 0.485 ;
    END
  END boot_addr_i[0]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 202.15 0.8 202.45 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  50.76 295.735 50.9 296.22 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  262.36 295.735 262.5 296.22 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.56 295.735 64.7 296.22 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  230.16 295.735 230.3 296.22 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.06 295.735 99.2 296.22 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.06 295.735 7.2 296.22 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  283.06 295.735 283.2 296.22 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  269.26 295.735 269.4 296.22 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  168.06 295.735 168.2 296.22 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  30.06 0 30.2 0.485 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.96 295.735 152.1 296.22 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  32.36 295.735 32.5 296.22 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 295.735 27.9 296.22 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  225.56 295.735 225.7 296.22 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  96.76 295.735 96.9 296.22 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  172.66 295.735 172.8 296.22 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  78.36 295.735 78.5 296.22 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  46.16 295.735 46.3 296.22 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 259.27 0.8 259.57 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.96 295.735 14.1 296.22 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 0 18.7 0.485 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  163.46 295.735 163.6 296.22 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  289.96 295.735 290.1 296.22 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  200.26 0 200.4 0.485 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.66 0 11.8 0.485 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.96 0 14.1 0.485 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  32.36 0 32.5 0.485 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  41.56 0 41.7 0.485 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 193.99 0.8 194.29 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 196.03 0.8 196.33 ;
    END
  END boot_addr_i[9]
  PIN branch_target_ex_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 0 37.1 0.485 ;
    END
  END branch_target_ex_i[0]
  PIN branch_target_ex_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 206.23 0.8 206.53 ;
    END
  END branch_target_ex_i[10]
  PIN branch_target_ex_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  55.36 295.735 55.5 296.22 ;
    END
  END branch_target_ex_i[11]
  PIN branch_target_ex_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  154.26 295.735 154.4 296.22 ;
    END
  END branch_target_ex_i[12]
  PIN branch_target_ex_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  43.86 295.735 44 296.22 ;
    END
  END branch_target_ex_i[13]
  PIN branch_target_ex_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  253.16 295.735 253.3 296.22 ;
    END
  END branch_target_ex_i[14]
  PIN branch_target_ex_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  207.16 295.735 207.3 296.22 ;
    END
  END branch_target_ex_i[15]
  PIN branch_target_ex_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  271.56 295.735 271.7 296.22 ;
    END
  END branch_target_ex_i[16]
  PIN branch_target_ex_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  260.06 295.735 260.2 296.22 ;
    END
  END branch_target_ex_i[17]
  PIN branch_target_ex_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 214.39 0.8 214.69 ;
    END
  END branch_target_ex_i[18]
  PIN branch_target_ex_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140.46 295.735 140.6 296.22 ;
    END
  END branch_target_ex_i[19]
  PIN branch_target_ex_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  248.56 295.735 248.7 296.22 ;
    END
  END branch_target_ex_i[1]
  PIN branch_target_ex_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.96 295.735 83.1 296.22 ;
    END
  END branch_target_ex_i[20]
  PIN branch_target_ex_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 232.75 0.8 233.05 ;
    END
  END branch_target_ex_i[21]
  PIN branch_target_ex_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  34.66 295.735 34.8 296.22 ;
    END
  END branch_target_ex_i[22]
  PIN branch_target_ex_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  128.96 295.735 129.1 296.22 ;
    END
  END branch_target_ex_i[23]
  PIN branch_target_ex_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.16 295.735 92.3 296.22 ;
    END
  END branch_target_ex_i[24]
  PIN branch_target_ex_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 295.735 73.9 296.22 ;
    END
  END branch_target_ex_i[25]
  PIN branch_target_ex_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  214.06 295.735 214.2 296.22 ;
    END
  END branch_target_ex_i[26]
  PIN branch_target_ex_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  39.26 295.735 39.4 296.22 ;
    END
  END branch_target_ex_i[27]
  PIN branch_target_ex_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.86 295.735 21 296.22 ;
    END
  END branch_target_ex_i[28]
  PIN branch_target_ex_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 238.87 0.8 239.17 ;
    END
  END branch_target_ex_i[29]
  PIN branch_target_ex_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  110.56 295.735 110.7 296.22 ;
    END
  END branch_target_ex_i[2]
  PIN branch_target_ex_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  191.06 295.735 191.2 296.22 ;
    END
  END branch_target_ex_i[30]
  PIN branch_target_ex_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  285.36 295.735 285.5 296.22 ;
    END
  END branch_target_ex_i[31]
  PIN branch_target_ex_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  119.76 295.735 119.9 296.22 ;
    END
  END branch_target_ex_i[3]
  PIN branch_target_ex_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  241.66 295.735 241.8 296.22 ;
    END
  END branch_target_ex_i[4]
  PIN branch_target_ex_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  184.16 295.735 184.3 296.22 ;
    END
  END branch_target_ex_i[5]
  PIN branch_target_ex_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  158.86 295.735 159 296.22 ;
    END
  END branch_target_ex_i[6]
  PIN branch_target_ex_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  179.56 295.735 179.7 296.22 ;
    END
  END branch_target_ex_i[7]
  PIN branch_target_ex_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.26 295.735 108.4 296.22 ;
    END
  END branch_target_ex_i[8]
  PIN branch_target_ex_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  177.26 295.735 177.4 296.22 ;
    END
  END branch_target_ex_i[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 271.51 0.8 271.81 ;
    END
  END clk_i
  PIN csr_depc_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  23.16 0 23.3 0.485 ;
    END
  END csr_depc_i[0]
  PIN csr_depc_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  145.06 295.735 145.2 296.22 ;
    END
  END csr_depc_i[10]
  PIN csr_depc_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48.46 295.735 48.6 296.22 ;
    END
  END csr_depc_i[11]
  PIN csr_depc_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 226.63 0.8 226.93 ;
    END
  END csr_depc_i[12]
  PIN csr_depc_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 220.51 0.8 220.81 ;
    END
  END csr_depc_i[13]
  PIN csr_depc_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  131.26 295.735 131.4 296.22 ;
    END
  END csr_depc_i[14]
  PIN csr_depc_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.66 295.735 103.8 296.22 ;
    END
  END csr_depc_i[15]
  PIN csr_depc_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  69.16 295.735 69.3 296.22 ;
    END
  END csr_depc_i[16]
  PIN csr_depc_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  264.66 295.735 264.8 296.22 ;
    END
  END csr_depc_i[17]
  PIN csr_depc_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  218.66 295.735 218.8 296.22 ;
    END
  END csr_depc_i[18]
  PIN csr_depc_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.96 295.735 175.1 296.22 ;
    END
  END csr_depc_i[19]
  PIN csr_depc_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  202.56 295.735 202.7 296.22 ;
    END
  END csr_depc_i[1]
  PIN csr_depc_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  126.66 295.735 126.8 296.22 ;
    END
  END csr_depc_i[20]
  PIN csr_depc_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  23.16 295.735 23.3 296.22 ;
    END
  END csr_depc_i[21]
  PIN csr_depc_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 295.735 37.1 296.22 ;
    END
  END csr_depc_i[22]
  PIN csr_depc_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  195.66 295.735 195.8 296.22 ;
    END
  END csr_depc_i[23]
  PIN csr_depc_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.96 295.735 60.1 296.22 ;
    END
  END csr_depc_i[24]
  PIN csr_depc_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  80.66 295.735 80.8 296.22 ;
    END
  END csr_depc_i[25]
  PIN csr_depc_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  280.76 295.735 280.9 296.22 ;
    END
  END csr_depc_i[26]
  PIN csr_depc_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  41.56 295.735 41.7 296.22 ;
    END
  END csr_depc_i[27]
  PIN csr_depc_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 257.23 0.8 257.53 ;
    END
  END csr_depc_i[28]
  PIN csr_depc_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 249.07 0.8 249.37 ;
    END
  END csr_depc_i[29]
  PIN csr_depc_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  188.76 295.735 188.9 296.22 ;
    END
  END csr_depc_i[2]
  PIN csr_depc_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  89.86 295.735 90 296.22 ;
    END
  END csr_depc_i[30]
  PIN csr_depc_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  227.86 295.735 228 296.22 ;
    END
  END csr_depc_i[31]
  PIN csr_depc_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  133.56 295.735 133.7 296.22 ;
    END
  END csr_depc_i[3]
  PIN csr_depc_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  250.86 295.735 251 296.22 ;
    END
  END csr_depc_i[4]
  PIN csr_depc_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  246.26 295.735 246.4 296.22 ;
    END
  END csr_depc_i[5]
  PIN csr_depc_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  161.16 295.735 161.3 296.22 ;
    END
  END csr_depc_i[6]
  PIN csr_depc_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  156.56 295.735 156.7 296.22 ;
    END
  END csr_depc_i[7]
  PIN csr_depc_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  216.36 295.735 216.5 296.22 ;
    END
  END csr_depc_i[8]
  PIN csr_depc_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  138.16 295.735 138.3 296.22 ;
    END
  END csr_depc_i[9]
  PIN csr_mepc_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.46 0 25.6 0.485 ;
    END
  END csr_mepc_i[0]
  PIN csr_mepc_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 208.27 0.8 208.57 ;
    END
  END csr_mepc_i[10]
  PIN csr_mepc_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.26 295.735 16.4 296.22 ;
    END
  END csr_mepc_i[11]
  PIN csr_mepc_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  237.06 295.735 237.2 296.22 ;
    END
  END csr_mepc_i[12]
  PIN csr_mepc_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 295.735 9.5 296.22 ;
    END
  END csr_mepc_i[13]
  PIN csr_mepc_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  243.96 295.735 244.1 296.22 ;
    END
  END csr_mepc_i[14]
  PIN csr_mepc_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  149.66 295.735 149.8 296.22 ;
    END
  END csr_mepc_i[15]
  PIN csr_mepc_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  53.06 295.735 53.2 296.22 ;
    END
  END csr_mepc_i[16]
  PIN csr_mepc_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  204.86 295.735 205 296.22 ;
    END
  END csr_mepc_i[17]
  PIN csr_mepc_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 212.35 0.8 212.65 ;
    END
  END csr_mepc_i[18]
  PIN csr_mepc_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  200.26 295.735 200.4 296.22 ;
    END
  END csr_mepc_i[19]
  PIN csr_mepc_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  255.46 295.735 255.6 296.22 ;
    END
  END csr_mepc_i[1]
  PIN csr_mepc_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  197.96 295.735 198.1 296.22 ;
    END
  END csr_mepc_i[20]
  PIN csr_mepc_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 234.79 0.8 235.09 ;
    END
  END csr_mepc_i[21]
  PIN csr_mepc_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  4.76 295.735 4.9 296.22 ;
    END
  END csr_mepc_i[22]
  PIN csr_mepc_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  135.86 295.735 136 296.22 ;
    END
  END csr_mepc_i[23]
  PIN csr_mepc_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94.46 295.735 94.6 296.22 ;
    END
  END csr_mepc_i[24]
  PIN csr_mepc_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71.46 295.735 71.6 296.22 ;
    END
  END csr_mepc_i[25]
  PIN csr_mepc_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  76.06 295.735 76.2 296.22 ;
    END
  END csr_mepc_i[26]
  PIN csr_mepc_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.66 295.735 11.8 296.22 ;
    END
  END csr_mepc_i[27]
  PIN csr_mepc_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 295.735 18.7 296.22 ;
    END
  END csr_mepc_i[28]
  PIN csr_mepc_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 242.95 0.8 243.25 ;
    END
  END csr_mepc_i[29]
  PIN csr_mepc_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  165.76 295.735 165.9 296.22 ;
    END
  END csr_mepc_i[2]
  PIN csr_mepc_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  85.26 295.735 85.4 296.22 ;
    END
  END csr_mepc_i[30]
  PIN csr_mepc_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  273.86 295.735 274 296.22 ;
    END
  END csr_mepc_i[31]
  PIN csr_mepc_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  257.76 295.735 257.9 296.22 ;
    END
  END csr_mepc_i[3]
  PIN csr_mepc_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  266.96 295.735 267.1 296.22 ;
    END
  END csr_mepc_i[4]
  PIN csr_mepc_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  124.36 295.735 124.5 296.22 ;
    END
  END csr_mepc_i[5]
  PIN csr_mepc_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  276.16 295.735 276.3 296.22 ;
    END
  END csr_mepc_i[6]
  PIN csr_mepc_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.86 295.735 113 296.22 ;
    END
  END csr_mepc_i[7]
  PIN csr_mepc_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  193.36 295.735 193.5 296.22 ;
    END
  END csr_mepc_i[8]
  PIN csr_mepc_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  115.16 295.735 115.3 296.22 ;
    END
  END csr_mepc_i[9]
  PIN csr_mtvec_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.96 0 60.1 0.485 ;
    END
  END csr_mtvec_i[0]
  PIN csr_mtvec_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  87.56 295.735 87.7 296.22 ;
    END
  END csr_mtvec_i[10]
  PIN csr_mtvec_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  57.66 295.735 57.8 296.22 ;
    END
  END csr_mtvec_i[11]
  PIN csr_mtvec_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 216.43 0.8 216.73 ;
    END
  END csr_mtvec_i[12]
  PIN csr_mtvec_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 218.47 0.8 218.77 ;
    END
  END csr_mtvec_i[13]
  PIN csr_mtvec_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  211.76 295.735 211.9 296.22 ;
    END
  END csr_mtvec_i[14]
  PIN csr_mtvec_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  105.96 295.735 106.1 296.22 ;
    END
  END csr_mtvec_i[15]
  PIN csr_mtvec_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  62.26 295.735 62.4 296.22 ;
    END
  END csr_mtvec_i[16]
  PIN csr_mtvec_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  234.76 295.735 234.9 296.22 ;
    END
  END csr_mtvec_i[17]
  PIN csr_mtvec_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  117.46 295.735 117.6 296.22 ;
    END
  END csr_mtvec_i[18]
  PIN csr_mtvec_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  181.86 295.735 182 296.22 ;
    END
  END csr_mtvec_i[19]
  PIN csr_mtvec_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  39.26 0 39.4 0.485 ;
    END
  END csr_mtvec_i[1]
  PIN csr_mtvec_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  186.46 295.735 186.6 296.22 ;
    END
  END csr_mtvec_i[20]
  PIN csr_mtvec_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 230.71 0.8 231.01 ;
    END
  END csr_mtvec_i[21]
  PIN csr_mtvec_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2.46 295.735 2.6 296.22 ;
    END
  END csr_mtvec_i[22]
  PIN csr_mtvec_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  170.36 295.735 170.5 296.22 ;
    END
  END csr_mtvec_i[23]
  PIN csr_mtvec_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  287.66 295.735 287.8 296.22 ;
    END
  END csr_mtvec_i[24]
  PIN csr_mtvec_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  232.46 295.735 232.6 296.22 ;
    END
  END csr_mtvec_i[25]
  PIN csr_mtvec_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.86 295.735 67 296.22 ;
    END
  END csr_mtvec_i[26]
  PIN csr_mtvec_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.46 295.735 25.6 296.22 ;
    END
  END csr_mtvec_i[27]
  PIN csr_mtvec_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  30.06 295.735 30.2 296.22 ;
    END
  END csr_mtvec_i[28]
  PIN csr_mtvec_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 240.91 0.8 241.21 ;
    END
  END csr_mtvec_i[29]
  PIN csr_mtvec_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  43.86 0 44 0.485 ;
    END
  END csr_mtvec_i[2]
  PIN csr_mtvec_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  147.36 295.735 147.5 296.22 ;
    END
  END csr_mtvec_i[30]
  PIN csr_mtvec_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  122.06 295.735 122.2 296.22 ;
    END
  END csr_mtvec_i[31]
  PIN csr_mtvec_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  34.66 0 34.8 0.485 ;
    END
  END csr_mtvec_i[3]
  PIN csr_mtvec_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  53.06 0 53.2 0.485 ;
    END
  END csr_mtvec_i[4]
  PIN csr_mtvec_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  188.76 0 188.9 0.485 ;
    END
  END csr_mtvec_i[5]
  PIN csr_mtvec_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  202.56 0 202.7 0.485 ;
    END
  END csr_mtvec_i[6]
  PIN csr_mtvec_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48.46 0 48.6 0.485 ;
    END
  END csr_mtvec_i[7]
  PIN csr_mtvec_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  239.36 295.735 239.5 296.22 ;
    END
  END csr_mtvec_i[8]
  PIN csr_mtvec_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  223.26 295.735 223.4 296.22 ;
    END
  END csr_mtvec_i[9]
  PIN csr_mtvec_init_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  101.36 295.735 101.5 296.22 ;
    END
  END csr_mtvec_init_o
  PIN dummy_instr_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  46.16 0 46.3 0.485 ;
    END
  END dummy_instr_en_i
  PIN dummy_instr_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 77.71 0.8 78.01 ;
    END
  END dummy_instr_id_o
  PIN dummy_instr_mask_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  126.66 0 126.8 0.485 ;
    END
  END dummy_instr_mask_i[0]
  PIN dummy_instr_mask_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  207.16 0 207.3 0.485 ;
    END
  END dummy_instr_mask_i[1]
  PIN dummy_instr_mask_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  69.16 0 69.3 0.485 ;
    END
  END dummy_instr_mask_i[2]
  PIN dummy_instr_seed_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  55.36 0 55.5 0.485 ;
    END
  END dummy_instr_seed_en_i
  PIN dummy_instr_seed_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  57.66 0 57.8 0.485 ;
    END
  END dummy_instr_seed_i[0]
  PIN dummy_instr_seed_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.96 0 83.1 0.485 ;
    END
  END dummy_instr_seed_i[10]
  PIN dummy_instr_seed_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  62.26 0 62.4 0.485 ;
    END
  END dummy_instr_seed_i[11]
  PIN dummy_instr_seed_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.56 0 64.7 0.485 ;
    END
  END dummy_instr_seed_i[12]
  PIN dummy_instr_seed_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.86 0 67 0.485 ;
    END
  END dummy_instr_seed_i[13]
  PIN dummy_instr_seed_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  85.26 0 85.4 0.485 ;
    END
  END dummy_instr_seed_i[14]
  PIN dummy_instr_seed_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71.46 0 71.6 0.485 ;
    END
  END dummy_instr_seed_i[15]
  PIN dummy_instr_seed_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 0 73.9 0.485 ;
    END
  END dummy_instr_seed_i[16]
  PIN dummy_instr_seed_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  76.06 0 76.2 0.485 ;
    END
  END dummy_instr_seed_i[17]
  PIN dummy_instr_seed_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  78.36 0 78.5 0.485 ;
    END
  END dummy_instr_seed_i[18]
  PIN dummy_instr_seed_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  80.66 0 80.8 0.485 ;
    END
  END dummy_instr_seed_i[19]
  PIN dummy_instr_seed_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.26 0 108.4 0.485 ;
    END
  END dummy_instr_seed_i[1]
  PIN dummy_instr_seed_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  119.76 0 119.9 0.485 ;
    END
  END dummy_instr_seed_i[20]
  PIN dummy_instr_seed_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  87.56 0 87.7 0.485 ;
    END
  END dummy_instr_seed_i[21]
  PIN dummy_instr_seed_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  193.36 0 193.5 0.485 ;
    END
  END dummy_instr_seed_i[22]
  PIN dummy_instr_seed_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.16 0 92.3 0.485 ;
    END
  END dummy_instr_seed_i[23]
  PIN dummy_instr_seed_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94.46 0 94.6 0.485 ;
    END
  END dummy_instr_seed_i[24]
  PIN dummy_instr_seed_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  96.76 0 96.9 0.485 ;
    END
  END dummy_instr_seed_i[25]
  PIN dummy_instr_seed_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  4.76 0 4.9 0.485 ;
    END
  END dummy_instr_seed_i[26]
  PIN dummy_instr_seed_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  101.36 0 101.5 0.485 ;
    END
  END dummy_instr_seed_i[27]
  PIN dummy_instr_seed_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 0 27.9 0.485 ;
    END
  END dummy_instr_seed_i[28]
  PIN dummy_instr_seed_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.86 0 21 0.485 ;
    END
  END dummy_instr_seed_i[29]
  PIN dummy_instr_seed_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  211.76 0 211.9 0.485 ;
    END
  END dummy_instr_seed_i[2]
  PIN dummy_instr_seed_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  110.56 0 110.7 0.485 ;
    END
  END dummy_instr_seed_i[30]
  PIN dummy_instr_seed_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.96 0 175.1 0.485 ;
    END
  END dummy_instr_seed_i[31]
  PIN dummy_instr_seed_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  115.16 0 115.3 0.485 ;
    END
  END dummy_instr_seed_i[3]
  PIN dummy_instr_seed_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.06 0 7.2 0.485 ;
    END
  END dummy_instr_seed_i[4]
  PIN dummy_instr_seed_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2.46 0 2.6 0.485 ;
    END
  END dummy_instr_seed_i[5]
  PIN dummy_instr_seed_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  122.06 0 122.2 0.485 ;
    END
  END dummy_instr_seed_i[6]
  PIN dummy_instr_seed_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  177.26 0 177.4 0.485 ;
    END
  END dummy_instr_seed_i[7]
  PIN dummy_instr_seed_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  204.86 0 205 0.485 ;
    END
  END dummy_instr_seed_i[8]
  PIN dummy_instr_seed_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  128.96 0 129.1 0.485 ;
    END
  END dummy_instr_seed_i[9]
  PIN exc_cause[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  209.46 295.735 209.6 296.22 ;
    END
  END exc_cause[0]
  PIN exc_cause[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  142.76 295.735 142.9 296.22 ;
    END
  END exc_cause[1]
  PIN exc_cause[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 183.79 0.8 184.09 ;
    END
  END exc_cause[2]
  PIN exc_cause[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  278.46 295.735 278.6 296.22 ;
    END
  END exc_cause[3]
  PIN exc_cause[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  220.96 295.735 221.1 296.22 ;
    END
  END exc_cause[4]
  PIN exc_cause[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 0 9.5 0.485 ;
    END
  END exc_cause[5]
  PIN exc_pc_mux_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  292.26 295.735 292.4 296.22 ;
    END
  END exc_pc_mux_i[0]
  PIN exc_pc_mux_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 255.19 0.8 255.49 ;
    END
  END exc_pc_mux_i[1]
  PIN icache_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  197.96 0 198.1 0.485 ;
    END
  END icache_enable_i
  PIN icache_inval_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  50.76 0 50.9 0.485 ;
    END
  END icache_inval_i
  PIN id_in_ready_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  124.36 0 124.5 0.485 ;
    END
  END id_in_ready_i
  PIN if_busy_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 91.99 0.8 92.29 ;
    END
  END if_busy_o
  PIN illegal_c_insn_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 291.91 296.22 292.21 ;
    END
  END illegal_c_insn_id_o
  PIN instr_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 87.91 0.8 88.21 ;
    END
  END instr_addr_o[0]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 136.87 0.8 137.17 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 100.15 0.8 100.45 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 106.27 0.8 106.57 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 122.59 0.8 122.89 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 114.43 0.8 114.73 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 102.19 0.8 102.49 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 126.67 0.8 126.97 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 108.31 0.8 108.61 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 130.75 0.8 131.05 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 132.79 0.8 133.09 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 85.87 0.8 86.17 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 118.51 0.8 118.81 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 167.47 0.8 167.77 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 116.47 0.8 116.77 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 112.39 0.8 112.69 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 145.03 0.8 145.33 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 155.23 0.8 155.53 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 157.27 0.8 157.57 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 110.35 0.8 110.65 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 151.15 0.8 151.45 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 161.35 0.8 161.65 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 163.39 0.8 163.69 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 153.19 0.8 153.49 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 159.31 0.8 159.61 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 120.55 0.8 120.85 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 142.99 0.8 143.29 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 134.83 0.8 135.13 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 147.07 0.8 147.37 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 140.95 0.8 141.25 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 128.71 0.8 129.01 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 165.43 0.8 165.73 ;
    END
  END instr_addr_o[9]
  PIN instr_bp_taken_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 79.75 0.8 80.05 ;
    END
  END instr_bp_taken_o
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  117.46 0 117.6 0.485 ;
    END
  END instr_err_i
  PIN instr_fetch_err_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  138.16 0 138.3 0.485 ;
    END
  END instr_fetch_err_o
  PIN instr_fetch_err_plus2_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  133.56 0 133.7 0.485 ;
    END
  END instr_fetch_err_plus2_o
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 96.07 0.8 96.37 ;
    END
  END instr_gnt_i
  PIN instr_is_compressed_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 32.83 296.22 33.13 ;
    END
  END instr_is_compressed_id_o
  PIN instr_new_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  135.86 0 136 0.485 ;
    END
  END instr_new_id_o
  PIN instr_pmp_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 94.03 0.8 94.33 ;
    END
  END instr_pmp_err_i
  PIN instr_rdata_alu_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 69.55 296.22 69.85 ;
    END
  END instr_rdata_alu_id_o[0]
  PIN instr_rdata_alu_id_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 289.87 296.22 290.17 ;
    END
  END instr_rdata_alu_id_o[10]
  PIN instr_rdata_alu_id_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 287.83 296.22 288.13 ;
    END
  END instr_rdata_alu_id_o[11]
  PIN instr_rdata_alu_id_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 55.27 296.22 55.57 ;
    END
  END instr_rdata_alu_id_o[12]
  PIN instr_rdata_alu_id_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 200.11 296.22 200.41 ;
    END
  END instr_rdata_alu_id_o[13]
  PIN instr_rdata_alu_id_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 71.59 296.22 71.89 ;
    END
  END instr_rdata_alu_id_o[14]
  PIN instr_rdata_alu_id_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 196.03 296.22 196.33 ;
    END
  END instr_rdata_alu_id_o[15]
  PIN instr_rdata_alu_id_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 136.87 296.22 137.17 ;
    END
  END instr_rdata_alu_id_o[16]
  PIN instr_rdata_alu_id_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 132.79 296.22 133.09 ;
    END
  END instr_rdata_alu_id_o[17]
  PIN instr_rdata_alu_id_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 126.67 296.22 126.97 ;
    END
  END instr_rdata_alu_id_o[18]
  PIN instr_rdata_alu_id_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 147.07 296.22 147.37 ;
    END
  END instr_rdata_alu_id_o[19]
  PIN instr_rdata_alu_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 242.95 296.22 243.25 ;
    END
  END instr_rdata_alu_id_o[1]
  PIN instr_rdata_alu_id_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  158.86 0 159 0.485 ;
    END
  END instr_rdata_alu_id_o[20]
  PIN instr_rdata_alu_id_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 124.63 296.22 124.93 ;
    END
  END instr_rdata_alu_id_o[21]
  PIN instr_rdata_alu_id_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 116.47 296.22 116.77 ;
    END
  END instr_rdata_alu_id_o[22]
  PIN instr_rdata_alu_id_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 98.11 296.22 98.41 ;
    END
  END instr_rdata_alu_id_o[23]
  PIN instr_rdata_alu_id_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 120.55 296.22 120.85 ;
    END
  END instr_rdata_alu_id_o[24]
  PIN instr_rdata_alu_id_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 114.43 296.22 114.73 ;
    END
  END instr_rdata_alu_id_o[25]
  PIN instr_rdata_alu_id_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 102.19 296.22 102.49 ;
    END
  END instr_rdata_alu_id_o[26]
  PIN instr_rdata_alu_id_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 73.63 296.22 73.93 ;
    END
  END instr_rdata_alu_id_o[27]
  PIN instr_rdata_alu_id_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 85.87 296.22 86.17 ;
    END
  END instr_rdata_alu_id_o[28]
  PIN instr_rdata_alu_id_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 77.71 296.22 78.01 ;
    END
  END instr_rdata_alu_id_o[29]
  PIN instr_rdata_alu_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 204.19 296.22 204.49 ;
    END
  END instr_rdata_alu_id_o[2]
  PIN instr_rdata_alu_id_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 87.91 296.22 88.21 ;
    END
  END instr_rdata_alu_id_o[30]
  PIN instr_rdata_alu_id_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 79.75 296.22 80.05 ;
    END
  END instr_rdata_alu_id_o[31]
  PIN instr_rdata_alu_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 63.43 296.22 63.73 ;
    END
  END instr_rdata_alu_id_o[3]
  PIN instr_rdata_alu_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 198.07 296.22 198.37 ;
    END
  END instr_rdata_alu_id_o[4]
  PIN instr_rdata_alu_id_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 57.31 296.22 57.61 ;
    END
  END instr_rdata_alu_id_o[5]
  PIN instr_rdata_alu_id_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 157.27 296.22 157.57 ;
    END
  END instr_rdata_alu_id_o[6]
  PIN instr_rdata_alu_id_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 34.87 296.22 35.17 ;
    END
  END instr_rdata_alu_id_o[7]
  PIN instr_rdata_alu_id_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 226.63 296.22 226.93 ;
    END
  END instr_rdata_alu_id_o[8]
  PIN instr_rdata_alu_id_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 47.11 296.22 47.41 ;
    END
  END instr_rdata_alu_id_o[9]
  PIN instr_rdata_c_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 36.91 296.22 37.21 ;
    END
  END instr_rdata_c_id_o[0]
  PIN instr_rdata_c_id_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 43.03 296.22 43.33 ;
    END
  END instr_rdata_c_id_o[10]
  PIN instr_rdata_c_id_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 53.23 296.22 53.53 ;
    END
  END instr_rdata_c_id_o[11]
  PIN instr_rdata_c_id_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 104.23 296.22 104.53 ;
    END
  END instr_rdata_c_id_o[12]
  PIN instr_rdata_c_id_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 183.79 296.22 184.09 ;
    END
  END instr_rdata_c_id_o[13]
  PIN instr_rdata_c_id_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 173.59 296.22 173.89 ;
    END
  END instr_rdata_c_id_o[14]
  PIN instr_rdata_c_id_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 40.99 296.22 41.29 ;
    END
  END instr_rdata_c_id_o[15]
  PIN instr_rdata_c_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 175.63 296.22 175.93 ;
    END
  END instr_rdata_c_id_o[1]
  PIN instr_rdata_c_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 167.47 296.22 167.77 ;
    END
  END instr_rdata_c_id_o[2]
  PIN instr_rdata_c_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 67.51 296.22 67.81 ;
    END
  END instr_rdata_c_id_o[3]
  PIN instr_rdata_c_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 149.11 296.22 149.41 ;
    END
  END instr_rdata_c_id_o[4]
  PIN instr_rdata_c_id_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 138.91 296.22 139.21 ;
    END
  END instr_rdata_c_id_o[5]
  PIN instr_rdata_c_id_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 130.75 296.22 131.05 ;
    END
  END instr_rdata_c_id_o[6]
  PIN instr_rdata_c_id_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 179.71 296.22 180.01 ;
    END
  END instr_rdata_c_id_o[7]
  PIN instr_rdata_c_id_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 285.79 296.22 286.09 ;
    END
  END instr_rdata_c_id_o[8]
  PIN instr_rdata_c_id_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 81.79 296.22 82.09 ;
    END
  END instr_rdata_c_id_o[9]
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.06 0 99.2 0.485 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  181.86 0 182 0.485 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  184.16 0 184.3 0.485 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 75.67 296.22 75.97 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 45.07 296.22 45.37 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  195.66 0 195.8 0.485 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  214.06 0 214.2 0.485 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  105.96 0 106.1 0.485 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.86 0 113 0.485 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  142.76 0 142.9 0.485 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  145.06 0 145.2 0.485 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.66 0 103.8 0.485 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  149.66 0 149.8 0.485 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.96 0 152.1 0.485 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  179.56 0 179.7 0.485 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  216.36 0 216.5 0.485 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  163.46 0 163.6 0.485 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  191.06 0 191.2 0.485 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  168.06 0 168.2 0.485 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  186.46 0 186.6 0.485 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  246.26 0 246.4 0.485 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  248.56 0 248.7 0.485 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140.46 0 140.6 0.485 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  209.46 0 209.6 0.485 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  227.86 0 228 0.485 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  154.26 0 154.4 0.485 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  156.56 0 156.7 0.485 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  165.76 0 165.9 0.485 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  170.36 0 170.5 0.485 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  225.56 0 225.7 0.485 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  172.66 0 172.8 0.485 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 61.39 296.22 61.69 ;
    END
  END instr_rdata_i[9]
  PIN instr_rdata_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 145.03 296.22 145.33 ;
    END
  END instr_rdata_id_o[0]
  PIN instr_rdata_id_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 216.43 296.22 216.73 ;
    END
  END instr_rdata_id_o[10]
  PIN instr_rdata_id_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 189.91 296.22 190.21 ;
    END
  END instr_rdata_id_o[11]
  PIN instr_rdata_id_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 159.31 296.22 159.61 ;
    END
  END instr_rdata_id_o[12]
  PIN instr_rdata_id_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 191.95 296.22 192.25 ;
    END
  END instr_rdata_id_o[13]
  PIN instr_rdata_id_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 110.35 296.22 110.65 ;
    END
  END instr_rdata_id_o[14]
  PIN instr_rdata_id_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 202.15 296.22 202.45 ;
    END
  END instr_rdata_id_o[15]
  PIN instr_rdata_id_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 140.95 296.22 141.25 ;
    END
  END instr_rdata_id_o[16]
  PIN instr_rdata_id_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 128.71 296.22 129.01 ;
    END
  END instr_rdata_id_o[17]
  PIN instr_rdata_id_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 100.15 296.22 100.45 ;
    END
  END instr_rdata_id_o[18]
  PIN instr_rdata_id_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 65.47 296.22 65.77 ;
    END
  END instr_rdata_id_o[19]
  PIN instr_rdata_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 259.27 296.22 259.57 ;
    END
  END instr_rdata_id_o[1]
  PIN instr_rdata_id_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  161.16 0 161.3 0.485 ;
    END
  END instr_rdata_id_o[20]
  PIN instr_rdata_id_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 108.31 296.22 108.61 ;
    END
  END instr_rdata_id_o[21]
  PIN instr_rdata_id_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 118.51 296.22 118.81 ;
    END
  END instr_rdata_id_o[22]
  PIN instr_rdata_id_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 134.83 296.22 135.13 ;
    END
  END instr_rdata_id_o[23]
  PIN instr_rdata_id_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 122.59 296.22 122.89 ;
    END
  END instr_rdata_id_o[24]
  PIN instr_rdata_id_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 112.39 296.22 112.69 ;
    END
  END instr_rdata_id_o[25]
  PIN instr_rdata_id_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 106.27 296.22 106.57 ;
    END
  END instr_rdata_id_o[26]
  PIN instr_rdata_id_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 94.03 296.22 94.33 ;
    END
  END instr_rdata_id_o[27]
  PIN instr_rdata_id_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 91.99 296.22 92.29 ;
    END
  END instr_rdata_id_o[28]
  PIN instr_rdata_id_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 96.07 296.22 96.37 ;
    END
  END instr_rdata_id_o[29]
  PIN instr_rdata_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 206.23 296.22 206.53 ;
    END
  END instr_rdata_id_o[2]
  PIN instr_rdata_id_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 89.95 296.22 90.25 ;
    END
  END instr_rdata_id_o[30]
  PIN instr_rdata_id_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 83.83 296.22 84.13 ;
    END
  END instr_rdata_id_o[31]
  PIN instr_rdata_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 59.35 296.22 59.65 ;
    END
  END instr_rdata_id_o[3]
  PIN instr_rdata_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 269.47 296.22 269.77 ;
    END
  END instr_rdata_id_o[4]
  PIN instr_rdata_id_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 153.19 296.22 153.49 ;
    END
  END instr_rdata_id_o[5]
  PIN instr_rdata_id_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 155.23 296.22 155.53 ;
    END
  END instr_rdata_id_o[6]
  PIN instr_rdata_id_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 181.75 296.22 182.05 ;
    END
  END instr_rdata_id_o[7]
  PIN instr_rdata_id_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 222.55 296.22 222.85 ;
    END
  END instr_rdata_id_o[8]
  PIN instr_rdata_id_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 161.35 296.22 161.65 ;
    END
  END instr_rdata_id_o[9]
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 98.11 0.8 98.41 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  89.86 0 90 0.485 ;
    END
  END instr_rvalid_i
  PIN instr_valid_clear_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 138.91 0.8 139.21 ;
    END
  END instr_valid_clear_i
  PIN instr_valid_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 124.63 0.8 124.93 ;
    END
  END instr_valid_id_o
  PIN nt_branch_mispredict_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 189.91 0.8 190.21 ;
    END
  END nt_branch_mispredict_i
  PIN pc_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 83.83 0.8 84.13 ;
    END
  END pc_id_o[0]
  PIN pc_id_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 212.35 296.22 212.65 ;
    END
  END pc_id_o[10]
  PIN pc_id_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 228.67 296.22 228.97 ;
    END
  END pc_id_o[11]
  PIN pc_id_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 283.75 296.22 284.05 ;
    END
  END pc_id_o[12]
  PIN pc_id_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 261.31 296.22 261.61 ;
    END
  END pc_id_o[13]
  PIN pc_id_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 230.71 296.22 231.01 ;
    END
  END pc_id_o[14]
  PIN pc_id_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 240.91 296.22 241.21 ;
    END
  END pc_id_o[15]
  PIN pc_id_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 210.31 296.22 210.61 ;
    END
  END pc_id_o[16]
  PIN pc_id_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 275.59 296.22 275.89 ;
    END
  END pc_id_o[17]
  PIN pc_id_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 279.67 0.8 279.97 ;
    END
  END pc_id_o[18]
  PIN pc_id_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 277.63 0.8 277.93 ;
    END
  END pc_id_o[19]
  PIN pc_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  147.36 0 147.5 0.485 ;
    END
  END pc_id_o[1]
  PIN pc_id_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 273.55 0.8 273.85 ;
    END
  END pc_id_o[20]
  PIN pc_id_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 275.59 0.8 275.89 ;
    END
  END pc_id_o[21]
  PIN pc_id_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 281.71 296.22 282.01 ;
    END
  END pc_id_o[22]
  PIN pc_id_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 247.03 296.22 247.33 ;
    END
  END pc_id_o[23]
  PIN pc_id_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 257.23 296.22 257.53 ;
    END
  END pc_id_o[24]
  PIN pc_id_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 255.19 296.22 255.49 ;
    END
  END pc_id_o[25]
  PIN pc_id_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 267.43 296.22 267.73 ;
    END
  END pc_id_o[26]
  PIN pc_id_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 273.55 296.22 273.85 ;
    END
  END pc_id_o[27]
  PIN pc_id_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 279.67 296.22 279.97 ;
    END
  END pc_id_o[28]
  PIN pc_id_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 238.87 296.22 239.17 ;
    END
  END pc_id_o[29]
  PIN pc_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 142.99 296.22 143.29 ;
    END
  END pc_id_o[2]
  PIN pc_id_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 244.99 296.22 245.29 ;
    END
  END pc_id_o[30]
  PIN pc_id_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 222.55 0.8 222.85 ;
    END
  END pc_id_o[31]
  PIN pc_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 151.15 296.22 151.45 ;
    END
  END pc_id_o[3]
  PIN pc_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 177.67 296.22 177.97 ;
    END
  END pc_id_o[4]
  PIN pc_id_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 165.43 296.22 165.73 ;
    END
  END pc_id_o[5]
  PIN pc_id_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 169.51 296.22 169.81 ;
    END
  END pc_id_o[6]
  PIN pc_id_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 51.19 296.22 51.49 ;
    END
  END pc_id_o[7]
  PIN pc_id_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 187.87 296.22 188.17 ;
    END
  END pc_id_o[8]
  PIN pc_id_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 185.83 296.22 186.13 ;
    END
  END pc_id_o[9]
  PIN pc_if_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 89.95 0.8 90.25 ;
    END
  END pc_if_o[0]
  PIN pc_if_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 263.35 296.22 263.65 ;
    END
  END pc_if_o[10]
  PIN pc_if_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 224.59 296.22 224.89 ;
    END
  END pc_if_o[11]
  PIN pc_if_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 218.47 296.22 218.77 ;
    END
  END pc_if_o[12]
  PIN pc_if_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 220.51 296.22 220.81 ;
    END
  END pc_if_o[13]
  PIN pc_if_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 214.39 296.22 214.69 ;
    END
  END pc_if_o[14]
  PIN pc_if_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 204.19 0.8 204.49 ;
    END
  END pc_if_o[15]
  PIN pc_if_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 234.79 296.22 235.09 ;
    END
  END pc_if_o[16]
  PIN pc_if_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 208.27 296.22 208.57 ;
    END
  END pc_if_o[17]
  PIN pc_if_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 267.43 0.8 267.73 ;
    END
  END pc_if_o[18]
  PIN pc_if_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 265.39 0.8 265.69 ;
    END
  END pc_if_o[19]
  PIN pc_if_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  131.26 0 131.4 0.485 ;
    END
  END pc_if_o[1]
  PIN pc_if_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 269.47 0.8 269.77 ;
    END
  END pc_if_o[20]
  PIN pc_if_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 263.35 0.8 263.65 ;
    END
  END pc_if_o[21]
  PIN pc_if_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 261.31 0.8 261.61 ;
    END
  END pc_if_o[22]
  PIN pc_if_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 249.07 296.22 249.37 ;
    END
  END pc_if_o[23]
  PIN pc_if_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 251.11 296.22 251.41 ;
    END
  END pc_if_o[24]
  PIN pc_if_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 253.15 296.22 253.45 ;
    END
  END pc_if_o[25]
  PIN pc_if_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 265.39 296.22 265.69 ;
    END
  END pc_if_o[26]
  PIN pc_if_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 271.51 296.22 271.81 ;
    END
  END pc_if_o[27]
  PIN pc_if_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 277.63 296.22 277.93 ;
    END
  END pc_if_o[28]
  PIN pc_if_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 236.83 296.22 237.13 ;
    END
  END pc_if_o[29]
  PIN pc_if_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 149.11 0.8 149.41 ;
    END
  END pc_if_o[2]
  PIN pc_if_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 232.75 296.22 233.05 ;
    END
  END pc_if_o[30]
  PIN pc_if_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 224.59 0.8 224.89 ;
    END
  END pc_if_o[31]
  PIN pc_if_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 175.63 0.8 175.93 ;
    END
  END pc_if_o[3]
  PIN pc_if_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 171.55 296.22 171.85 ;
    END
  END pc_if_o[4]
  PIN pc_if_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 163.39 296.22 163.69 ;
    END
  END pc_if_o[5]
  PIN pc_if_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 38.95 296.22 39.25 ;
    END
  END pc_if_o[6]
  PIN pc_if_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 49.15 296.22 49.45 ;
    END
  END pc_if_o[7]
  PIN pc_if_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 187.87 0.8 188.17 ;
    END
  END pc_if_o[8]
  PIN pc_if_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  295.42 193.99 296.22 194.29 ;
    END
  END pc_if_o[9]
  PIN pc_mismatch_alert_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 81.79 0.8 82.09 ;
    END
  END pc_mismatch_alert_o
  PIN pc_mux_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 283.75 0.8 284.05 ;
    END
  END pc_mux_i[0]
  PIN pc_mux_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 287.83 0.8 288.13 ;
    END
  END pc_mux_i[1]
  PIN pc_mux_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 281.71 0.8 282.01 ;
    END
  END pc_mux_i[2]
  PIN pc_set_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 210.31 0.8 210.61 ;
    END
  END pc_set_i
  PIN pc_set_spec_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 181.75 0.8 182.05 ;
    END
  END pc_set_spec_i
  PIN req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 104.23 0.8 104.53 ;
    END
  END req_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 75.67 0.8 75.97 ;
    END
  END rst_ni
  OBS
    LAYER nwell ;
     RECT  0 0 296.22 296.22 ;
    LAYER pwell ;
     RECT  0 0 296.22 296.22 ;
    LAYER li1 ;
     RECT  0 0 296.22 296.22 ;
    LAYER met1 ;
     RECT  0 0 296.22 296.22 ;
    LAYER met2 ;
     RECT  0 0 296.22 296.22 ;
    LAYER met3 ;
     RECT  0 0 296.22 296.22 ;
    LAYER met4 ;
     RECT  0 0 296.22 296.22 ;
    LAYER met5 ;
     RECT  0 0 296.22 296.22 ;
  END
END ibex_if_stage
END LIBRARY
