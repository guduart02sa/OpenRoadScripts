module ibex_wb_stage (clk_i,
    en_wb_i,
    instr_done_wb_o,
    instr_is_compressed_id_i,
    instr_perf_count_id_i,
    lsu_resp_err_i,
    lsu_resp_valid_i,
    outstanding_load_wb_o,
    outstanding_store_wb_o,
    perf_instr_ret_compressed_wb_o,
    perf_instr_ret_wb_o,
    ready_wb_o,
    rf_we_id_i,
    rf_we_lsu_i,
    rf_we_wb_o,
    rf_write_wb_o,
    rst_ni,
    instr_type_wb_i,
    pc_id_i,
    pc_wb_o,
    rf_waddr_id_i,
    rf_waddr_wb_o,
    rf_wdata_fwd_wb_o,
    rf_wdata_id_i,
    rf_wdata_lsu_i,
    rf_wdata_wb_o);
 input clk_i;
 input en_wb_i;
 output instr_done_wb_o;
 input instr_is_compressed_id_i;
 input instr_perf_count_id_i;
 input lsu_resp_err_i;
 input lsu_resp_valid_i;
 output outstanding_load_wb_o;
 output outstanding_store_wb_o;
 output perf_instr_ret_compressed_wb_o;
 output perf_instr_ret_wb_o;
 output ready_wb_o;
 input rf_we_id_i;
 input rf_we_lsu_i;
 output rf_we_wb_o;
 output rf_write_wb_o;
 input rst_ni;
 input [1:0] instr_type_wb_i;
 input [31:0] pc_id_i;
 output [31:0] pc_wb_o;
 input [4:0] rf_waddr_id_i;
 output [4:0] rf_waddr_wb_o;
 output [31:0] rf_wdata_fwd_wb_o;
 input [31:0] rf_wdata_id_i;
 input [31:0] rf_wdata_lsu_i;
 output [31:0] rf_wdata_wb_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire net179;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;

 sky130_fd_sc_hd__nand2_1 _008_ (.A(net1),
    .B(net3),
    .Y(_000_));
 sky130_fd_sc_hd__a21oi_1 _009_ (.A1(net4),
    .A2(net5),
    .B1(_000_),
    .Y(net72));
 sky130_fd_sc_hd__inv_1 _010_ (.A(net2),
    .Y(_001_));
 sky130_fd_sc_hd__a211oi_1 _011_ (.A1(net4),
    .A2(net5),
    .B1(_001_),
    .C1(_000_),
    .Y(net71));
 sky130_fd_sc_hd__buf_6 _012_ (.A(rf_we_id_i),
    .X(_002_));
 sky130_fd_sc_hd__buf_6 _013_ (.A(_002_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _014_ (.A0(net38),
    .A1(net6),
    .S(_003_),
    .X(net78));
 sky130_fd_sc_hd__mux2_1 _015_ (.A0(net39),
    .A1(net7),
    .S(_003_),
    .X(net79));
 sky130_fd_sc_hd__mux2_1 _016_ (.A0(net40),
    .A1(net8),
    .S(_003_),
    .X(net80));
 sky130_fd_sc_hd__mux2_1 _017_ (.A0(net41),
    .A1(net9),
    .S(_003_),
    .X(net81));
 sky130_fd_sc_hd__mux2_1 _018_ (.A0(net42),
    .A1(net10),
    .S(_003_),
    .X(net82));
 sky130_fd_sc_hd__mux2_1 _019_ (.A0(net43),
    .A1(net11),
    .S(_003_),
    .X(net83));
 sky130_fd_sc_hd__mux2_1 _020_ (.A0(net44),
    .A1(net12),
    .S(_003_),
    .X(net84));
 sky130_fd_sc_hd__mux2_1 _021_ (.A0(net45),
    .A1(net13),
    .S(_003_),
    .X(net85));
 sky130_fd_sc_hd__mux2_1 _022_ (.A0(net46),
    .A1(net14),
    .S(_003_),
    .X(net86));
 sky130_fd_sc_hd__buf_6 _023_ (.A(_002_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _024_ (.A0(net47),
    .A1(net15),
    .S(_004_),
    .X(net87));
 sky130_fd_sc_hd__mux2_1 _025_ (.A0(net48),
    .A1(net16),
    .S(_004_),
    .X(net88));
 sky130_fd_sc_hd__mux2_1 _026_ (.A0(net49),
    .A1(net17),
    .S(_004_),
    .X(net89));
 sky130_fd_sc_hd__mux2_1 _027_ (.A0(net50),
    .A1(net18),
    .S(_004_),
    .X(net90));
 sky130_fd_sc_hd__mux2_1 _028_ (.A0(net51),
    .A1(net19),
    .S(_004_),
    .X(net91));
 sky130_fd_sc_hd__mux2_1 _029_ (.A0(net52),
    .A1(net20),
    .S(_004_),
    .X(net92));
 sky130_fd_sc_hd__mux2_1 _030_ (.A0(net53),
    .A1(net21),
    .S(_004_),
    .X(net93));
 sky130_fd_sc_hd__mux2_1 _031_ (.A0(net54),
    .A1(net22),
    .S(_004_),
    .X(net94));
 sky130_fd_sc_hd__mux2_1 _032_ (.A0(net55),
    .A1(net23),
    .S(_004_),
    .X(net95));
 sky130_fd_sc_hd__mux2_1 _033_ (.A0(net56),
    .A1(net24),
    .S(_004_),
    .X(net96));
 sky130_fd_sc_hd__buf_6 _034_ (.A(_002_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _035_ (.A0(net57),
    .A1(net25),
    .S(_005_),
    .X(net97));
 sky130_fd_sc_hd__mux2_1 _036_ (.A0(net58),
    .A1(net26),
    .S(_005_),
    .X(net98));
 sky130_fd_sc_hd__mux2_1 _037_ (.A0(net59),
    .A1(net27),
    .S(_005_),
    .X(net99));
 sky130_fd_sc_hd__mux2_1 _038_ (.A0(net60),
    .A1(net28),
    .S(_005_),
    .X(net100));
 sky130_fd_sc_hd__mux2_1 _039_ (.A0(net61),
    .A1(net29),
    .S(_005_),
    .X(net101));
 sky130_fd_sc_hd__mux2_1 _040_ (.A0(net62),
    .A1(net30),
    .S(_005_),
    .X(net102));
 sky130_fd_sc_hd__mux2_1 _041_ (.A0(net63),
    .A1(net31),
    .S(_005_),
    .X(net103));
 sky130_fd_sc_hd__mux2_1 _042_ (.A0(net64),
    .A1(net32),
    .S(_005_),
    .X(net104));
 sky130_fd_sc_hd__mux2_1 _043_ (.A0(net65),
    .A1(net33),
    .S(_005_),
    .X(net105));
 sky130_fd_sc_hd__mux2_1 _044_ (.A0(net66),
    .A1(net34),
    .S(_005_),
    .X(net106));
 sky130_fd_sc_hd__mux2_1 _045_ (.A0(net67),
    .A1(net35),
    .S(_002_),
    .X(net107));
 sky130_fd_sc_hd__mux2_1 _046_ (.A0(net68),
    .A1(net36),
    .S(_002_),
    .X(net108));
 sky130_fd_sc_hd__mux2_1 _047_ (.A0(net69),
    .A1(net37),
    .S(_002_),
    .X(net109));
 sky130_fd_sc_hd__or2_0 _048_ (.A(_003_),
    .B(net70),
    .X(net110));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__conb_1 _086__179 (.HI(net179));
 sky130_fd_sc_hd__buf_4 _051_ (.A(net111),
    .X(instr_done_wb_o));
 sky130_fd_sc_hd__buf_4 _052_ (.A(net112),
    .X(outstanding_load_wb_o));
 sky130_fd_sc_hd__buf_4 _053_ (.A(net113),
    .X(outstanding_store_wb_o));
 sky130_fd_sc_hd__buf_4 _054_ (.A(net114),
    .X(pc_wb_o[0]));
 sky130_fd_sc_hd__buf_4 _055_ (.A(net115),
    .X(pc_wb_o[1]));
 sky130_fd_sc_hd__buf_4 _056_ (.A(net116),
    .X(pc_wb_o[2]));
 sky130_fd_sc_hd__buf_4 _057_ (.A(net117),
    .X(pc_wb_o[3]));
 sky130_fd_sc_hd__buf_4 _058_ (.A(net118),
    .X(pc_wb_o[4]));
 sky130_fd_sc_hd__buf_4 _059_ (.A(net119),
    .X(pc_wb_o[5]));
 sky130_fd_sc_hd__buf_4 _060_ (.A(net120),
    .X(pc_wb_o[6]));
 sky130_fd_sc_hd__buf_4 _061_ (.A(net121),
    .X(pc_wb_o[7]));
 sky130_fd_sc_hd__buf_4 _062_ (.A(net122),
    .X(pc_wb_o[8]));
 sky130_fd_sc_hd__buf_4 _063_ (.A(net123),
    .X(pc_wb_o[9]));
 sky130_fd_sc_hd__buf_4 _064_ (.A(net124),
    .X(pc_wb_o[10]));
 sky130_fd_sc_hd__buf_4 _065_ (.A(net125),
    .X(pc_wb_o[11]));
 sky130_fd_sc_hd__buf_4 _066_ (.A(net126),
    .X(pc_wb_o[12]));
 sky130_fd_sc_hd__buf_4 _067_ (.A(net127),
    .X(pc_wb_o[13]));
 sky130_fd_sc_hd__buf_4 _068_ (.A(net128),
    .X(pc_wb_o[14]));
 sky130_fd_sc_hd__buf_4 _069_ (.A(net129),
    .X(pc_wb_o[15]));
 sky130_fd_sc_hd__buf_4 _070_ (.A(net130),
    .X(pc_wb_o[16]));
 sky130_fd_sc_hd__buf_4 _071_ (.A(net131),
    .X(pc_wb_o[17]));
 sky130_fd_sc_hd__buf_4 _072_ (.A(net132),
    .X(pc_wb_o[18]));
 sky130_fd_sc_hd__buf_4 _073_ (.A(net133),
    .X(pc_wb_o[19]));
 sky130_fd_sc_hd__buf_4 _074_ (.A(net134),
    .X(pc_wb_o[20]));
 sky130_fd_sc_hd__buf_4 _075_ (.A(net135),
    .X(pc_wb_o[21]));
 sky130_fd_sc_hd__buf_4 _076_ (.A(net136),
    .X(pc_wb_o[22]));
 sky130_fd_sc_hd__buf_4 _077_ (.A(net137),
    .X(pc_wb_o[23]));
 sky130_fd_sc_hd__buf_4 _078_ (.A(net138),
    .X(pc_wb_o[24]));
 sky130_fd_sc_hd__buf_4 _079_ (.A(net139),
    .X(pc_wb_o[25]));
 sky130_fd_sc_hd__buf_4 _080_ (.A(net140),
    .X(pc_wb_o[26]));
 sky130_fd_sc_hd__buf_4 _081_ (.A(net141),
    .X(pc_wb_o[27]));
 sky130_fd_sc_hd__buf_4 _082_ (.A(net142),
    .X(pc_wb_o[28]));
 sky130_fd_sc_hd__buf_4 _083_ (.A(net143),
    .X(pc_wb_o[29]));
 sky130_fd_sc_hd__buf_4 _084_ (.A(net144),
    .X(pc_wb_o[30]));
 sky130_fd_sc_hd__buf_4 _085_ (.A(net145),
    .X(pc_wb_o[31]));
 sky130_fd_sc_hd__buf_4 _086_ (.A(net179),
    .X(ready_wb_o));
 sky130_fd_sc_hd__clkbuf_1 _087_ (.A(rf_waddr_id_i[0]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(rf_waddr_id_i[1]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(rf_waddr_id_i[2]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(rf_waddr_id_i[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(rf_waddr_id_i[4]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 _092_ (.A(net146),
    .X(rf_wdata_fwd_wb_o[0]));
 sky130_fd_sc_hd__buf_4 _093_ (.A(net147),
    .X(rf_wdata_fwd_wb_o[1]));
 sky130_fd_sc_hd__buf_4 _094_ (.A(net148),
    .X(rf_wdata_fwd_wb_o[2]));
 sky130_fd_sc_hd__buf_4 _095_ (.A(net149),
    .X(rf_wdata_fwd_wb_o[3]));
 sky130_fd_sc_hd__buf_4 _096_ (.A(net150),
    .X(rf_wdata_fwd_wb_o[4]));
 sky130_fd_sc_hd__buf_4 _097_ (.A(net151),
    .X(rf_wdata_fwd_wb_o[5]));
 sky130_fd_sc_hd__buf_4 _098_ (.A(net152),
    .X(rf_wdata_fwd_wb_o[6]));
 sky130_fd_sc_hd__buf_4 _099_ (.A(net153),
    .X(rf_wdata_fwd_wb_o[7]));
 sky130_fd_sc_hd__buf_4 _100_ (.A(net154),
    .X(rf_wdata_fwd_wb_o[8]));
 sky130_fd_sc_hd__buf_4 _101_ (.A(net155),
    .X(rf_wdata_fwd_wb_o[9]));
 sky130_fd_sc_hd__buf_4 _102_ (.A(net156),
    .X(rf_wdata_fwd_wb_o[10]));
 sky130_fd_sc_hd__buf_4 _103_ (.A(net157),
    .X(rf_wdata_fwd_wb_o[11]));
 sky130_fd_sc_hd__buf_4 _104_ (.A(net158),
    .X(rf_wdata_fwd_wb_o[12]));
 sky130_fd_sc_hd__buf_4 _105_ (.A(net159),
    .X(rf_wdata_fwd_wb_o[13]));
 sky130_fd_sc_hd__buf_4 _106_ (.A(net160),
    .X(rf_wdata_fwd_wb_o[14]));
 sky130_fd_sc_hd__buf_4 _107_ (.A(net161),
    .X(rf_wdata_fwd_wb_o[15]));
 sky130_fd_sc_hd__buf_4 _108_ (.A(net162),
    .X(rf_wdata_fwd_wb_o[16]));
 sky130_fd_sc_hd__buf_4 _109_ (.A(net163),
    .X(rf_wdata_fwd_wb_o[17]));
 sky130_fd_sc_hd__buf_4 _110_ (.A(net164),
    .X(rf_wdata_fwd_wb_o[18]));
 sky130_fd_sc_hd__buf_4 _111_ (.A(net165),
    .X(rf_wdata_fwd_wb_o[19]));
 sky130_fd_sc_hd__buf_4 _112_ (.A(net166),
    .X(rf_wdata_fwd_wb_o[20]));
 sky130_fd_sc_hd__buf_4 _113_ (.A(net167),
    .X(rf_wdata_fwd_wb_o[21]));
 sky130_fd_sc_hd__buf_4 _114_ (.A(net168),
    .X(rf_wdata_fwd_wb_o[22]));
 sky130_fd_sc_hd__buf_4 _115_ (.A(net169),
    .X(rf_wdata_fwd_wb_o[23]));
 sky130_fd_sc_hd__buf_4 _116_ (.A(net170),
    .X(rf_wdata_fwd_wb_o[24]));
 sky130_fd_sc_hd__buf_4 _117_ (.A(net171),
    .X(rf_wdata_fwd_wb_o[25]));
 sky130_fd_sc_hd__buf_4 _118_ (.A(net172),
    .X(rf_wdata_fwd_wb_o[26]));
 sky130_fd_sc_hd__buf_4 _119_ (.A(net173),
    .X(rf_wdata_fwd_wb_o[27]));
 sky130_fd_sc_hd__buf_4 _120_ (.A(net174),
    .X(rf_wdata_fwd_wb_o[28]));
 sky130_fd_sc_hd__buf_4 _121_ (.A(net175),
    .X(rf_wdata_fwd_wb_o[29]));
 sky130_fd_sc_hd__buf_4 _122_ (.A(net176),
    .X(rf_wdata_fwd_wb_o[30]));
 sky130_fd_sc_hd__buf_4 _123_ (.A(net177),
    .X(rf_wdata_fwd_wb_o[31]));
 sky130_fd_sc_hd__buf_4 _124_ (.A(net178),
    .X(rf_write_wb_o));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_93 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(en_wb_i),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(instr_is_compressed_id_i),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(instr_perf_count_id_i),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(lsu_resp_err_i),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(lsu_resp_valid_i),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(rf_wdata_id_i[0]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(rf_wdata_id_i[10]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(rf_wdata_id_i[11]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(rf_wdata_id_i[12]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(rf_wdata_id_i[13]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(rf_wdata_id_i[14]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(rf_wdata_id_i[15]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(rf_wdata_id_i[16]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(rf_wdata_id_i[17]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(rf_wdata_id_i[18]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(rf_wdata_id_i[19]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(rf_wdata_id_i[1]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(rf_wdata_id_i[20]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(rf_wdata_id_i[21]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(rf_wdata_id_i[22]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(rf_wdata_id_i[23]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(rf_wdata_id_i[24]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(rf_wdata_id_i[25]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(rf_wdata_id_i[26]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(rf_wdata_id_i[27]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(rf_wdata_id_i[28]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(rf_wdata_id_i[29]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(rf_wdata_id_i[2]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(rf_wdata_id_i[30]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(rf_wdata_id_i[31]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(rf_wdata_id_i[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(rf_wdata_id_i[4]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(rf_wdata_id_i[5]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(rf_wdata_id_i[6]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(rf_wdata_id_i[7]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(rf_wdata_id_i[8]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(rf_wdata_id_i[9]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(rf_wdata_lsu_i[0]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(rf_wdata_lsu_i[10]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(rf_wdata_lsu_i[11]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(rf_wdata_lsu_i[12]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(rf_wdata_lsu_i[13]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(rf_wdata_lsu_i[14]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(rf_wdata_lsu_i[15]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(rf_wdata_lsu_i[16]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(rf_wdata_lsu_i[17]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(rf_wdata_lsu_i[18]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(rf_wdata_lsu_i[19]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(rf_wdata_lsu_i[1]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(rf_wdata_lsu_i[20]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(rf_wdata_lsu_i[21]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(rf_wdata_lsu_i[22]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(rf_wdata_lsu_i[23]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(rf_wdata_lsu_i[24]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(rf_wdata_lsu_i[25]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(rf_wdata_lsu_i[26]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(rf_wdata_lsu_i[27]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(rf_wdata_lsu_i[28]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(rf_wdata_lsu_i[29]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(rf_wdata_lsu_i[2]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(rf_wdata_lsu_i[30]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(rf_wdata_lsu_i[31]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(rf_wdata_lsu_i[3]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(rf_wdata_lsu_i[4]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(rf_wdata_lsu_i[5]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(rf_wdata_lsu_i[6]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(rf_wdata_lsu_i[7]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(rf_wdata_lsu_i[8]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(rf_wdata_lsu_i[9]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(rf_we_lsu_i),
    .X(net70));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(perf_instr_ret_compressed_wb_o));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(perf_instr_ret_wb_o));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(rf_waddr_wb_o[0]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(rf_waddr_wb_o[1]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(rf_waddr_wb_o[2]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(rf_waddr_wb_o[3]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(rf_waddr_wb_o[4]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(rf_wdata_wb_o[0]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(rf_wdata_wb_o[10]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(rf_wdata_wb_o[11]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(rf_wdata_wb_o[12]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(rf_wdata_wb_o[13]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(rf_wdata_wb_o[14]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(rf_wdata_wb_o[15]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(rf_wdata_wb_o[16]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(rf_wdata_wb_o[17]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(rf_wdata_wb_o[18]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(rf_wdata_wb_o[19]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(rf_wdata_wb_o[1]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(rf_wdata_wb_o[20]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(rf_wdata_wb_o[21]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(rf_wdata_wb_o[22]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(rf_wdata_wb_o[23]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(rf_wdata_wb_o[24]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(rf_wdata_wb_o[25]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(rf_wdata_wb_o[26]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(rf_wdata_wb_o[27]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(rf_wdata_wb_o[28]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(rf_wdata_wb_o[29]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(rf_wdata_wb_o[2]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(rf_wdata_wb_o[30]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(rf_wdata_wb_o[31]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(rf_wdata_wb_o[3]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(rf_wdata_wb_o[4]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(rf_wdata_wb_o[5]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(rf_wdata_wb_o[6]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(rf_wdata_wb_o[7]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(rf_wdata_wb_o[8]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(rf_wdata_wb_o[9]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(rf_we_wb_o));
 sky130_fd_sc_hd__conb_1 _051__111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 _052__112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 _053__113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 _054__114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 _055__115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 _056__116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 _057__117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 _058__118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 _059__119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 _060__120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 _061__121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 _062__122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 _063__123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 _064__124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 _065__125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 _066__126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 _067__127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 _068__128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 _069__129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 _070__130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 _071__131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 _072__132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 _073__133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 _074__134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 _075__135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 _076__136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 _077__137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 _078__138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 _079__139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 _080__140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 _081__141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 _082__142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 _083__143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 _084__144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 _085__145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 _092__146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 _093__147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 _094__148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 _095__149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 _096__150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 _097__151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 _098__152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 _099__153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 _100__154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 _101__155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 _102__156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 _103__157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 _104__158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 _105__159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 _106__160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 _107__161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 _108__162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 _109__163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 _110__164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 _111__165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 _112__166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 _113__167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 _114__168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 _115__169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 _116__170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 _117__171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 _118__172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 _119__173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 _120__174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 _121__175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 _122__176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 _123__177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 _124__178 (.LO(net178));
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_119 ();
endmodule
