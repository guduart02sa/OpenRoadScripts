VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA fakeram7_256x32_via1_2_3132_18_1_87_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 87 ;
END fakeram7_256x32_via1_2_3132_18_1_87_36_36

VIA fakeram7_256x32_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END fakeram7_256x32_VIA23_1_3_36_36

VIA fakeram7_256x32_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END fakeram7_256x32_VIA34_1_2_58_52

VIA fakeram7_256x32_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END fakeram7_256x32_VIA45_1_2_58_58

VIA fakeram7_256x32_VIA45_2_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.06 0.052 0.06 ;
    LAYER M5 ;
      RECT  -0.06 -0.052 0.06 0.052 ;
    LAYER V4 ;
      RECT  0.017 0.017 0.041 0.041 ;
      RECT  -0.041 0.017 -0.017 0.041 ;
      RECT  0.017 -0.041 0.041 -0.017 ;
      RECT  -0.041 -0.041 -0.017 -0.017 ;
END fakeram7_256x32_VIA45_2_2_58_58

MACRO fakeram7_256x32
  FOREIGN fakeram7_256x32 0 0 ;
  CLASS BLOCK ;
  SIZE 5.163 BY 27.304 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M5 ;
        RECT  2.658 0.684 2.778 26.586 ;
      LAYER M2 ;
        RECT  1.026 26.181 4.158 26.199 ;
        RECT  1.026 25.641 4.158 25.659 ;
        RECT  1.026 25.101 4.158 25.119 ;
        RECT  1.026 24.561 4.158 24.579 ;
        RECT  1.026 24.021 4.158 24.039 ;
        RECT  1.026 23.481 4.158 23.499 ;
        RECT  1.026 22.941 4.158 22.959 ;
        RECT  1.026 22.401 4.158 22.419 ;
        RECT  1.026 21.861 4.158 21.879 ;
        RECT  1.026 21.321 4.158 21.339 ;
        RECT  1.026 20.781 4.158 20.799 ;
        RECT  1.026 20.241 4.158 20.259 ;
        RECT  1.026 19.701 4.158 19.719 ;
        RECT  1.026 19.161 4.158 19.179 ;
        RECT  1.026 18.621 4.158 18.639 ;
        RECT  1.026 18.081 4.158 18.099 ;
        RECT  1.026 17.541 4.158 17.559 ;
        RECT  1.026 17.001 4.158 17.019 ;
        RECT  1.026 16.461 4.158 16.479 ;
        RECT  1.026 15.921 4.158 15.939 ;
        RECT  1.026 15.381 4.158 15.399 ;
        RECT  1.026 14.841 4.158 14.859 ;
        RECT  1.026 14.301 4.158 14.319 ;
        RECT  1.026 13.761 4.158 13.779 ;
        RECT  1.026 13.221 4.158 13.239 ;
        RECT  1.026 12.681 4.158 12.699 ;
        RECT  1.026 12.141 4.158 12.159 ;
        RECT  1.026 11.601 4.158 11.619 ;
        RECT  1.026 11.061 4.158 11.079 ;
        RECT  1.026 10.521 4.158 10.539 ;
        RECT  1.026 9.981 4.158 9.999 ;
        RECT  1.026 9.441 4.158 9.459 ;
        RECT  1.026 8.901 4.158 8.919 ;
        RECT  1.026 8.361 4.158 8.379 ;
        RECT  1.026 7.821 4.158 7.839 ;
        RECT  1.026 7.281 4.158 7.299 ;
        RECT  1.026 6.741 4.158 6.759 ;
        RECT  1.026 6.201 4.158 6.219 ;
        RECT  1.026 5.661 4.158 5.679 ;
        RECT  1.026 5.121 4.158 5.139 ;
        RECT  1.026 4.581 4.158 4.599 ;
        RECT  1.026 4.041 4.158 4.059 ;
        RECT  1.026 3.501 4.158 3.519 ;
        RECT  1.026 2.961 4.158 2.979 ;
        RECT  1.026 2.421 4.158 2.439 ;
        RECT  1.026 1.881 4.158 1.899 ;
        RECT  1.026 1.341 4.158 1.359 ;
      LAYER M1 ;
        RECT  1.026 26.181 4.158 26.199 ;
        RECT  1.026 25.641 4.158 25.659 ;
        RECT  1.026 25.101 4.158 25.119 ;
        RECT  1.026 24.561 4.158 24.579 ;
        RECT  1.026 24.021 4.158 24.039 ;
        RECT  1.026 23.481 4.158 23.499 ;
        RECT  1.026 22.941 4.158 22.959 ;
        RECT  1.026 22.401 4.158 22.419 ;
        RECT  1.026 21.861 4.158 21.879 ;
        RECT  1.026 21.321 4.158 21.339 ;
        RECT  1.026 20.781 4.158 20.799 ;
        RECT  1.026 20.241 4.158 20.259 ;
        RECT  1.026 19.701 4.158 19.719 ;
        RECT  1.026 19.161 4.158 19.179 ;
        RECT  1.026 18.621 4.158 18.639 ;
        RECT  1.026 18.081 4.158 18.099 ;
        RECT  1.026 17.541 4.158 17.559 ;
        RECT  1.026 17.001 4.158 17.019 ;
        RECT  1.026 16.461 4.158 16.479 ;
        RECT  1.026 15.921 4.158 15.939 ;
        RECT  1.026 15.381 4.158 15.399 ;
        RECT  1.026 14.841 4.158 14.859 ;
        RECT  1.026 14.301 4.158 14.319 ;
        RECT  1.026 13.761 4.158 13.779 ;
        RECT  1.026 13.221 4.158 13.239 ;
        RECT  1.026 12.681 4.158 12.699 ;
        RECT  1.026 12.141 4.158 12.159 ;
        RECT  1.026 11.601 4.158 11.619 ;
        RECT  1.026 11.061 4.158 11.079 ;
        RECT  1.026 10.521 4.158 10.539 ;
        RECT  1.026 9.981 4.158 9.999 ;
        RECT  1.026 9.441 4.158 9.459 ;
        RECT  1.026 8.901 4.158 8.919 ;
        RECT  1.026 8.361 4.158 8.379 ;
        RECT  1.026 7.821 4.158 7.839 ;
        RECT  1.026 7.281 4.158 7.299 ;
        RECT  1.026 6.741 4.158 6.759 ;
        RECT  1.026 6.201 4.158 6.219 ;
        RECT  1.026 5.661 4.158 5.679 ;
        RECT  1.026 5.121 4.158 5.139 ;
        RECT  1.026 4.581 4.158 4.599 ;
        RECT  1.026 4.041 4.158 4.059 ;
        RECT  1.026 3.501 4.158 3.519 ;
        RECT  1.026 2.961 4.158 2.979 ;
        RECT  1.026 2.421 4.158 2.439 ;
        RECT  1.026 1.881 4.158 1.899 ;
        RECT  1.026 1.341 4.158 1.359 ;
      LAYER M5 ;
        RECT  4.434 0.684 4.554 26.586 ;
      LAYER M4 ;
        RECT  0.63 26.466 4.554 26.586 ;
        RECT  0.63 0.684 4.554 0.804 ;
      LAYER M5 ;
        RECT  0.63 0.684 0.75 26.586 ;
      VIA 4.494 26.526 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 4.494 0.744 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 2.718 26.526 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 2.718 0.744 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 0.69 26.526 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 0.69 0.744 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 2.718 26.19 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 26.173 2.763 26.207 ;
      VIA 2.718 26.19 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 26.19 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 25.65 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 25.633 2.763 25.667 ;
      VIA 2.718 25.65 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 25.65 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 25.11 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 25.093 2.763 25.127 ;
      VIA 2.718 25.11 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 25.11 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 24.57 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 24.553 2.763 24.587 ;
      VIA 2.718 24.57 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 24.57 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 24.03 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 24.013 2.763 24.047 ;
      VIA 2.718 24.03 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 24.03 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 23.49 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 23.473 2.763 23.507 ;
      VIA 2.718 23.49 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 23.49 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 22.95 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 22.933 2.763 22.967 ;
      VIA 2.718 22.95 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 22.95 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 22.41 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 22.393 2.763 22.427 ;
      VIA 2.718 22.41 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 22.41 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 21.87 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 21.853 2.763 21.887 ;
      VIA 2.718 21.87 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 21.87 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 21.33 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 21.313 2.763 21.347 ;
      VIA 2.718 21.33 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 21.33 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 20.79 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 20.773 2.763 20.807 ;
      VIA 2.718 20.79 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 20.79 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 20.25 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 20.233 2.763 20.267 ;
      VIA 2.718 20.25 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 20.25 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 19.71 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 19.693 2.763 19.727 ;
      VIA 2.718 19.71 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 19.71 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 19.17 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 19.153 2.763 19.187 ;
      VIA 2.718 19.17 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 19.17 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 18.63 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 18.613 2.763 18.647 ;
      VIA 2.718 18.63 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 18.63 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 18.09 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 18.073 2.763 18.107 ;
      VIA 2.718 18.09 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 18.09 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 17.55 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 17.533 2.763 17.567 ;
      VIA 2.718 17.55 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 17.55 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 17.01 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 16.993 2.763 17.027 ;
      VIA 2.718 17.01 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 17.01 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 16.47 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 16.453 2.763 16.487 ;
      VIA 2.718 16.47 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 16.47 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 15.93 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 15.913 2.763 15.947 ;
      VIA 2.718 15.93 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 15.93 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 15.39 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 15.373 2.763 15.407 ;
      VIA 2.718 15.39 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 15.39 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 14.85 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 14.833 2.763 14.867 ;
      VIA 2.718 14.85 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 14.85 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 14.31 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 14.293 2.763 14.327 ;
      VIA 2.718 14.31 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 14.31 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 13.77 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 13.753 2.763 13.787 ;
      VIA 2.718 13.77 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 13.77 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 13.23 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 13.213 2.763 13.247 ;
      VIA 2.718 13.23 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 13.23 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 12.69 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 12.673 2.763 12.707 ;
      VIA 2.718 12.69 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 12.69 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 12.15 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 12.133 2.763 12.167 ;
      VIA 2.718 12.15 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 12.15 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 11.61 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 11.593 2.763 11.627 ;
      VIA 2.718 11.61 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 11.61 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 11.07 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 11.053 2.763 11.087 ;
      VIA 2.718 11.07 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 11.07 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 10.53 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 10.513 2.763 10.547 ;
      VIA 2.718 10.53 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 10.53 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 9.99 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 9.973 2.763 10.007 ;
      VIA 2.718 9.99 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 9.99 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 9.45 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 9.433 2.763 9.467 ;
      VIA 2.718 9.45 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 9.45 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 8.91 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 8.893 2.763 8.927 ;
      VIA 2.718 8.91 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 8.91 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 8.37 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 8.353 2.763 8.387 ;
      VIA 2.718 8.37 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 8.37 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 7.83 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 7.813 2.763 7.847 ;
      VIA 2.718 7.83 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 7.83 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 7.29 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 7.273 2.763 7.307 ;
      VIA 2.718 7.29 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 7.29 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 6.75 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 6.733 2.763 6.767 ;
      VIA 2.718 6.75 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 6.75 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 6.21 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 6.193 2.763 6.227 ;
      VIA 2.718 6.21 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 6.21 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 5.67 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 5.653 2.763 5.687 ;
      VIA 2.718 5.67 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 5.67 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 5.13 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 5.113 2.763 5.147 ;
      VIA 2.718 5.13 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 5.13 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 4.59 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 4.573 2.763 4.607 ;
      VIA 2.718 4.59 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 4.59 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 4.05 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 4.033 2.763 4.067 ;
      VIA 2.718 4.05 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 4.05 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 3.51 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 3.493 2.763 3.527 ;
      VIA 2.718 3.51 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 3.51 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 2.97 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 2.953 2.763 2.987 ;
      VIA 2.718 2.97 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 2.97 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 2.43 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 2.413 2.763 2.447 ;
      VIA 2.718 2.43 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 2.43 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 1.89 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 1.873 2.763 1.907 ;
      VIA 2.718 1.89 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 1.89 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.718 1.35 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.673 1.333 2.763 1.367 ;
      VIA 2.718 1.35 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.718 1.35 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.592 26.19 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 25.65 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 25.11 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 24.57 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 24.03 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 23.49 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 22.95 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 22.41 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 21.87 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 21.33 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 20.79 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 20.25 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 19.71 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 19.17 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 18.63 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 18.09 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 17.55 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 17.01 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 16.47 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 15.93 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 15.39 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 14.85 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 14.31 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 13.77 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 13.23 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 12.69 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 12.15 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 11.61 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 11.07 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 10.53 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 9.99 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 9.45 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 8.91 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 8.37 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 7.83 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 7.29 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 6.75 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 6.21 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 5.67 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 5.13 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 4.59 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 4.05 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 3.51 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 2.97 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 2.43 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 1.89 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 1.35 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M5 ;
        RECT  2.466 0.876 2.586 26.394 ;
      LAYER M2 ;
        RECT  1.026 25.911 4.158 25.929 ;
        RECT  1.026 25.371 4.158 25.389 ;
        RECT  1.026 24.831 4.158 24.849 ;
        RECT  1.026 24.291 4.158 24.309 ;
        RECT  1.026 23.751 4.158 23.769 ;
        RECT  1.026 23.211 4.158 23.229 ;
        RECT  1.026 22.671 4.158 22.689 ;
        RECT  1.026 22.131 4.158 22.149 ;
        RECT  1.026 21.591 4.158 21.609 ;
        RECT  1.026 21.051 4.158 21.069 ;
        RECT  1.026 20.511 4.158 20.529 ;
        RECT  1.026 19.971 4.158 19.989 ;
        RECT  1.026 19.431 4.158 19.449 ;
        RECT  1.026 18.891 4.158 18.909 ;
        RECT  1.026 18.351 4.158 18.369 ;
        RECT  1.026 17.811 4.158 17.829 ;
        RECT  1.026 17.271 4.158 17.289 ;
        RECT  1.026 16.731 4.158 16.749 ;
        RECT  1.026 16.191 4.158 16.209 ;
        RECT  1.026 15.651 4.158 15.669 ;
        RECT  1.026 15.111 4.158 15.129 ;
        RECT  1.026 14.571 4.158 14.589 ;
        RECT  1.026 14.031 4.158 14.049 ;
        RECT  1.026 13.491 4.158 13.509 ;
        RECT  1.026 12.951 4.158 12.969 ;
        RECT  1.026 12.411 4.158 12.429 ;
        RECT  1.026 11.871 4.158 11.889 ;
        RECT  1.026 11.331 4.158 11.349 ;
        RECT  1.026 10.791 4.158 10.809 ;
        RECT  1.026 10.251 4.158 10.269 ;
        RECT  1.026 9.711 4.158 9.729 ;
        RECT  1.026 9.171 4.158 9.189 ;
        RECT  1.026 8.631 4.158 8.649 ;
        RECT  1.026 8.091 4.158 8.109 ;
        RECT  1.026 7.551 4.158 7.569 ;
        RECT  1.026 7.011 4.158 7.029 ;
        RECT  1.026 6.471 4.158 6.489 ;
        RECT  1.026 5.931 4.158 5.949 ;
        RECT  1.026 5.391 4.158 5.409 ;
        RECT  1.026 4.851 4.158 4.869 ;
        RECT  1.026 4.311 4.158 4.329 ;
        RECT  1.026 3.771 4.158 3.789 ;
        RECT  1.026 3.231 4.158 3.249 ;
        RECT  1.026 2.691 4.158 2.709 ;
        RECT  1.026 2.151 4.158 2.169 ;
        RECT  1.026 1.611 4.158 1.629 ;
        RECT  1.026 1.071 4.158 1.089 ;
      LAYER M1 ;
        RECT  1.026 25.911 4.158 25.929 ;
        RECT  1.026 25.371 4.158 25.389 ;
        RECT  1.026 24.831 4.158 24.849 ;
        RECT  1.026 24.291 4.158 24.309 ;
        RECT  1.026 23.751 4.158 23.769 ;
        RECT  1.026 23.211 4.158 23.229 ;
        RECT  1.026 22.671 4.158 22.689 ;
        RECT  1.026 22.131 4.158 22.149 ;
        RECT  1.026 21.591 4.158 21.609 ;
        RECT  1.026 21.051 4.158 21.069 ;
        RECT  1.026 20.511 4.158 20.529 ;
        RECT  1.026 19.971 4.158 19.989 ;
        RECT  1.026 19.431 4.158 19.449 ;
        RECT  1.026 18.891 4.158 18.909 ;
        RECT  1.026 18.351 4.158 18.369 ;
        RECT  1.026 17.811 4.158 17.829 ;
        RECT  1.026 17.271 4.158 17.289 ;
        RECT  1.026 16.731 4.158 16.749 ;
        RECT  1.026 16.191 4.158 16.209 ;
        RECT  1.026 15.651 4.158 15.669 ;
        RECT  1.026 15.111 4.158 15.129 ;
        RECT  1.026 14.571 4.158 14.589 ;
        RECT  1.026 14.031 4.158 14.049 ;
        RECT  1.026 13.491 4.158 13.509 ;
        RECT  1.026 12.951 4.158 12.969 ;
        RECT  1.026 12.411 4.158 12.429 ;
        RECT  1.026 11.871 4.158 11.889 ;
        RECT  1.026 11.331 4.158 11.349 ;
        RECT  1.026 10.791 4.158 10.809 ;
        RECT  1.026 10.251 4.158 10.269 ;
        RECT  1.026 9.711 4.158 9.729 ;
        RECT  1.026 9.171 4.158 9.189 ;
        RECT  1.026 8.631 4.158 8.649 ;
        RECT  1.026 8.091 4.158 8.109 ;
        RECT  1.026 7.551 4.158 7.569 ;
        RECT  1.026 7.011 4.158 7.029 ;
        RECT  1.026 6.471 4.158 6.489 ;
        RECT  1.026 5.931 4.158 5.949 ;
        RECT  1.026 5.391 4.158 5.409 ;
        RECT  1.026 4.851 4.158 4.869 ;
        RECT  1.026 4.311 4.158 4.329 ;
        RECT  1.026 3.771 4.158 3.789 ;
        RECT  1.026 3.231 4.158 3.249 ;
        RECT  1.026 2.691 4.158 2.709 ;
        RECT  1.026 2.151 4.158 2.169 ;
        RECT  1.026 1.611 4.158 1.629 ;
        RECT  1.026 1.071 4.158 1.089 ;
      LAYER M5 ;
        RECT  4.242 0.876 4.362 26.394 ;
      LAYER M4 ;
        RECT  0.822 26.274 4.362 26.394 ;
        RECT  0.822 0.876 4.362 0.996 ;
      LAYER M5 ;
        RECT  0.822 0.876 0.942 26.394 ;
      VIA 4.302 26.334 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 4.302 0.936 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 2.526 26.334 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 2.526 0.936 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 0.882 26.334 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 0.882 0.936 fakeram7_256x32_VIA45_2_2_58_58 ;
      VIA 2.526 25.92 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 25.903 2.571 25.937 ;
      VIA 2.526 25.92 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 25.92 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 25.38 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 25.363 2.571 25.397 ;
      VIA 2.526 25.38 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 25.38 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 24.84 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 24.823 2.571 24.857 ;
      VIA 2.526 24.84 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 24.84 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 24.3 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 24.283 2.571 24.317 ;
      VIA 2.526 24.3 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 24.3 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 23.76 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 23.743 2.571 23.777 ;
      VIA 2.526 23.76 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 23.76 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 23.22 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 23.203 2.571 23.237 ;
      VIA 2.526 23.22 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 23.22 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 22.68 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 22.663 2.571 22.697 ;
      VIA 2.526 22.68 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 22.68 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 22.14 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 22.123 2.571 22.157 ;
      VIA 2.526 22.14 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 22.14 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 21.6 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 21.583 2.571 21.617 ;
      VIA 2.526 21.6 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 21.6 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 21.06 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 21.043 2.571 21.077 ;
      VIA 2.526 21.06 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 21.06 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 20.52 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 20.503 2.571 20.537 ;
      VIA 2.526 20.52 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 20.52 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 19.98 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 19.963 2.571 19.997 ;
      VIA 2.526 19.98 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 19.98 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 19.44 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 19.423 2.571 19.457 ;
      VIA 2.526 19.44 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 19.44 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 18.9 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 18.883 2.571 18.917 ;
      VIA 2.526 18.9 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 18.9 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 18.36 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 18.343 2.571 18.377 ;
      VIA 2.526 18.36 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 18.36 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 17.82 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 17.803 2.571 17.837 ;
      VIA 2.526 17.82 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 17.82 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 17.28 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 17.263 2.571 17.297 ;
      VIA 2.526 17.28 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 17.28 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 16.74 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 16.723 2.571 16.757 ;
      VIA 2.526 16.74 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 16.74 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 16.2 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 16.183 2.571 16.217 ;
      VIA 2.526 16.2 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 16.2 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 15.66 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 15.643 2.571 15.677 ;
      VIA 2.526 15.66 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 15.66 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 15.12 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 15.103 2.571 15.137 ;
      VIA 2.526 15.12 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 15.12 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 14.58 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 14.563 2.571 14.597 ;
      VIA 2.526 14.58 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 14.58 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 14.04 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 14.023 2.571 14.057 ;
      VIA 2.526 14.04 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 14.04 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 13.5 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 13.483 2.571 13.517 ;
      VIA 2.526 13.5 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 13.5 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 12.96 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 12.943 2.571 12.977 ;
      VIA 2.526 12.96 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 12.96 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 12.42 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 12.403 2.571 12.437 ;
      VIA 2.526 12.42 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 12.42 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 11.88 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 11.863 2.571 11.897 ;
      VIA 2.526 11.88 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 11.88 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 11.34 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 11.323 2.571 11.357 ;
      VIA 2.526 11.34 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 11.34 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 10.8 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 10.783 2.571 10.817 ;
      VIA 2.526 10.8 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 10.8 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 10.26 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 10.243 2.571 10.277 ;
      VIA 2.526 10.26 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 10.26 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 9.72 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 9.703 2.571 9.737 ;
      VIA 2.526 9.72 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 9.72 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 9.18 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 9.163 2.571 9.197 ;
      VIA 2.526 9.18 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 9.18 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 8.64 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 8.623 2.571 8.657 ;
      VIA 2.526 8.64 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 8.64 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 8.1 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 8.083 2.571 8.117 ;
      VIA 2.526 8.1 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 8.1 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 7.56 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 7.543 2.571 7.577 ;
      VIA 2.526 7.56 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 7.56 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 7.02 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 7.003 2.571 7.037 ;
      VIA 2.526 7.02 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 7.02 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 6.48 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 6.463 2.571 6.497 ;
      VIA 2.526 6.48 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 6.48 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 5.94 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 5.923 2.571 5.957 ;
      VIA 2.526 5.94 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 5.94 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 5.4 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 5.383 2.571 5.417 ;
      VIA 2.526 5.4 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 5.4 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 4.86 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 4.843 2.571 4.877 ;
      VIA 2.526 4.86 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 4.86 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 4.32 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 4.303 2.571 4.337 ;
      VIA 2.526 4.32 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 4.32 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 3.78 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 3.763 2.571 3.797 ;
      VIA 2.526 3.78 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 3.78 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 3.24 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 3.223 2.571 3.257 ;
      VIA 2.526 3.24 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 3.24 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 2.7 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 2.683 2.571 2.717 ;
      VIA 2.526 2.7 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 2.7 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 2.16 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 2.143 2.571 2.177 ;
      VIA 2.526 2.16 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 2.16 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 1.62 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 1.603 2.571 1.637 ;
      VIA 2.526 1.62 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 1.62 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.526 1.08 fakeram7_256x32_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.481 1.063 2.571 1.097 ;
      VIA 2.526 1.08 fakeram7_256x32_VIA34_1_2_58_52 ;
      VIA 2.526 1.08 fakeram7_256x32_VIA23_1_3_36_36 ;
      VIA 2.592 25.92 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 25.38 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 24.84 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 24.3 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 23.76 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 23.22 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 22.68 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 22.14 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 21.6 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 21.06 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 20.52 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 19.98 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 19.44 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 18.9 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 18.36 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 17.82 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 17.28 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 16.74 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 16.2 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 15.66 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 15.12 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 14.58 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 14.04 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 13.5 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 12.96 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 12.42 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 11.88 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 11.34 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 10.8 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 10.26 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 9.72 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 9.18 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 8.64 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 8.1 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 7.56 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 7.02 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 6.48 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 5.94 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 5.4 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 4.86 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 4.32 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 3.78 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 3.24 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 2.7 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 2.16 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 1.62 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
      VIA 2.592 1.08 fakeram7_256x32_via1_2_3132_18_1_87_36_36 ;
    END
  END VSS
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 10.656 5.163 10.68 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 11.808 5.163 11.832 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 0.864 5.163 0.888 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 1.152 5.163 1.176 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 1.44 5.163 1.464 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 1.728 5.163 1.752 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 2.016 5.163 2.04 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 2.304 5.163 2.328 ;
    END
  END addr_in[7]
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 10.944 5.163 10.968 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 23.616 5.163 23.64 ;
    END
  END clk
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 4.32 5.163 4.344 ;
    END
  END rd_out[0]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 4.896 5.163 4.92 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 6.336 5.163 6.36 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 7.488 5.163 7.512 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 7.776 5.163 7.8 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 6.624 5.163 6.648 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 5.76 5.163 5.784 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 5.472 5.163 5.496 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 9.504 5.163 9.528 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 9.792 5.163 9.816 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 12.096 5.163 12.12 ;
    END
  END rd_out[19]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 13.248 5.163 13.272 ;
    END
  END rd_out[1]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 17.28 5.163 17.304 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 16.704 5.163 16.728 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 15.552 5.163 15.576 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 14.976 5.163 15 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 14.688 5.163 14.712 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 17.568 5.163 17.592 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 17.856 5.163 17.88 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 19.008 5.163 19.032 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 19.872 5.163 19.896 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 21.024 5.163 21.048 ;
    END
  END rd_out[29]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 22.752 5.163 22.776 ;
    END
  END rd_out[2]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 19.584 5.163 19.608 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 19.296 5.163 19.32 ;
    END
  END rd_out[31]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 23.04 5.163 23.064 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 22.464 5.163 22.488 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 22.176 5.163 22.2 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 12.672 5.163 12.696 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 14.4 5.163 14.424 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 8.64 5.163 8.664 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 8.928 5.163 8.952 ;
    END
  END rd_out[9]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 9.216 5.163 9.24 ;
    END
  END wd_in[0]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 5.184 5.163 5.208 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 8.064 5.163 8.088 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 6.912 5.163 6.936 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 8.352 5.163 8.376 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 7.2 5.163 7.224 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 4.608 5.163 4.632 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 6.048 5.163 6.072 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 11.52 5.163 11.544 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 11.232 5.163 11.256 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 12.384 5.163 12.408 ;
    END
  END wd_in[19]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 13.536 5.163 13.56 ;
    END
  END wd_in[1]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 16.128 5.163 16.152 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 16.992 5.163 17.016 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 15.264 5.163 15.288 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 15.84 5.163 15.864 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 14.112 5.163 14.136 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 16.416 5.163 16.44 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 18.144 5.163 18.168 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 18.432 5.163 18.456 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 20.448 5.163 20.472 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 20.16 5.163 20.184 ;
    END
  END wd_in[29]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 21.888 5.163 21.912 ;
    END
  END wd_in[2]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 20.736 5.163 20.76 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 18.72 5.163 18.744 ;
    END
  END wd_in[31]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 21.6 5.163 21.624 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 21.312 5.163 21.336 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 23.328 5.163 23.352 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 12.96 5.163 12.984 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 13.824 5.163 13.848 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 10.368 5.163 10.392 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 10.08 5.163 10.104 ;
    END
  END wd_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  5.079 2.592 5.163 2.616 ;
    END
  END we_in
  OBS
    LAYER M1 ;
     RECT  0.63 0.684 5.163 26.586 ;
    LAYER M2 ;
     RECT  0.63 0.684 5.163 26.586 ;
    LAYER M3 ;
     RECT  0.63 0.684 5.163 26.586 ;
    LAYER M4 ;
     RECT  0.63 0.684 5.163 26.586 ;
    LAYER M5 ;
     RECT  0.63 0.684 5.163 26.586 ;
  END
END fakeram7_256x32
END LIBRARY
