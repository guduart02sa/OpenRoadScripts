VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA ibex_ex_block_via2_3_1600_480_1_5_320_320
  VIARULE M1M2_PR ;
  CUTSIZE 0.15 0.15 ;
  LAYERS met1 via met2 ;
  CUTSPACING 0.17 0.17 ;
  ENCLOSURE 0.085 0.165 0.055 0.085 ;
  ROWCOL 1 5 ;
END ibex_ex_block_via2_3_1600_480_1_5_320_320

VIA ibex_ex_block_via3_4_1600_480_1_4_400_400
  VIARULE M2M3_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met2 via2 met3 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.04 0.085 0.065 0.065 ;
  ROWCOL 1 4 ;
END ibex_ex_block_via3_4_1600_480_1_4_400_400

VIA ibex_ex_block_via4_5_1600_480_1_4_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.06 0.1 0.065 ;
  ROWCOL 1 4 ;
END ibex_ex_block_via4_5_1600_480_1_4_400_400

VIA ibex_ex_block_via5_6_1600_1600_1_1_1600_1600
  VIARULE M4M5_PR ;
  CUTSIZE 0.8 0.8 ;
  LAYERS met4 via4 met5 ;
  CUTSPACING 0.8 0.8 ;
  ENCLOSURE 0.4 0.19 0.31 0.4 ;
END ibex_ex_block_via5_6_1600_1600_1_1_1600_1600

MACRO ibex_ex_block
  FOREIGN ibex_ex_block 0 0 ;
  CLASS BLOCK ;
  SIZE 262.08 BY 782.24 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  27.78 764.13 246.5 765.73 ;
        RECT  27.78 736.93 246.5 738.53 ;
        RECT  27.78 709.73 246.5 711.33 ;
        RECT  27.78 682.53 246.5 684.13 ;
        RECT  27.78 655.33 246.5 656.93 ;
        RECT  27.78 628.13 246.5 629.73 ;
        RECT  27.78 600.93 246.5 602.53 ;
        RECT  27.78 573.73 246.5 575.33 ;
        RECT  27.78 546.53 246.5 548.13 ;
        RECT  27.78 519.33 246.5 520.93 ;
        RECT  27.78 492.13 246.5 493.73 ;
        RECT  27.78 464.93 246.5 466.53 ;
        RECT  27.78 437.73 246.5 439.33 ;
        RECT  27.78 410.53 246.5 412.13 ;
        RECT  27.78 383.33 246.5 384.93 ;
        RECT  27.78 356.13 246.5 357.73 ;
        RECT  27.78 328.93 246.5 330.53 ;
        RECT  27.78 301.73 246.5 303.33 ;
        RECT  27.78 274.53 246.5 276.13 ;
        RECT  27.78 247.33 246.5 248.93 ;
        RECT  27.78 220.13 246.5 221.73 ;
        RECT  27.78 192.93 246.5 194.53 ;
        RECT  27.78 165.73 246.5 167.33 ;
        RECT  27.78 138.53 246.5 140.13 ;
        RECT  27.78 111.33 246.5 112.93 ;
        RECT  27.78 84.13 246.5 85.73 ;
        RECT  27.78 56.93 246.5 58.53 ;
        RECT  27.78 29.73 246.5 31.33 ;
      LAYER met4 ;
        RECT  244.9 6.42 246.5 779.46 ;
        RECT  217.76 6.42 219.36 779.46 ;
        RECT  190.62 6.42 192.22 779.46 ;
        RECT  163.48 6.42 165.08 779.46 ;
        RECT  136.34 6.42 137.94 779.46 ;
        RECT  109.2 6.42 110.8 779.46 ;
        RECT  82.06 6.42 83.66 779.46 ;
        RECT  54.92 6.42 56.52 779.46 ;
        RECT  27.78 6.42 29.38 779.46 ;
      LAYER met1 ;
        RECT  1.44 778.98 260.64 779.46 ;
        RECT  1.44 772.32 260.64 772.8 ;
        RECT  1.44 765.66 260.64 766.14 ;
        RECT  1.44 759 260.64 759.48 ;
        RECT  1.44 752.34 260.64 752.82 ;
        RECT  1.44 745.68 260.64 746.16 ;
        RECT  1.44 739.02 260.64 739.5 ;
        RECT  1.44 732.36 260.64 732.84 ;
        RECT  1.44 725.7 260.64 726.18 ;
        RECT  1.44 719.04 260.64 719.52 ;
        RECT  1.44 712.38 260.64 712.86 ;
        RECT  1.44 705.72 260.64 706.2 ;
        RECT  1.44 699.06 260.64 699.54 ;
        RECT  1.44 692.4 260.64 692.88 ;
        RECT  1.44 685.74 260.64 686.22 ;
        RECT  1.44 679.08 260.64 679.56 ;
        RECT  1.44 672.42 260.64 672.9 ;
        RECT  1.44 665.76 260.64 666.24 ;
        RECT  1.44 659.1 260.64 659.58 ;
        RECT  1.44 652.44 260.64 652.92 ;
        RECT  1.44 645.78 260.64 646.26 ;
        RECT  1.44 639.12 260.64 639.6 ;
        RECT  1.44 632.46 260.64 632.94 ;
        RECT  1.44 625.8 260.64 626.28 ;
        RECT  1.44 619.14 260.64 619.62 ;
        RECT  1.44 612.48 260.64 612.96 ;
        RECT  1.44 605.82 260.64 606.3 ;
        RECT  1.44 599.16 260.64 599.64 ;
        RECT  1.44 592.5 260.64 592.98 ;
        RECT  1.44 585.84 260.64 586.32 ;
        RECT  1.44 579.18 260.64 579.66 ;
        RECT  1.44 572.52 260.64 573 ;
        RECT  1.44 565.86 260.64 566.34 ;
        RECT  1.44 559.2 260.64 559.68 ;
        RECT  1.44 552.54 260.64 553.02 ;
        RECT  1.44 545.88 260.64 546.36 ;
        RECT  1.44 539.22 260.64 539.7 ;
        RECT  1.44 532.56 260.64 533.04 ;
        RECT  1.44 525.9 260.64 526.38 ;
        RECT  1.44 519.24 260.64 519.72 ;
        RECT  1.44 512.58 260.64 513.06 ;
        RECT  1.44 505.92 260.64 506.4 ;
        RECT  1.44 499.26 260.64 499.74 ;
        RECT  1.44 492.6 260.64 493.08 ;
        RECT  1.44 485.94 260.64 486.42 ;
        RECT  1.44 479.28 260.64 479.76 ;
        RECT  1.44 472.62 260.64 473.1 ;
        RECT  1.44 465.96 260.64 466.44 ;
        RECT  1.44 459.3 260.64 459.78 ;
        RECT  1.44 452.64 260.64 453.12 ;
        RECT  1.44 445.98 260.64 446.46 ;
        RECT  1.44 439.32 260.64 439.8 ;
        RECT  1.44 432.66 260.64 433.14 ;
        RECT  1.44 426 260.64 426.48 ;
        RECT  1.44 419.34 260.64 419.82 ;
        RECT  1.44 412.68 260.64 413.16 ;
        RECT  1.44 406.02 260.64 406.5 ;
        RECT  1.44 399.36 260.64 399.84 ;
        RECT  1.44 392.7 260.64 393.18 ;
        RECT  1.44 386.04 260.64 386.52 ;
        RECT  1.44 379.38 260.64 379.86 ;
        RECT  1.44 372.72 260.64 373.2 ;
        RECT  1.44 366.06 260.64 366.54 ;
        RECT  1.44 359.4 260.64 359.88 ;
        RECT  1.44 352.74 260.64 353.22 ;
        RECT  1.44 346.08 260.64 346.56 ;
        RECT  1.44 339.42 260.64 339.9 ;
        RECT  1.44 332.76 260.64 333.24 ;
        RECT  1.44 326.1 260.64 326.58 ;
        RECT  1.44 319.44 260.64 319.92 ;
        RECT  1.44 312.78 260.64 313.26 ;
        RECT  1.44 306.12 260.64 306.6 ;
        RECT  1.44 299.46 260.64 299.94 ;
        RECT  1.44 292.8 260.64 293.28 ;
        RECT  1.44 286.14 260.64 286.62 ;
        RECT  1.44 279.48 260.64 279.96 ;
        RECT  1.44 272.82 260.64 273.3 ;
        RECT  1.44 266.16 260.64 266.64 ;
        RECT  1.44 259.5 260.64 259.98 ;
        RECT  1.44 252.84 260.64 253.32 ;
        RECT  1.44 246.18 260.64 246.66 ;
        RECT  1.44 239.52 260.64 240 ;
        RECT  1.44 232.86 260.64 233.34 ;
        RECT  1.44 226.2 260.64 226.68 ;
        RECT  1.44 219.54 260.64 220.02 ;
        RECT  1.44 212.88 260.64 213.36 ;
        RECT  1.44 206.22 260.64 206.7 ;
        RECT  1.44 199.56 260.64 200.04 ;
        RECT  1.44 192.9 260.64 193.38 ;
        RECT  1.44 186.24 260.64 186.72 ;
        RECT  1.44 179.58 260.64 180.06 ;
        RECT  1.44 172.92 260.64 173.4 ;
        RECT  1.44 166.26 260.64 166.74 ;
        RECT  1.44 159.6 260.64 160.08 ;
        RECT  1.44 152.94 260.64 153.42 ;
        RECT  1.44 146.28 260.64 146.76 ;
        RECT  1.44 139.62 260.64 140.1 ;
        RECT  1.44 132.96 260.64 133.44 ;
        RECT  1.44 126.3 260.64 126.78 ;
        RECT  1.44 119.64 260.64 120.12 ;
        RECT  1.44 112.98 260.64 113.46 ;
        RECT  1.44 106.32 260.64 106.8 ;
        RECT  1.44 99.66 260.64 100.14 ;
        RECT  1.44 93 260.64 93.48 ;
        RECT  1.44 86.34 260.64 86.82 ;
        RECT  1.44 79.68 260.64 80.16 ;
        RECT  1.44 73.02 260.64 73.5 ;
        RECT  1.44 66.36 260.64 66.84 ;
        RECT  1.44 59.7 260.64 60.18 ;
        RECT  1.44 53.04 260.64 53.52 ;
        RECT  1.44 46.38 260.64 46.86 ;
        RECT  1.44 39.72 260.64 40.2 ;
        RECT  1.44 33.06 260.64 33.54 ;
        RECT  1.44 26.4 260.64 26.88 ;
        RECT  1.44 19.74 260.64 20.22 ;
        RECT  1.44 13.08 260.64 13.56 ;
        RECT  1.44 6.42 260.64 6.9 ;
      VIA 245.7 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 245.7 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 218.56 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 191.42 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.28 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.14 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 110 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.86 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.72 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 764.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 737.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 710.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 683.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 656.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 628.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 601.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 574.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 547.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 520.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 492.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 465.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 438.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 411.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 384.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 356.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 329.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 302.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 275.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 248.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 220.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 193.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 166.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 139.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 112.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 84.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 57.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.58 30.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  244.91 779.055 246.49 779.385 ;
      VIA 245.7 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 779.035 246.47 779.405 ;
      VIA 245.7 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 772.395 246.49 772.725 ;
      VIA 245.7 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 772.375 246.47 772.745 ;
      VIA 245.7 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 765.735 246.49 766.065 ;
      VIA 245.7 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 765.715 246.47 766.085 ;
      VIA 245.7 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 759.075 246.49 759.405 ;
      VIA 245.7 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 759.055 246.47 759.425 ;
      VIA 245.7 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 752.415 246.49 752.745 ;
      VIA 245.7 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 752.395 246.47 752.765 ;
      VIA 245.7 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 745.755 246.49 746.085 ;
      VIA 245.7 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 745.735 246.47 746.105 ;
      VIA 245.7 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 739.095 246.49 739.425 ;
      VIA 245.7 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 739.075 246.47 739.445 ;
      VIA 245.7 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 732.435 246.49 732.765 ;
      VIA 245.7 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 732.415 246.47 732.785 ;
      VIA 245.7 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 725.775 246.49 726.105 ;
      VIA 245.7 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 725.755 246.47 726.125 ;
      VIA 245.7 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 719.115 246.49 719.445 ;
      VIA 245.7 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 719.095 246.47 719.465 ;
      VIA 245.7 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 712.455 246.49 712.785 ;
      VIA 245.7 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 712.435 246.47 712.805 ;
      VIA 245.7 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 705.795 246.49 706.125 ;
      VIA 245.7 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 705.775 246.47 706.145 ;
      VIA 245.7 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 699.135 246.49 699.465 ;
      VIA 245.7 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 699.115 246.47 699.485 ;
      VIA 245.7 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 692.475 246.49 692.805 ;
      VIA 245.7 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 692.455 246.47 692.825 ;
      VIA 245.7 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 685.815 246.49 686.145 ;
      VIA 245.7 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 685.795 246.47 686.165 ;
      VIA 245.7 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 679.155 246.49 679.485 ;
      VIA 245.7 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 679.135 246.47 679.505 ;
      VIA 245.7 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 672.495 246.49 672.825 ;
      VIA 245.7 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 672.475 246.47 672.845 ;
      VIA 245.7 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 665.835 246.49 666.165 ;
      VIA 245.7 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 665.815 246.47 666.185 ;
      VIA 245.7 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 659.175 246.49 659.505 ;
      VIA 245.7 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 659.155 246.47 659.525 ;
      VIA 245.7 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 652.515 246.49 652.845 ;
      VIA 245.7 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 652.495 246.47 652.865 ;
      VIA 245.7 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 645.855 246.49 646.185 ;
      VIA 245.7 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 645.835 246.47 646.205 ;
      VIA 245.7 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 639.195 246.49 639.525 ;
      VIA 245.7 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 639.175 246.47 639.545 ;
      VIA 245.7 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 632.535 246.49 632.865 ;
      VIA 245.7 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 632.515 246.47 632.885 ;
      VIA 245.7 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 625.875 246.49 626.205 ;
      VIA 245.7 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 625.855 246.47 626.225 ;
      VIA 245.7 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 619.215 246.49 619.545 ;
      VIA 245.7 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 619.195 246.47 619.565 ;
      VIA 245.7 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 612.555 246.49 612.885 ;
      VIA 245.7 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 612.535 246.47 612.905 ;
      VIA 245.7 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 605.895 246.49 606.225 ;
      VIA 245.7 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 605.875 246.47 606.245 ;
      VIA 245.7 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 599.235 246.49 599.565 ;
      VIA 245.7 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 599.215 246.47 599.585 ;
      VIA 245.7 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 592.575 246.49 592.905 ;
      VIA 245.7 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 592.555 246.47 592.925 ;
      VIA 245.7 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 585.915 246.49 586.245 ;
      VIA 245.7 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 585.895 246.47 586.265 ;
      VIA 245.7 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 579.255 246.49 579.585 ;
      VIA 245.7 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 579.235 246.47 579.605 ;
      VIA 245.7 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 572.595 246.49 572.925 ;
      VIA 245.7 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 572.575 246.47 572.945 ;
      VIA 245.7 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 565.935 246.49 566.265 ;
      VIA 245.7 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 565.915 246.47 566.285 ;
      VIA 245.7 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 559.275 246.49 559.605 ;
      VIA 245.7 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 559.255 246.47 559.625 ;
      VIA 245.7 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 552.615 246.49 552.945 ;
      VIA 245.7 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 552.595 246.47 552.965 ;
      VIA 245.7 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 545.955 246.49 546.285 ;
      VIA 245.7 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 545.935 246.47 546.305 ;
      VIA 245.7 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 539.295 246.49 539.625 ;
      VIA 245.7 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 539.275 246.47 539.645 ;
      VIA 245.7 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 532.635 246.49 532.965 ;
      VIA 245.7 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 532.615 246.47 532.985 ;
      VIA 245.7 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 525.975 246.49 526.305 ;
      VIA 245.7 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 525.955 246.47 526.325 ;
      VIA 245.7 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 519.315 246.49 519.645 ;
      VIA 245.7 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 519.295 246.47 519.665 ;
      VIA 245.7 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 512.655 246.49 512.985 ;
      VIA 245.7 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 512.635 246.47 513.005 ;
      VIA 245.7 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 505.995 246.49 506.325 ;
      VIA 245.7 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 505.975 246.47 506.345 ;
      VIA 245.7 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 499.335 246.49 499.665 ;
      VIA 245.7 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 499.315 246.47 499.685 ;
      VIA 245.7 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 492.675 246.49 493.005 ;
      VIA 245.7 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 492.655 246.47 493.025 ;
      VIA 245.7 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 486.015 246.49 486.345 ;
      VIA 245.7 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 485.995 246.47 486.365 ;
      VIA 245.7 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 479.355 246.49 479.685 ;
      VIA 245.7 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 479.335 246.47 479.705 ;
      VIA 245.7 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 472.695 246.49 473.025 ;
      VIA 245.7 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 472.675 246.47 473.045 ;
      VIA 245.7 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 466.035 246.49 466.365 ;
      VIA 245.7 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 466.015 246.47 466.385 ;
      VIA 245.7 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 459.375 246.49 459.705 ;
      VIA 245.7 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 459.355 246.47 459.725 ;
      VIA 245.7 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 452.715 246.49 453.045 ;
      VIA 245.7 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 452.695 246.47 453.065 ;
      VIA 245.7 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 446.055 246.49 446.385 ;
      VIA 245.7 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 446.035 246.47 446.405 ;
      VIA 245.7 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 439.395 246.49 439.725 ;
      VIA 245.7 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 439.375 246.47 439.745 ;
      VIA 245.7 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 432.735 246.49 433.065 ;
      VIA 245.7 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 432.715 246.47 433.085 ;
      VIA 245.7 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 426.075 246.49 426.405 ;
      VIA 245.7 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 426.055 246.47 426.425 ;
      VIA 245.7 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 419.415 246.49 419.745 ;
      VIA 245.7 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 419.395 246.47 419.765 ;
      VIA 245.7 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 412.755 246.49 413.085 ;
      VIA 245.7 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 412.735 246.47 413.105 ;
      VIA 245.7 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 406.095 246.49 406.425 ;
      VIA 245.7 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 406.075 246.47 406.445 ;
      VIA 245.7 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 399.435 246.49 399.765 ;
      VIA 245.7 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 399.415 246.47 399.785 ;
      VIA 245.7 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 392.775 246.49 393.105 ;
      VIA 245.7 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 392.755 246.47 393.125 ;
      VIA 245.7 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 386.115 246.49 386.445 ;
      VIA 245.7 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 386.095 246.47 386.465 ;
      VIA 245.7 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 379.455 246.49 379.785 ;
      VIA 245.7 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 379.435 246.47 379.805 ;
      VIA 245.7 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 372.795 246.49 373.125 ;
      VIA 245.7 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 372.775 246.47 373.145 ;
      VIA 245.7 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 366.135 246.49 366.465 ;
      VIA 245.7 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 366.115 246.47 366.485 ;
      VIA 245.7 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 359.475 246.49 359.805 ;
      VIA 245.7 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 359.455 246.47 359.825 ;
      VIA 245.7 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 352.815 246.49 353.145 ;
      VIA 245.7 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 352.795 246.47 353.165 ;
      VIA 245.7 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 346.155 246.49 346.485 ;
      VIA 245.7 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 346.135 246.47 346.505 ;
      VIA 245.7 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 339.495 246.49 339.825 ;
      VIA 245.7 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 339.475 246.47 339.845 ;
      VIA 245.7 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 332.835 246.49 333.165 ;
      VIA 245.7 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 332.815 246.47 333.185 ;
      VIA 245.7 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 326.175 246.49 326.505 ;
      VIA 245.7 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 326.155 246.47 326.525 ;
      VIA 245.7 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 319.515 246.49 319.845 ;
      VIA 245.7 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 319.495 246.47 319.865 ;
      VIA 245.7 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 312.855 246.49 313.185 ;
      VIA 245.7 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 312.835 246.47 313.205 ;
      VIA 245.7 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 306.195 246.49 306.525 ;
      VIA 245.7 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 306.175 246.47 306.545 ;
      VIA 245.7 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 299.535 246.49 299.865 ;
      VIA 245.7 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 299.515 246.47 299.885 ;
      VIA 245.7 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 292.875 246.49 293.205 ;
      VIA 245.7 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 292.855 246.47 293.225 ;
      VIA 245.7 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 286.215 246.49 286.545 ;
      VIA 245.7 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 286.195 246.47 286.565 ;
      VIA 245.7 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 279.555 246.49 279.885 ;
      VIA 245.7 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 279.535 246.47 279.905 ;
      VIA 245.7 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 272.895 246.49 273.225 ;
      VIA 245.7 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 272.875 246.47 273.245 ;
      VIA 245.7 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 266.235 246.49 266.565 ;
      VIA 245.7 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 266.215 246.47 266.585 ;
      VIA 245.7 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 259.575 246.49 259.905 ;
      VIA 245.7 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 259.555 246.47 259.925 ;
      VIA 245.7 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 252.915 246.49 253.245 ;
      VIA 245.7 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 252.895 246.47 253.265 ;
      VIA 245.7 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 246.255 246.49 246.585 ;
      VIA 245.7 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 246.235 246.47 246.605 ;
      VIA 245.7 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 239.595 246.49 239.925 ;
      VIA 245.7 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 239.575 246.47 239.945 ;
      VIA 245.7 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 232.935 246.49 233.265 ;
      VIA 245.7 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 232.915 246.47 233.285 ;
      VIA 245.7 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 226.275 246.49 226.605 ;
      VIA 245.7 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 226.255 246.47 226.625 ;
      VIA 245.7 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 219.615 246.49 219.945 ;
      VIA 245.7 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 219.595 246.47 219.965 ;
      VIA 245.7 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 212.955 246.49 213.285 ;
      VIA 245.7 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 212.935 246.47 213.305 ;
      VIA 245.7 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 206.295 246.49 206.625 ;
      VIA 245.7 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 206.275 246.47 206.645 ;
      VIA 245.7 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 199.635 246.49 199.965 ;
      VIA 245.7 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 199.615 246.47 199.985 ;
      VIA 245.7 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 192.975 246.49 193.305 ;
      VIA 245.7 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 192.955 246.47 193.325 ;
      VIA 245.7 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 186.315 246.49 186.645 ;
      VIA 245.7 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 186.295 246.47 186.665 ;
      VIA 245.7 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 179.655 246.49 179.985 ;
      VIA 245.7 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 179.635 246.47 180.005 ;
      VIA 245.7 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 172.995 246.49 173.325 ;
      VIA 245.7 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 172.975 246.47 173.345 ;
      VIA 245.7 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 166.335 246.49 166.665 ;
      VIA 245.7 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 166.315 246.47 166.685 ;
      VIA 245.7 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 159.675 246.49 160.005 ;
      VIA 245.7 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 159.655 246.47 160.025 ;
      VIA 245.7 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 153.015 246.49 153.345 ;
      VIA 245.7 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 152.995 246.47 153.365 ;
      VIA 245.7 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 146.355 246.49 146.685 ;
      VIA 245.7 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 146.335 246.47 146.705 ;
      VIA 245.7 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 139.695 246.49 140.025 ;
      VIA 245.7 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 139.675 246.47 140.045 ;
      VIA 245.7 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 133.035 246.49 133.365 ;
      VIA 245.7 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 133.015 246.47 133.385 ;
      VIA 245.7 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 126.375 246.49 126.705 ;
      VIA 245.7 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 126.355 246.47 126.725 ;
      VIA 245.7 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 119.715 246.49 120.045 ;
      VIA 245.7 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 119.695 246.47 120.065 ;
      VIA 245.7 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 113.055 246.49 113.385 ;
      VIA 245.7 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 113.035 246.47 113.405 ;
      VIA 245.7 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 106.395 246.49 106.725 ;
      VIA 245.7 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 106.375 246.47 106.745 ;
      VIA 245.7 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 99.735 246.49 100.065 ;
      VIA 245.7 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 99.715 246.47 100.085 ;
      VIA 245.7 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 93.075 246.49 93.405 ;
      VIA 245.7 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 93.055 246.47 93.425 ;
      VIA 245.7 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 86.415 246.49 86.745 ;
      VIA 245.7 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 86.395 246.47 86.765 ;
      VIA 245.7 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 79.755 246.49 80.085 ;
      VIA 245.7 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 79.735 246.47 80.105 ;
      VIA 245.7 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 73.095 246.49 73.425 ;
      VIA 245.7 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 73.075 246.47 73.445 ;
      VIA 245.7 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 66.435 246.49 66.765 ;
      VIA 245.7 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 66.415 246.47 66.785 ;
      VIA 245.7 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 59.775 246.49 60.105 ;
      VIA 245.7 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 59.755 246.47 60.125 ;
      VIA 245.7 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 53.115 246.49 53.445 ;
      VIA 245.7 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 53.095 246.47 53.465 ;
      VIA 245.7 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 46.455 246.49 46.785 ;
      VIA 245.7 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 46.435 246.47 46.805 ;
      VIA 245.7 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 39.795 246.49 40.125 ;
      VIA 245.7 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 39.775 246.47 40.145 ;
      VIA 245.7 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 33.135 246.49 33.465 ;
      VIA 245.7 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 33.115 246.47 33.485 ;
      VIA 245.7 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 26.475 246.49 26.805 ;
      VIA 245.7 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 26.455 246.47 26.825 ;
      VIA 245.7 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 19.815 246.49 20.145 ;
      VIA 245.7 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 19.795 246.47 20.165 ;
      VIA 245.7 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 13.155 246.49 13.485 ;
      VIA 245.7 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 13.135 246.47 13.505 ;
      VIA 245.7 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  244.91 6.495 246.49 6.825 ;
      VIA 245.7 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  244.93 6.475 246.47 6.845 ;
      VIA 245.7 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 245.7 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 779.055 219.35 779.385 ;
      VIA 218.56 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 779.035 219.33 779.405 ;
      VIA 218.56 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 772.395 219.35 772.725 ;
      VIA 218.56 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 772.375 219.33 772.745 ;
      VIA 218.56 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 765.735 219.35 766.065 ;
      VIA 218.56 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 765.715 219.33 766.085 ;
      VIA 218.56 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 759.075 219.35 759.405 ;
      VIA 218.56 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 759.055 219.33 759.425 ;
      VIA 218.56 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 752.415 219.35 752.745 ;
      VIA 218.56 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 752.395 219.33 752.765 ;
      VIA 218.56 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 745.755 219.35 746.085 ;
      VIA 218.56 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 745.735 219.33 746.105 ;
      VIA 218.56 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 739.095 219.35 739.425 ;
      VIA 218.56 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 739.075 219.33 739.445 ;
      VIA 218.56 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 732.435 219.35 732.765 ;
      VIA 218.56 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 732.415 219.33 732.785 ;
      VIA 218.56 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 725.775 219.35 726.105 ;
      VIA 218.56 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 725.755 219.33 726.125 ;
      VIA 218.56 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 719.115 219.35 719.445 ;
      VIA 218.56 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 719.095 219.33 719.465 ;
      VIA 218.56 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 712.455 219.35 712.785 ;
      VIA 218.56 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 712.435 219.33 712.805 ;
      VIA 218.56 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 705.795 219.35 706.125 ;
      VIA 218.56 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 705.775 219.33 706.145 ;
      VIA 218.56 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 699.135 219.35 699.465 ;
      VIA 218.56 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 699.115 219.33 699.485 ;
      VIA 218.56 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 692.475 219.35 692.805 ;
      VIA 218.56 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 692.455 219.33 692.825 ;
      VIA 218.56 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 685.815 219.35 686.145 ;
      VIA 218.56 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 685.795 219.33 686.165 ;
      VIA 218.56 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 679.155 219.35 679.485 ;
      VIA 218.56 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 679.135 219.33 679.505 ;
      VIA 218.56 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 672.495 219.35 672.825 ;
      VIA 218.56 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 672.475 219.33 672.845 ;
      VIA 218.56 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 665.835 219.35 666.165 ;
      VIA 218.56 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 665.815 219.33 666.185 ;
      VIA 218.56 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 659.175 219.35 659.505 ;
      VIA 218.56 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 659.155 219.33 659.525 ;
      VIA 218.56 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 652.515 219.35 652.845 ;
      VIA 218.56 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 652.495 219.33 652.865 ;
      VIA 218.56 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 645.855 219.35 646.185 ;
      VIA 218.56 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 645.835 219.33 646.205 ;
      VIA 218.56 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 639.195 219.35 639.525 ;
      VIA 218.56 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 639.175 219.33 639.545 ;
      VIA 218.56 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 632.535 219.35 632.865 ;
      VIA 218.56 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 632.515 219.33 632.885 ;
      VIA 218.56 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 625.875 219.35 626.205 ;
      VIA 218.56 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 625.855 219.33 626.225 ;
      VIA 218.56 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 619.215 219.35 619.545 ;
      VIA 218.56 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 619.195 219.33 619.565 ;
      VIA 218.56 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 612.555 219.35 612.885 ;
      VIA 218.56 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 612.535 219.33 612.905 ;
      VIA 218.56 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 605.895 219.35 606.225 ;
      VIA 218.56 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 605.875 219.33 606.245 ;
      VIA 218.56 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 599.235 219.35 599.565 ;
      VIA 218.56 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 599.215 219.33 599.585 ;
      VIA 218.56 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 592.575 219.35 592.905 ;
      VIA 218.56 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 592.555 219.33 592.925 ;
      VIA 218.56 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 585.915 219.35 586.245 ;
      VIA 218.56 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 585.895 219.33 586.265 ;
      VIA 218.56 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 579.255 219.35 579.585 ;
      VIA 218.56 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 579.235 219.33 579.605 ;
      VIA 218.56 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 572.595 219.35 572.925 ;
      VIA 218.56 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 572.575 219.33 572.945 ;
      VIA 218.56 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 565.935 219.35 566.265 ;
      VIA 218.56 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 565.915 219.33 566.285 ;
      VIA 218.56 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 559.275 219.35 559.605 ;
      VIA 218.56 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 559.255 219.33 559.625 ;
      VIA 218.56 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 552.615 219.35 552.945 ;
      VIA 218.56 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 552.595 219.33 552.965 ;
      VIA 218.56 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 545.955 219.35 546.285 ;
      VIA 218.56 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 545.935 219.33 546.305 ;
      VIA 218.56 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 539.295 219.35 539.625 ;
      VIA 218.56 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 539.275 219.33 539.645 ;
      VIA 218.56 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 532.635 219.35 532.965 ;
      VIA 218.56 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 532.615 219.33 532.985 ;
      VIA 218.56 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 525.975 219.35 526.305 ;
      VIA 218.56 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 525.955 219.33 526.325 ;
      VIA 218.56 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 519.315 219.35 519.645 ;
      VIA 218.56 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 519.295 219.33 519.665 ;
      VIA 218.56 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 512.655 219.35 512.985 ;
      VIA 218.56 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 512.635 219.33 513.005 ;
      VIA 218.56 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 505.995 219.35 506.325 ;
      VIA 218.56 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 505.975 219.33 506.345 ;
      VIA 218.56 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 499.335 219.35 499.665 ;
      VIA 218.56 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 499.315 219.33 499.685 ;
      VIA 218.56 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 492.675 219.35 493.005 ;
      VIA 218.56 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 492.655 219.33 493.025 ;
      VIA 218.56 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 486.015 219.35 486.345 ;
      VIA 218.56 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 485.995 219.33 486.365 ;
      VIA 218.56 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 479.355 219.35 479.685 ;
      VIA 218.56 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 479.335 219.33 479.705 ;
      VIA 218.56 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 472.695 219.35 473.025 ;
      VIA 218.56 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 472.675 219.33 473.045 ;
      VIA 218.56 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 466.035 219.35 466.365 ;
      VIA 218.56 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 466.015 219.33 466.385 ;
      VIA 218.56 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 459.375 219.35 459.705 ;
      VIA 218.56 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 459.355 219.33 459.725 ;
      VIA 218.56 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 452.715 219.35 453.045 ;
      VIA 218.56 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 452.695 219.33 453.065 ;
      VIA 218.56 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 446.055 219.35 446.385 ;
      VIA 218.56 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 446.035 219.33 446.405 ;
      VIA 218.56 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 439.395 219.35 439.725 ;
      VIA 218.56 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 439.375 219.33 439.745 ;
      VIA 218.56 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 432.735 219.35 433.065 ;
      VIA 218.56 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 432.715 219.33 433.085 ;
      VIA 218.56 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 426.075 219.35 426.405 ;
      VIA 218.56 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 426.055 219.33 426.425 ;
      VIA 218.56 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 419.415 219.35 419.745 ;
      VIA 218.56 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 419.395 219.33 419.765 ;
      VIA 218.56 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 412.755 219.35 413.085 ;
      VIA 218.56 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 412.735 219.33 413.105 ;
      VIA 218.56 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 406.095 219.35 406.425 ;
      VIA 218.56 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 406.075 219.33 406.445 ;
      VIA 218.56 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 399.435 219.35 399.765 ;
      VIA 218.56 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 399.415 219.33 399.785 ;
      VIA 218.56 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 392.775 219.35 393.105 ;
      VIA 218.56 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 392.755 219.33 393.125 ;
      VIA 218.56 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 386.115 219.35 386.445 ;
      VIA 218.56 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 386.095 219.33 386.465 ;
      VIA 218.56 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 379.455 219.35 379.785 ;
      VIA 218.56 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 379.435 219.33 379.805 ;
      VIA 218.56 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 372.795 219.35 373.125 ;
      VIA 218.56 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 372.775 219.33 373.145 ;
      VIA 218.56 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 366.135 219.35 366.465 ;
      VIA 218.56 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 366.115 219.33 366.485 ;
      VIA 218.56 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 359.475 219.35 359.805 ;
      VIA 218.56 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 359.455 219.33 359.825 ;
      VIA 218.56 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 352.815 219.35 353.145 ;
      VIA 218.56 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 352.795 219.33 353.165 ;
      VIA 218.56 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 346.155 219.35 346.485 ;
      VIA 218.56 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 346.135 219.33 346.505 ;
      VIA 218.56 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 339.495 219.35 339.825 ;
      VIA 218.56 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 339.475 219.33 339.845 ;
      VIA 218.56 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 332.835 219.35 333.165 ;
      VIA 218.56 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 332.815 219.33 333.185 ;
      VIA 218.56 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 326.175 219.35 326.505 ;
      VIA 218.56 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 326.155 219.33 326.525 ;
      VIA 218.56 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 319.515 219.35 319.845 ;
      VIA 218.56 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 319.495 219.33 319.865 ;
      VIA 218.56 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 312.855 219.35 313.185 ;
      VIA 218.56 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 312.835 219.33 313.205 ;
      VIA 218.56 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 306.195 219.35 306.525 ;
      VIA 218.56 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 306.175 219.33 306.545 ;
      VIA 218.56 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 299.535 219.35 299.865 ;
      VIA 218.56 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 299.515 219.33 299.885 ;
      VIA 218.56 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 292.875 219.35 293.205 ;
      VIA 218.56 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 292.855 219.33 293.225 ;
      VIA 218.56 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 286.215 219.35 286.545 ;
      VIA 218.56 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 286.195 219.33 286.565 ;
      VIA 218.56 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 279.555 219.35 279.885 ;
      VIA 218.56 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 279.535 219.33 279.905 ;
      VIA 218.56 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 272.895 219.35 273.225 ;
      VIA 218.56 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 272.875 219.33 273.245 ;
      VIA 218.56 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 266.235 219.35 266.565 ;
      VIA 218.56 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 266.215 219.33 266.585 ;
      VIA 218.56 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 259.575 219.35 259.905 ;
      VIA 218.56 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 259.555 219.33 259.925 ;
      VIA 218.56 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 252.915 219.35 253.245 ;
      VIA 218.56 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 252.895 219.33 253.265 ;
      VIA 218.56 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 246.255 219.35 246.585 ;
      VIA 218.56 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 246.235 219.33 246.605 ;
      VIA 218.56 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 239.595 219.35 239.925 ;
      VIA 218.56 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 239.575 219.33 239.945 ;
      VIA 218.56 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 232.935 219.35 233.265 ;
      VIA 218.56 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 232.915 219.33 233.285 ;
      VIA 218.56 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 226.275 219.35 226.605 ;
      VIA 218.56 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 226.255 219.33 226.625 ;
      VIA 218.56 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 219.615 219.35 219.945 ;
      VIA 218.56 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 219.595 219.33 219.965 ;
      VIA 218.56 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 212.955 219.35 213.285 ;
      VIA 218.56 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 212.935 219.33 213.305 ;
      VIA 218.56 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 206.295 219.35 206.625 ;
      VIA 218.56 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 206.275 219.33 206.645 ;
      VIA 218.56 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 199.635 219.35 199.965 ;
      VIA 218.56 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 199.615 219.33 199.985 ;
      VIA 218.56 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 192.975 219.35 193.305 ;
      VIA 218.56 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 192.955 219.33 193.325 ;
      VIA 218.56 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 186.315 219.35 186.645 ;
      VIA 218.56 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 186.295 219.33 186.665 ;
      VIA 218.56 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 179.655 219.35 179.985 ;
      VIA 218.56 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 179.635 219.33 180.005 ;
      VIA 218.56 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 172.995 219.35 173.325 ;
      VIA 218.56 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 172.975 219.33 173.345 ;
      VIA 218.56 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 166.335 219.35 166.665 ;
      VIA 218.56 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 166.315 219.33 166.685 ;
      VIA 218.56 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 159.675 219.35 160.005 ;
      VIA 218.56 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 159.655 219.33 160.025 ;
      VIA 218.56 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 153.015 219.35 153.345 ;
      VIA 218.56 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 152.995 219.33 153.365 ;
      VIA 218.56 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 146.355 219.35 146.685 ;
      VIA 218.56 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 146.335 219.33 146.705 ;
      VIA 218.56 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 139.695 219.35 140.025 ;
      VIA 218.56 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 139.675 219.33 140.045 ;
      VIA 218.56 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 133.035 219.35 133.365 ;
      VIA 218.56 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 133.015 219.33 133.385 ;
      VIA 218.56 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 126.375 219.35 126.705 ;
      VIA 218.56 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 126.355 219.33 126.725 ;
      VIA 218.56 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 119.715 219.35 120.045 ;
      VIA 218.56 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 119.695 219.33 120.065 ;
      VIA 218.56 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 113.055 219.35 113.385 ;
      VIA 218.56 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 113.035 219.33 113.405 ;
      VIA 218.56 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 106.395 219.35 106.725 ;
      VIA 218.56 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 106.375 219.33 106.745 ;
      VIA 218.56 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 99.735 219.35 100.065 ;
      VIA 218.56 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 99.715 219.33 100.085 ;
      VIA 218.56 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 93.075 219.35 93.405 ;
      VIA 218.56 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 93.055 219.33 93.425 ;
      VIA 218.56 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 86.415 219.35 86.745 ;
      VIA 218.56 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 86.395 219.33 86.765 ;
      VIA 218.56 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 79.755 219.35 80.085 ;
      VIA 218.56 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 79.735 219.33 80.105 ;
      VIA 218.56 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 73.095 219.35 73.425 ;
      VIA 218.56 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 73.075 219.33 73.445 ;
      VIA 218.56 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 66.435 219.35 66.765 ;
      VIA 218.56 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 66.415 219.33 66.785 ;
      VIA 218.56 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 59.775 219.35 60.105 ;
      VIA 218.56 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 59.755 219.33 60.125 ;
      VIA 218.56 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 53.115 219.35 53.445 ;
      VIA 218.56 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 53.095 219.33 53.465 ;
      VIA 218.56 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 46.455 219.35 46.785 ;
      VIA 218.56 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 46.435 219.33 46.805 ;
      VIA 218.56 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 39.795 219.35 40.125 ;
      VIA 218.56 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 39.775 219.33 40.145 ;
      VIA 218.56 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 33.135 219.35 33.465 ;
      VIA 218.56 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 33.115 219.33 33.485 ;
      VIA 218.56 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 26.475 219.35 26.805 ;
      VIA 218.56 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 26.455 219.33 26.825 ;
      VIA 218.56 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 19.815 219.35 20.145 ;
      VIA 218.56 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 19.795 219.33 20.165 ;
      VIA 218.56 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 13.155 219.35 13.485 ;
      VIA 218.56 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 13.135 219.33 13.505 ;
      VIA 218.56 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  217.77 6.495 219.35 6.825 ;
      VIA 218.56 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  217.79 6.475 219.33 6.845 ;
      VIA 218.56 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 218.56 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 779.055 192.21 779.385 ;
      VIA 191.42 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 779.035 192.19 779.405 ;
      VIA 191.42 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 772.395 192.21 772.725 ;
      VIA 191.42 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 772.375 192.19 772.745 ;
      VIA 191.42 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 765.735 192.21 766.065 ;
      VIA 191.42 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 765.715 192.19 766.085 ;
      VIA 191.42 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 759.075 192.21 759.405 ;
      VIA 191.42 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 759.055 192.19 759.425 ;
      VIA 191.42 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 752.415 192.21 752.745 ;
      VIA 191.42 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 752.395 192.19 752.765 ;
      VIA 191.42 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 745.755 192.21 746.085 ;
      VIA 191.42 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 745.735 192.19 746.105 ;
      VIA 191.42 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 739.095 192.21 739.425 ;
      VIA 191.42 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 739.075 192.19 739.445 ;
      VIA 191.42 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 732.435 192.21 732.765 ;
      VIA 191.42 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 732.415 192.19 732.785 ;
      VIA 191.42 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 725.775 192.21 726.105 ;
      VIA 191.42 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 725.755 192.19 726.125 ;
      VIA 191.42 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 719.115 192.21 719.445 ;
      VIA 191.42 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 719.095 192.19 719.465 ;
      VIA 191.42 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 712.455 192.21 712.785 ;
      VIA 191.42 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 712.435 192.19 712.805 ;
      VIA 191.42 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 705.795 192.21 706.125 ;
      VIA 191.42 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 705.775 192.19 706.145 ;
      VIA 191.42 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 699.135 192.21 699.465 ;
      VIA 191.42 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 699.115 192.19 699.485 ;
      VIA 191.42 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 692.475 192.21 692.805 ;
      VIA 191.42 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 692.455 192.19 692.825 ;
      VIA 191.42 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 685.815 192.21 686.145 ;
      VIA 191.42 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 685.795 192.19 686.165 ;
      VIA 191.42 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 679.155 192.21 679.485 ;
      VIA 191.42 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 679.135 192.19 679.505 ;
      VIA 191.42 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 672.495 192.21 672.825 ;
      VIA 191.42 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 672.475 192.19 672.845 ;
      VIA 191.42 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 665.835 192.21 666.165 ;
      VIA 191.42 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 665.815 192.19 666.185 ;
      VIA 191.42 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 659.175 192.21 659.505 ;
      VIA 191.42 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 659.155 192.19 659.525 ;
      VIA 191.42 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 652.515 192.21 652.845 ;
      VIA 191.42 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 652.495 192.19 652.865 ;
      VIA 191.42 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 645.855 192.21 646.185 ;
      VIA 191.42 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 645.835 192.19 646.205 ;
      VIA 191.42 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 639.195 192.21 639.525 ;
      VIA 191.42 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 639.175 192.19 639.545 ;
      VIA 191.42 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 632.535 192.21 632.865 ;
      VIA 191.42 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 632.515 192.19 632.885 ;
      VIA 191.42 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 625.875 192.21 626.205 ;
      VIA 191.42 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 625.855 192.19 626.225 ;
      VIA 191.42 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 619.215 192.21 619.545 ;
      VIA 191.42 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 619.195 192.19 619.565 ;
      VIA 191.42 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 612.555 192.21 612.885 ;
      VIA 191.42 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 612.535 192.19 612.905 ;
      VIA 191.42 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 605.895 192.21 606.225 ;
      VIA 191.42 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 605.875 192.19 606.245 ;
      VIA 191.42 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 599.235 192.21 599.565 ;
      VIA 191.42 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 599.215 192.19 599.585 ;
      VIA 191.42 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 592.575 192.21 592.905 ;
      VIA 191.42 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 592.555 192.19 592.925 ;
      VIA 191.42 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 585.915 192.21 586.245 ;
      VIA 191.42 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 585.895 192.19 586.265 ;
      VIA 191.42 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 579.255 192.21 579.585 ;
      VIA 191.42 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 579.235 192.19 579.605 ;
      VIA 191.42 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 572.595 192.21 572.925 ;
      VIA 191.42 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 572.575 192.19 572.945 ;
      VIA 191.42 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 565.935 192.21 566.265 ;
      VIA 191.42 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 565.915 192.19 566.285 ;
      VIA 191.42 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 559.275 192.21 559.605 ;
      VIA 191.42 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 559.255 192.19 559.625 ;
      VIA 191.42 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 552.615 192.21 552.945 ;
      VIA 191.42 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 552.595 192.19 552.965 ;
      VIA 191.42 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 545.955 192.21 546.285 ;
      VIA 191.42 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 545.935 192.19 546.305 ;
      VIA 191.42 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 539.295 192.21 539.625 ;
      VIA 191.42 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 539.275 192.19 539.645 ;
      VIA 191.42 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 532.635 192.21 532.965 ;
      VIA 191.42 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 532.615 192.19 532.985 ;
      VIA 191.42 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 525.975 192.21 526.305 ;
      VIA 191.42 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 525.955 192.19 526.325 ;
      VIA 191.42 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 519.315 192.21 519.645 ;
      VIA 191.42 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 519.295 192.19 519.665 ;
      VIA 191.42 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 512.655 192.21 512.985 ;
      VIA 191.42 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 512.635 192.19 513.005 ;
      VIA 191.42 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 505.995 192.21 506.325 ;
      VIA 191.42 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 505.975 192.19 506.345 ;
      VIA 191.42 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 499.335 192.21 499.665 ;
      VIA 191.42 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 499.315 192.19 499.685 ;
      VIA 191.42 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 492.675 192.21 493.005 ;
      VIA 191.42 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 492.655 192.19 493.025 ;
      VIA 191.42 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 486.015 192.21 486.345 ;
      VIA 191.42 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 485.995 192.19 486.365 ;
      VIA 191.42 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 479.355 192.21 479.685 ;
      VIA 191.42 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 479.335 192.19 479.705 ;
      VIA 191.42 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 472.695 192.21 473.025 ;
      VIA 191.42 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 472.675 192.19 473.045 ;
      VIA 191.42 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 466.035 192.21 466.365 ;
      VIA 191.42 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 466.015 192.19 466.385 ;
      VIA 191.42 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 459.375 192.21 459.705 ;
      VIA 191.42 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 459.355 192.19 459.725 ;
      VIA 191.42 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 452.715 192.21 453.045 ;
      VIA 191.42 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 452.695 192.19 453.065 ;
      VIA 191.42 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 446.055 192.21 446.385 ;
      VIA 191.42 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 446.035 192.19 446.405 ;
      VIA 191.42 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 439.395 192.21 439.725 ;
      VIA 191.42 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 439.375 192.19 439.745 ;
      VIA 191.42 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 432.735 192.21 433.065 ;
      VIA 191.42 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 432.715 192.19 433.085 ;
      VIA 191.42 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 426.075 192.21 426.405 ;
      VIA 191.42 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 426.055 192.19 426.425 ;
      VIA 191.42 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 419.415 192.21 419.745 ;
      VIA 191.42 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 419.395 192.19 419.765 ;
      VIA 191.42 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 412.755 192.21 413.085 ;
      VIA 191.42 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 412.735 192.19 413.105 ;
      VIA 191.42 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 406.095 192.21 406.425 ;
      VIA 191.42 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 406.075 192.19 406.445 ;
      VIA 191.42 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 399.435 192.21 399.765 ;
      VIA 191.42 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 399.415 192.19 399.785 ;
      VIA 191.42 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 392.775 192.21 393.105 ;
      VIA 191.42 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 392.755 192.19 393.125 ;
      VIA 191.42 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 386.115 192.21 386.445 ;
      VIA 191.42 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 386.095 192.19 386.465 ;
      VIA 191.42 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 379.455 192.21 379.785 ;
      VIA 191.42 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 379.435 192.19 379.805 ;
      VIA 191.42 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 372.795 192.21 373.125 ;
      VIA 191.42 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 372.775 192.19 373.145 ;
      VIA 191.42 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 366.135 192.21 366.465 ;
      VIA 191.42 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 366.115 192.19 366.485 ;
      VIA 191.42 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 359.475 192.21 359.805 ;
      VIA 191.42 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 359.455 192.19 359.825 ;
      VIA 191.42 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 352.815 192.21 353.145 ;
      VIA 191.42 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 352.795 192.19 353.165 ;
      VIA 191.42 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 346.155 192.21 346.485 ;
      VIA 191.42 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 346.135 192.19 346.505 ;
      VIA 191.42 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 339.495 192.21 339.825 ;
      VIA 191.42 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 339.475 192.19 339.845 ;
      VIA 191.42 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 332.835 192.21 333.165 ;
      VIA 191.42 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 332.815 192.19 333.185 ;
      VIA 191.42 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 326.175 192.21 326.505 ;
      VIA 191.42 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 326.155 192.19 326.525 ;
      VIA 191.42 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 319.515 192.21 319.845 ;
      VIA 191.42 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 319.495 192.19 319.865 ;
      VIA 191.42 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 312.855 192.21 313.185 ;
      VIA 191.42 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 312.835 192.19 313.205 ;
      VIA 191.42 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 306.195 192.21 306.525 ;
      VIA 191.42 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 306.175 192.19 306.545 ;
      VIA 191.42 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 299.535 192.21 299.865 ;
      VIA 191.42 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 299.515 192.19 299.885 ;
      VIA 191.42 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 292.875 192.21 293.205 ;
      VIA 191.42 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 292.855 192.19 293.225 ;
      VIA 191.42 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 286.215 192.21 286.545 ;
      VIA 191.42 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 286.195 192.19 286.565 ;
      VIA 191.42 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 279.555 192.21 279.885 ;
      VIA 191.42 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 279.535 192.19 279.905 ;
      VIA 191.42 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 272.895 192.21 273.225 ;
      VIA 191.42 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 272.875 192.19 273.245 ;
      VIA 191.42 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 266.235 192.21 266.565 ;
      VIA 191.42 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 266.215 192.19 266.585 ;
      VIA 191.42 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 259.575 192.21 259.905 ;
      VIA 191.42 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 259.555 192.19 259.925 ;
      VIA 191.42 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 252.915 192.21 253.245 ;
      VIA 191.42 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 252.895 192.19 253.265 ;
      VIA 191.42 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 246.255 192.21 246.585 ;
      VIA 191.42 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 246.235 192.19 246.605 ;
      VIA 191.42 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 239.595 192.21 239.925 ;
      VIA 191.42 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 239.575 192.19 239.945 ;
      VIA 191.42 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 232.935 192.21 233.265 ;
      VIA 191.42 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 232.915 192.19 233.285 ;
      VIA 191.42 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 226.275 192.21 226.605 ;
      VIA 191.42 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 226.255 192.19 226.625 ;
      VIA 191.42 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 219.615 192.21 219.945 ;
      VIA 191.42 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 219.595 192.19 219.965 ;
      VIA 191.42 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 212.955 192.21 213.285 ;
      VIA 191.42 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 212.935 192.19 213.305 ;
      VIA 191.42 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 206.295 192.21 206.625 ;
      VIA 191.42 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 206.275 192.19 206.645 ;
      VIA 191.42 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 199.635 192.21 199.965 ;
      VIA 191.42 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 199.615 192.19 199.985 ;
      VIA 191.42 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 192.975 192.21 193.305 ;
      VIA 191.42 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 192.955 192.19 193.325 ;
      VIA 191.42 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 186.315 192.21 186.645 ;
      VIA 191.42 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 186.295 192.19 186.665 ;
      VIA 191.42 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 179.655 192.21 179.985 ;
      VIA 191.42 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 179.635 192.19 180.005 ;
      VIA 191.42 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 172.995 192.21 173.325 ;
      VIA 191.42 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 172.975 192.19 173.345 ;
      VIA 191.42 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 166.335 192.21 166.665 ;
      VIA 191.42 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 166.315 192.19 166.685 ;
      VIA 191.42 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 159.675 192.21 160.005 ;
      VIA 191.42 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 159.655 192.19 160.025 ;
      VIA 191.42 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 153.015 192.21 153.345 ;
      VIA 191.42 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 152.995 192.19 153.365 ;
      VIA 191.42 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 146.355 192.21 146.685 ;
      VIA 191.42 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 146.335 192.19 146.705 ;
      VIA 191.42 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 139.695 192.21 140.025 ;
      VIA 191.42 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 139.675 192.19 140.045 ;
      VIA 191.42 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 133.035 192.21 133.365 ;
      VIA 191.42 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 133.015 192.19 133.385 ;
      VIA 191.42 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 126.375 192.21 126.705 ;
      VIA 191.42 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 126.355 192.19 126.725 ;
      VIA 191.42 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 119.715 192.21 120.045 ;
      VIA 191.42 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 119.695 192.19 120.065 ;
      VIA 191.42 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 113.055 192.21 113.385 ;
      VIA 191.42 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 113.035 192.19 113.405 ;
      VIA 191.42 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 106.395 192.21 106.725 ;
      VIA 191.42 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 106.375 192.19 106.745 ;
      VIA 191.42 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 99.735 192.21 100.065 ;
      VIA 191.42 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 99.715 192.19 100.085 ;
      VIA 191.42 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 93.075 192.21 93.405 ;
      VIA 191.42 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 93.055 192.19 93.425 ;
      VIA 191.42 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 86.415 192.21 86.745 ;
      VIA 191.42 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 86.395 192.19 86.765 ;
      VIA 191.42 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 79.755 192.21 80.085 ;
      VIA 191.42 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 79.735 192.19 80.105 ;
      VIA 191.42 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 73.095 192.21 73.425 ;
      VIA 191.42 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 73.075 192.19 73.445 ;
      VIA 191.42 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 66.435 192.21 66.765 ;
      VIA 191.42 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 66.415 192.19 66.785 ;
      VIA 191.42 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 59.775 192.21 60.105 ;
      VIA 191.42 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 59.755 192.19 60.125 ;
      VIA 191.42 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 53.115 192.21 53.445 ;
      VIA 191.42 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 53.095 192.19 53.465 ;
      VIA 191.42 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 46.455 192.21 46.785 ;
      VIA 191.42 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 46.435 192.19 46.805 ;
      VIA 191.42 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 39.795 192.21 40.125 ;
      VIA 191.42 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 39.775 192.19 40.145 ;
      VIA 191.42 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 33.135 192.21 33.465 ;
      VIA 191.42 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 33.115 192.19 33.485 ;
      VIA 191.42 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 26.475 192.21 26.805 ;
      VIA 191.42 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 26.455 192.19 26.825 ;
      VIA 191.42 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 19.815 192.21 20.145 ;
      VIA 191.42 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 19.795 192.19 20.165 ;
      VIA 191.42 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 13.155 192.21 13.485 ;
      VIA 191.42 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 13.135 192.19 13.505 ;
      VIA 191.42 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  190.63 6.495 192.21 6.825 ;
      VIA 191.42 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  190.65 6.475 192.19 6.845 ;
      VIA 191.42 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 191.42 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 779.055 165.07 779.385 ;
      VIA 164.28 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 779.035 165.05 779.405 ;
      VIA 164.28 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 772.395 165.07 772.725 ;
      VIA 164.28 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 772.375 165.05 772.745 ;
      VIA 164.28 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 765.735 165.07 766.065 ;
      VIA 164.28 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 765.715 165.05 766.085 ;
      VIA 164.28 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 759.075 165.07 759.405 ;
      VIA 164.28 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 759.055 165.05 759.425 ;
      VIA 164.28 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 752.415 165.07 752.745 ;
      VIA 164.28 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 752.395 165.05 752.765 ;
      VIA 164.28 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 745.755 165.07 746.085 ;
      VIA 164.28 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 745.735 165.05 746.105 ;
      VIA 164.28 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 739.095 165.07 739.425 ;
      VIA 164.28 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 739.075 165.05 739.445 ;
      VIA 164.28 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 732.435 165.07 732.765 ;
      VIA 164.28 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 732.415 165.05 732.785 ;
      VIA 164.28 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 725.775 165.07 726.105 ;
      VIA 164.28 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 725.755 165.05 726.125 ;
      VIA 164.28 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 719.115 165.07 719.445 ;
      VIA 164.28 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 719.095 165.05 719.465 ;
      VIA 164.28 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 712.455 165.07 712.785 ;
      VIA 164.28 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 712.435 165.05 712.805 ;
      VIA 164.28 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 705.795 165.07 706.125 ;
      VIA 164.28 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 705.775 165.05 706.145 ;
      VIA 164.28 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 699.135 165.07 699.465 ;
      VIA 164.28 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 699.115 165.05 699.485 ;
      VIA 164.28 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 692.475 165.07 692.805 ;
      VIA 164.28 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 692.455 165.05 692.825 ;
      VIA 164.28 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 685.815 165.07 686.145 ;
      VIA 164.28 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 685.795 165.05 686.165 ;
      VIA 164.28 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 679.155 165.07 679.485 ;
      VIA 164.28 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 679.135 165.05 679.505 ;
      VIA 164.28 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 672.495 165.07 672.825 ;
      VIA 164.28 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 672.475 165.05 672.845 ;
      VIA 164.28 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 665.835 165.07 666.165 ;
      VIA 164.28 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 665.815 165.05 666.185 ;
      VIA 164.28 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 659.175 165.07 659.505 ;
      VIA 164.28 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 659.155 165.05 659.525 ;
      VIA 164.28 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 652.515 165.07 652.845 ;
      VIA 164.28 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 652.495 165.05 652.865 ;
      VIA 164.28 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 645.855 165.07 646.185 ;
      VIA 164.28 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 645.835 165.05 646.205 ;
      VIA 164.28 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 639.195 165.07 639.525 ;
      VIA 164.28 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 639.175 165.05 639.545 ;
      VIA 164.28 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 632.535 165.07 632.865 ;
      VIA 164.28 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 632.515 165.05 632.885 ;
      VIA 164.28 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 625.875 165.07 626.205 ;
      VIA 164.28 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 625.855 165.05 626.225 ;
      VIA 164.28 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 619.215 165.07 619.545 ;
      VIA 164.28 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 619.195 165.05 619.565 ;
      VIA 164.28 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 612.555 165.07 612.885 ;
      VIA 164.28 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 612.535 165.05 612.905 ;
      VIA 164.28 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 605.895 165.07 606.225 ;
      VIA 164.28 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 605.875 165.05 606.245 ;
      VIA 164.28 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 599.235 165.07 599.565 ;
      VIA 164.28 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 599.215 165.05 599.585 ;
      VIA 164.28 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 592.575 165.07 592.905 ;
      VIA 164.28 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 592.555 165.05 592.925 ;
      VIA 164.28 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 585.915 165.07 586.245 ;
      VIA 164.28 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 585.895 165.05 586.265 ;
      VIA 164.28 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 579.255 165.07 579.585 ;
      VIA 164.28 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 579.235 165.05 579.605 ;
      VIA 164.28 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 572.595 165.07 572.925 ;
      VIA 164.28 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 572.575 165.05 572.945 ;
      VIA 164.28 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 565.935 165.07 566.265 ;
      VIA 164.28 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 565.915 165.05 566.285 ;
      VIA 164.28 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 559.275 165.07 559.605 ;
      VIA 164.28 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 559.255 165.05 559.625 ;
      VIA 164.28 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 552.615 165.07 552.945 ;
      VIA 164.28 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 552.595 165.05 552.965 ;
      VIA 164.28 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 545.955 165.07 546.285 ;
      VIA 164.28 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 545.935 165.05 546.305 ;
      VIA 164.28 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 539.295 165.07 539.625 ;
      VIA 164.28 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 539.275 165.05 539.645 ;
      VIA 164.28 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 532.635 165.07 532.965 ;
      VIA 164.28 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 532.615 165.05 532.985 ;
      VIA 164.28 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 525.975 165.07 526.305 ;
      VIA 164.28 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 525.955 165.05 526.325 ;
      VIA 164.28 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 519.315 165.07 519.645 ;
      VIA 164.28 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 519.295 165.05 519.665 ;
      VIA 164.28 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 512.655 165.07 512.985 ;
      VIA 164.28 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 512.635 165.05 513.005 ;
      VIA 164.28 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 505.995 165.07 506.325 ;
      VIA 164.28 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 505.975 165.05 506.345 ;
      VIA 164.28 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 499.335 165.07 499.665 ;
      VIA 164.28 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 499.315 165.05 499.685 ;
      VIA 164.28 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 492.675 165.07 493.005 ;
      VIA 164.28 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 492.655 165.05 493.025 ;
      VIA 164.28 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 486.015 165.07 486.345 ;
      VIA 164.28 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 485.995 165.05 486.365 ;
      VIA 164.28 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 479.355 165.07 479.685 ;
      VIA 164.28 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 479.335 165.05 479.705 ;
      VIA 164.28 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 472.695 165.07 473.025 ;
      VIA 164.28 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 472.675 165.05 473.045 ;
      VIA 164.28 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 466.035 165.07 466.365 ;
      VIA 164.28 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 466.015 165.05 466.385 ;
      VIA 164.28 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 459.375 165.07 459.705 ;
      VIA 164.28 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 459.355 165.05 459.725 ;
      VIA 164.28 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 452.715 165.07 453.045 ;
      VIA 164.28 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 452.695 165.05 453.065 ;
      VIA 164.28 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 446.055 165.07 446.385 ;
      VIA 164.28 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 446.035 165.05 446.405 ;
      VIA 164.28 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 439.395 165.07 439.725 ;
      VIA 164.28 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 439.375 165.05 439.745 ;
      VIA 164.28 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 432.735 165.07 433.065 ;
      VIA 164.28 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 432.715 165.05 433.085 ;
      VIA 164.28 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 426.075 165.07 426.405 ;
      VIA 164.28 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 426.055 165.05 426.425 ;
      VIA 164.28 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 419.415 165.07 419.745 ;
      VIA 164.28 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 419.395 165.05 419.765 ;
      VIA 164.28 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 412.755 165.07 413.085 ;
      VIA 164.28 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 412.735 165.05 413.105 ;
      VIA 164.28 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 406.095 165.07 406.425 ;
      VIA 164.28 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 406.075 165.05 406.445 ;
      VIA 164.28 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 399.435 165.07 399.765 ;
      VIA 164.28 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 399.415 165.05 399.785 ;
      VIA 164.28 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 392.775 165.07 393.105 ;
      VIA 164.28 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 392.755 165.05 393.125 ;
      VIA 164.28 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 386.115 165.07 386.445 ;
      VIA 164.28 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 386.095 165.05 386.465 ;
      VIA 164.28 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 379.455 165.07 379.785 ;
      VIA 164.28 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 379.435 165.05 379.805 ;
      VIA 164.28 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 372.795 165.07 373.125 ;
      VIA 164.28 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 372.775 165.05 373.145 ;
      VIA 164.28 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 366.135 165.07 366.465 ;
      VIA 164.28 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 366.115 165.05 366.485 ;
      VIA 164.28 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 359.475 165.07 359.805 ;
      VIA 164.28 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 359.455 165.05 359.825 ;
      VIA 164.28 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 352.815 165.07 353.145 ;
      VIA 164.28 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 352.795 165.05 353.165 ;
      VIA 164.28 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 346.155 165.07 346.485 ;
      VIA 164.28 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 346.135 165.05 346.505 ;
      VIA 164.28 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 339.495 165.07 339.825 ;
      VIA 164.28 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 339.475 165.05 339.845 ;
      VIA 164.28 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 332.835 165.07 333.165 ;
      VIA 164.28 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 332.815 165.05 333.185 ;
      VIA 164.28 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 326.175 165.07 326.505 ;
      VIA 164.28 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 326.155 165.05 326.525 ;
      VIA 164.28 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 319.515 165.07 319.845 ;
      VIA 164.28 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 319.495 165.05 319.865 ;
      VIA 164.28 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 312.855 165.07 313.185 ;
      VIA 164.28 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 312.835 165.05 313.205 ;
      VIA 164.28 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 306.195 165.07 306.525 ;
      VIA 164.28 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 306.175 165.05 306.545 ;
      VIA 164.28 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 299.535 165.07 299.865 ;
      VIA 164.28 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 299.515 165.05 299.885 ;
      VIA 164.28 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 292.875 165.07 293.205 ;
      VIA 164.28 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 292.855 165.05 293.225 ;
      VIA 164.28 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 286.215 165.07 286.545 ;
      VIA 164.28 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 286.195 165.05 286.565 ;
      VIA 164.28 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 279.555 165.07 279.885 ;
      VIA 164.28 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 279.535 165.05 279.905 ;
      VIA 164.28 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 272.895 165.07 273.225 ;
      VIA 164.28 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 272.875 165.05 273.245 ;
      VIA 164.28 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 266.235 165.07 266.565 ;
      VIA 164.28 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 266.215 165.05 266.585 ;
      VIA 164.28 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 259.575 165.07 259.905 ;
      VIA 164.28 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 259.555 165.05 259.925 ;
      VIA 164.28 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 252.915 165.07 253.245 ;
      VIA 164.28 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 252.895 165.05 253.265 ;
      VIA 164.28 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 246.255 165.07 246.585 ;
      VIA 164.28 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 246.235 165.05 246.605 ;
      VIA 164.28 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 239.595 165.07 239.925 ;
      VIA 164.28 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 239.575 165.05 239.945 ;
      VIA 164.28 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 232.935 165.07 233.265 ;
      VIA 164.28 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 232.915 165.05 233.285 ;
      VIA 164.28 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 226.275 165.07 226.605 ;
      VIA 164.28 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 226.255 165.05 226.625 ;
      VIA 164.28 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 219.615 165.07 219.945 ;
      VIA 164.28 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 219.595 165.05 219.965 ;
      VIA 164.28 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 212.955 165.07 213.285 ;
      VIA 164.28 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 212.935 165.05 213.305 ;
      VIA 164.28 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 206.295 165.07 206.625 ;
      VIA 164.28 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 206.275 165.05 206.645 ;
      VIA 164.28 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 199.635 165.07 199.965 ;
      VIA 164.28 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 199.615 165.05 199.985 ;
      VIA 164.28 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 192.975 165.07 193.305 ;
      VIA 164.28 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 192.955 165.05 193.325 ;
      VIA 164.28 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 186.315 165.07 186.645 ;
      VIA 164.28 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 186.295 165.05 186.665 ;
      VIA 164.28 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 179.655 165.07 179.985 ;
      VIA 164.28 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 179.635 165.05 180.005 ;
      VIA 164.28 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 172.995 165.07 173.325 ;
      VIA 164.28 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 172.975 165.05 173.345 ;
      VIA 164.28 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 166.335 165.07 166.665 ;
      VIA 164.28 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 166.315 165.05 166.685 ;
      VIA 164.28 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 159.675 165.07 160.005 ;
      VIA 164.28 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 159.655 165.05 160.025 ;
      VIA 164.28 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 153.015 165.07 153.345 ;
      VIA 164.28 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 152.995 165.05 153.365 ;
      VIA 164.28 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 146.355 165.07 146.685 ;
      VIA 164.28 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 146.335 165.05 146.705 ;
      VIA 164.28 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 139.695 165.07 140.025 ;
      VIA 164.28 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 139.675 165.05 140.045 ;
      VIA 164.28 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 133.035 165.07 133.365 ;
      VIA 164.28 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 133.015 165.05 133.385 ;
      VIA 164.28 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 126.375 165.07 126.705 ;
      VIA 164.28 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 126.355 165.05 126.725 ;
      VIA 164.28 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 119.715 165.07 120.045 ;
      VIA 164.28 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 119.695 165.05 120.065 ;
      VIA 164.28 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 113.055 165.07 113.385 ;
      VIA 164.28 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 113.035 165.05 113.405 ;
      VIA 164.28 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 106.395 165.07 106.725 ;
      VIA 164.28 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 106.375 165.05 106.745 ;
      VIA 164.28 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 99.735 165.07 100.065 ;
      VIA 164.28 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 99.715 165.05 100.085 ;
      VIA 164.28 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 93.075 165.07 93.405 ;
      VIA 164.28 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 93.055 165.05 93.425 ;
      VIA 164.28 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 86.415 165.07 86.745 ;
      VIA 164.28 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 86.395 165.05 86.765 ;
      VIA 164.28 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 79.755 165.07 80.085 ;
      VIA 164.28 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 79.735 165.05 80.105 ;
      VIA 164.28 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 73.095 165.07 73.425 ;
      VIA 164.28 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 73.075 165.05 73.445 ;
      VIA 164.28 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 66.435 165.07 66.765 ;
      VIA 164.28 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 66.415 165.05 66.785 ;
      VIA 164.28 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 59.775 165.07 60.105 ;
      VIA 164.28 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 59.755 165.05 60.125 ;
      VIA 164.28 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 53.115 165.07 53.445 ;
      VIA 164.28 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 53.095 165.05 53.465 ;
      VIA 164.28 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 46.455 165.07 46.785 ;
      VIA 164.28 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 46.435 165.05 46.805 ;
      VIA 164.28 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 39.795 165.07 40.125 ;
      VIA 164.28 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 39.775 165.05 40.145 ;
      VIA 164.28 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 33.135 165.07 33.465 ;
      VIA 164.28 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 33.115 165.05 33.485 ;
      VIA 164.28 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 26.475 165.07 26.805 ;
      VIA 164.28 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 26.455 165.05 26.825 ;
      VIA 164.28 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 19.815 165.07 20.145 ;
      VIA 164.28 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 19.795 165.05 20.165 ;
      VIA 164.28 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 13.155 165.07 13.485 ;
      VIA 164.28 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 13.135 165.05 13.505 ;
      VIA 164.28 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.49 6.495 165.07 6.825 ;
      VIA 164.28 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.51 6.475 165.05 6.845 ;
      VIA 164.28 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 164.28 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 779.055 137.93 779.385 ;
      VIA 137.14 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 779.035 137.91 779.405 ;
      VIA 137.14 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 772.395 137.93 772.725 ;
      VIA 137.14 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 772.375 137.91 772.745 ;
      VIA 137.14 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 765.735 137.93 766.065 ;
      VIA 137.14 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 765.715 137.91 766.085 ;
      VIA 137.14 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 759.075 137.93 759.405 ;
      VIA 137.14 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 759.055 137.91 759.425 ;
      VIA 137.14 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 752.415 137.93 752.745 ;
      VIA 137.14 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 752.395 137.91 752.765 ;
      VIA 137.14 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 745.755 137.93 746.085 ;
      VIA 137.14 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 745.735 137.91 746.105 ;
      VIA 137.14 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 739.095 137.93 739.425 ;
      VIA 137.14 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 739.075 137.91 739.445 ;
      VIA 137.14 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 732.435 137.93 732.765 ;
      VIA 137.14 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 732.415 137.91 732.785 ;
      VIA 137.14 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 725.775 137.93 726.105 ;
      VIA 137.14 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 725.755 137.91 726.125 ;
      VIA 137.14 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 719.115 137.93 719.445 ;
      VIA 137.14 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 719.095 137.91 719.465 ;
      VIA 137.14 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 712.455 137.93 712.785 ;
      VIA 137.14 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 712.435 137.91 712.805 ;
      VIA 137.14 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 705.795 137.93 706.125 ;
      VIA 137.14 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 705.775 137.91 706.145 ;
      VIA 137.14 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 699.135 137.93 699.465 ;
      VIA 137.14 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 699.115 137.91 699.485 ;
      VIA 137.14 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 692.475 137.93 692.805 ;
      VIA 137.14 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 692.455 137.91 692.825 ;
      VIA 137.14 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 685.815 137.93 686.145 ;
      VIA 137.14 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 685.795 137.91 686.165 ;
      VIA 137.14 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 679.155 137.93 679.485 ;
      VIA 137.14 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 679.135 137.91 679.505 ;
      VIA 137.14 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 672.495 137.93 672.825 ;
      VIA 137.14 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 672.475 137.91 672.845 ;
      VIA 137.14 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 665.835 137.93 666.165 ;
      VIA 137.14 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 665.815 137.91 666.185 ;
      VIA 137.14 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 659.175 137.93 659.505 ;
      VIA 137.14 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 659.155 137.91 659.525 ;
      VIA 137.14 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 652.515 137.93 652.845 ;
      VIA 137.14 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 652.495 137.91 652.865 ;
      VIA 137.14 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 645.855 137.93 646.185 ;
      VIA 137.14 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 645.835 137.91 646.205 ;
      VIA 137.14 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 639.195 137.93 639.525 ;
      VIA 137.14 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 639.175 137.91 639.545 ;
      VIA 137.14 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 632.535 137.93 632.865 ;
      VIA 137.14 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 632.515 137.91 632.885 ;
      VIA 137.14 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 625.875 137.93 626.205 ;
      VIA 137.14 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 625.855 137.91 626.225 ;
      VIA 137.14 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 619.215 137.93 619.545 ;
      VIA 137.14 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 619.195 137.91 619.565 ;
      VIA 137.14 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 612.555 137.93 612.885 ;
      VIA 137.14 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 612.535 137.91 612.905 ;
      VIA 137.14 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 605.895 137.93 606.225 ;
      VIA 137.14 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 605.875 137.91 606.245 ;
      VIA 137.14 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 599.235 137.93 599.565 ;
      VIA 137.14 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 599.215 137.91 599.585 ;
      VIA 137.14 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 592.575 137.93 592.905 ;
      VIA 137.14 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 592.555 137.91 592.925 ;
      VIA 137.14 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 585.915 137.93 586.245 ;
      VIA 137.14 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 585.895 137.91 586.265 ;
      VIA 137.14 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 579.255 137.93 579.585 ;
      VIA 137.14 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 579.235 137.91 579.605 ;
      VIA 137.14 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 572.595 137.93 572.925 ;
      VIA 137.14 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 572.575 137.91 572.945 ;
      VIA 137.14 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 565.935 137.93 566.265 ;
      VIA 137.14 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 565.915 137.91 566.285 ;
      VIA 137.14 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 559.275 137.93 559.605 ;
      VIA 137.14 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 559.255 137.91 559.625 ;
      VIA 137.14 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 552.615 137.93 552.945 ;
      VIA 137.14 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 552.595 137.91 552.965 ;
      VIA 137.14 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 545.955 137.93 546.285 ;
      VIA 137.14 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 545.935 137.91 546.305 ;
      VIA 137.14 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 539.295 137.93 539.625 ;
      VIA 137.14 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 539.275 137.91 539.645 ;
      VIA 137.14 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 532.635 137.93 532.965 ;
      VIA 137.14 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 532.615 137.91 532.985 ;
      VIA 137.14 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 525.975 137.93 526.305 ;
      VIA 137.14 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 525.955 137.91 526.325 ;
      VIA 137.14 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 519.315 137.93 519.645 ;
      VIA 137.14 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 519.295 137.91 519.665 ;
      VIA 137.14 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 512.655 137.93 512.985 ;
      VIA 137.14 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 512.635 137.91 513.005 ;
      VIA 137.14 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 505.995 137.93 506.325 ;
      VIA 137.14 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 505.975 137.91 506.345 ;
      VIA 137.14 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 499.335 137.93 499.665 ;
      VIA 137.14 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 499.315 137.91 499.685 ;
      VIA 137.14 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 492.675 137.93 493.005 ;
      VIA 137.14 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 492.655 137.91 493.025 ;
      VIA 137.14 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 486.015 137.93 486.345 ;
      VIA 137.14 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 485.995 137.91 486.365 ;
      VIA 137.14 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 479.355 137.93 479.685 ;
      VIA 137.14 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 479.335 137.91 479.705 ;
      VIA 137.14 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 472.695 137.93 473.025 ;
      VIA 137.14 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 472.675 137.91 473.045 ;
      VIA 137.14 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 466.035 137.93 466.365 ;
      VIA 137.14 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 466.015 137.91 466.385 ;
      VIA 137.14 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 459.375 137.93 459.705 ;
      VIA 137.14 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 459.355 137.91 459.725 ;
      VIA 137.14 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 452.715 137.93 453.045 ;
      VIA 137.14 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 452.695 137.91 453.065 ;
      VIA 137.14 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 446.055 137.93 446.385 ;
      VIA 137.14 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 446.035 137.91 446.405 ;
      VIA 137.14 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 439.395 137.93 439.725 ;
      VIA 137.14 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 439.375 137.91 439.745 ;
      VIA 137.14 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 432.735 137.93 433.065 ;
      VIA 137.14 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 432.715 137.91 433.085 ;
      VIA 137.14 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 426.075 137.93 426.405 ;
      VIA 137.14 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 426.055 137.91 426.425 ;
      VIA 137.14 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 419.415 137.93 419.745 ;
      VIA 137.14 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 419.395 137.91 419.765 ;
      VIA 137.14 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 412.755 137.93 413.085 ;
      VIA 137.14 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 412.735 137.91 413.105 ;
      VIA 137.14 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 406.095 137.93 406.425 ;
      VIA 137.14 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 406.075 137.91 406.445 ;
      VIA 137.14 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 399.435 137.93 399.765 ;
      VIA 137.14 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 399.415 137.91 399.785 ;
      VIA 137.14 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 392.775 137.93 393.105 ;
      VIA 137.14 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 392.755 137.91 393.125 ;
      VIA 137.14 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 386.115 137.93 386.445 ;
      VIA 137.14 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 386.095 137.91 386.465 ;
      VIA 137.14 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 379.455 137.93 379.785 ;
      VIA 137.14 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 379.435 137.91 379.805 ;
      VIA 137.14 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 372.795 137.93 373.125 ;
      VIA 137.14 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 372.775 137.91 373.145 ;
      VIA 137.14 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 366.135 137.93 366.465 ;
      VIA 137.14 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 366.115 137.91 366.485 ;
      VIA 137.14 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 359.475 137.93 359.805 ;
      VIA 137.14 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 359.455 137.91 359.825 ;
      VIA 137.14 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 352.815 137.93 353.145 ;
      VIA 137.14 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 352.795 137.91 353.165 ;
      VIA 137.14 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 346.155 137.93 346.485 ;
      VIA 137.14 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 346.135 137.91 346.505 ;
      VIA 137.14 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 339.495 137.93 339.825 ;
      VIA 137.14 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 339.475 137.91 339.845 ;
      VIA 137.14 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 332.835 137.93 333.165 ;
      VIA 137.14 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 332.815 137.91 333.185 ;
      VIA 137.14 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 326.175 137.93 326.505 ;
      VIA 137.14 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 326.155 137.91 326.525 ;
      VIA 137.14 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 319.515 137.93 319.845 ;
      VIA 137.14 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 319.495 137.91 319.865 ;
      VIA 137.14 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 312.855 137.93 313.185 ;
      VIA 137.14 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 312.835 137.91 313.205 ;
      VIA 137.14 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 306.195 137.93 306.525 ;
      VIA 137.14 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 306.175 137.91 306.545 ;
      VIA 137.14 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 299.535 137.93 299.865 ;
      VIA 137.14 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 299.515 137.91 299.885 ;
      VIA 137.14 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 292.875 137.93 293.205 ;
      VIA 137.14 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 292.855 137.91 293.225 ;
      VIA 137.14 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 286.215 137.93 286.545 ;
      VIA 137.14 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 286.195 137.91 286.565 ;
      VIA 137.14 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 279.555 137.93 279.885 ;
      VIA 137.14 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 279.535 137.91 279.905 ;
      VIA 137.14 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 272.895 137.93 273.225 ;
      VIA 137.14 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 272.875 137.91 273.245 ;
      VIA 137.14 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 266.235 137.93 266.565 ;
      VIA 137.14 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 266.215 137.91 266.585 ;
      VIA 137.14 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 259.575 137.93 259.905 ;
      VIA 137.14 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 259.555 137.91 259.925 ;
      VIA 137.14 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 252.915 137.93 253.245 ;
      VIA 137.14 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 252.895 137.91 253.265 ;
      VIA 137.14 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 246.255 137.93 246.585 ;
      VIA 137.14 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 246.235 137.91 246.605 ;
      VIA 137.14 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 239.595 137.93 239.925 ;
      VIA 137.14 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 239.575 137.91 239.945 ;
      VIA 137.14 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 232.935 137.93 233.265 ;
      VIA 137.14 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 232.915 137.91 233.285 ;
      VIA 137.14 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 226.275 137.93 226.605 ;
      VIA 137.14 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 226.255 137.91 226.625 ;
      VIA 137.14 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 219.615 137.93 219.945 ;
      VIA 137.14 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 219.595 137.91 219.965 ;
      VIA 137.14 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 212.955 137.93 213.285 ;
      VIA 137.14 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 212.935 137.91 213.305 ;
      VIA 137.14 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 206.295 137.93 206.625 ;
      VIA 137.14 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 206.275 137.91 206.645 ;
      VIA 137.14 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 199.635 137.93 199.965 ;
      VIA 137.14 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 199.615 137.91 199.985 ;
      VIA 137.14 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 192.975 137.93 193.305 ;
      VIA 137.14 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 192.955 137.91 193.325 ;
      VIA 137.14 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 186.315 137.93 186.645 ;
      VIA 137.14 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 186.295 137.91 186.665 ;
      VIA 137.14 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 179.655 137.93 179.985 ;
      VIA 137.14 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 179.635 137.91 180.005 ;
      VIA 137.14 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 172.995 137.93 173.325 ;
      VIA 137.14 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 172.975 137.91 173.345 ;
      VIA 137.14 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 166.335 137.93 166.665 ;
      VIA 137.14 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 166.315 137.91 166.685 ;
      VIA 137.14 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 159.675 137.93 160.005 ;
      VIA 137.14 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 159.655 137.91 160.025 ;
      VIA 137.14 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 153.015 137.93 153.345 ;
      VIA 137.14 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 152.995 137.91 153.365 ;
      VIA 137.14 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 146.355 137.93 146.685 ;
      VIA 137.14 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 146.335 137.91 146.705 ;
      VIA 137.14 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 139.695 137.93 140.025 ;
      VIA 137.14 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 139.675 137.91 140.045 ;
      VIA 137.14 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 133.035 137.93 133.365 ;
      VIA 137.14 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 133.015 137.91 133.385 ;
      VIA 137.14 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 126.375 137.93 126.705 ;
      VIA 137.14 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 126.355 137.91 126.725 ;
      VIA 137.14 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 119.715 137.93 120.045 ;
      VIA 137.14 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 119.695 137.91 120.065 ;
      VIA 137.14 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 113.055 137.93 113.385 ;
      VIA 137.14 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 113.035 137.91 113.405 ;
      VIA 137.14 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 106.395 137.93 106.725 ;
      VIA 137.14 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 106.375 137.91 106.745 ;
      VIA 137.14 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 99.735 137.93 100.065 ;
      VIA 137.14 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 99.715 137.91 100.085 ;
      VIA 137.14 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 93.075 137.93 93.405 ;
      VIA 137.14 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 93.055 137.91 93.425 ;
      VIA 137.14 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 86.415 137.93 86.745 ;
      VIA 137.14 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 86.395 137.91 86.765 ;
      VIA 137.14 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 79.755 137.93 80.085 ;
      VIA 137.14 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 79.735 137.91 80.105 ;
      VIA 137.14 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 73.095 137.93 73.425 ;
      VIA 137.14 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 73.075 137.91 73.445 ;
      VIA 137.14 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 66.435 137.93 66.765 ;
      VIA 137.14 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 66.415 137.91 66.785 ;
      VIA 137.14 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 59.775 137.93 60.105 ;
      VIA 137.14 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 59.755 137.91 60.125 ;
      VIA 137.14 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 53.115 137.93 53.445 ;
      VIA 137.14 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 53.095 137.91 53.465 ;
      VIA 137.14 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 46.455 137.93 46.785 ;
      VIA 137.14 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 46.435 137.91 46.805 ;
      VIA 137.14 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 39.795 137.93 40.125 ;
      VIA 137.14 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 39.775 137.91 40.145 ;
      VIA 137.14 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 33.135 137.93 33.465 ;
      VIA 137.14 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 33.115 137.91 33.485 ;
      VIA 137.14 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 26.475 137.93 26.805 ;
      VIA 137.14 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 26.455 137.91 26.825 ;
      VIA 137.14 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 19.815 137.93 20.145 ;
      VIA 137.14 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 19.795 137.91 20.165 ;
      VIA 137.14 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 13.155 137.93 13.485 ;
      VIA 137.14 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 13.135 137.91 13.505 ;
      VIA 137.14 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.35 6.495 137.93 6.825 ;
      VIA 137.14 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.37 6.475 137.91 6.845 ;
      VIA 137.14 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 137.14 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 779.055 110.79 779.385 ;
      VIA 110 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 779.035 110.77 779.405 ;
      VIA 110 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 772.395 110.79 772.725 ;
      VIA 110 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 772.375 110.77 772.745 ;
      VIA 110 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 765.735 110.79 766.065 ;
      VIA 110 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 765.715 110.77 766.085 ;
      VIA 110 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 759.075 110.79 759.405 ;
      VIA 110 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 759.055 110.77 759.425 ;
      VIA 110 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 752.415 110.79 752.745 ;
      VIA 110 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 752.395 110.77 752.765 ;
      VIA 110 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 745.755 110.79 746.085 ;
      VIA 110 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 745.735 110.77 746.105 ;
      VIA 110 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 739.095 110.79 739.425 ;
      VIA 110 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 739.075 110.77 739.445 ;
      VIA 110 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 732.435 110.79 732.765 ;
      VIA 110 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 732.415 110.77 732.785 ;
      VIA 110 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 725.775 110.79 726.105 ;
      VIA 110 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 725.755 110.77 726.125 ;
      VIA 110 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 719.115 110.79 719.445 ;
      VIA 110 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 719.095 110.77 719.465 ;
      VIA 110 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 712.455 110.79 712.785 ;
      VIA 110 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 712.435 110.77 712.805 ;
      VIA 110 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 705.795 110.79 706.125 ;
      VIA 110 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 705.775 110.77 706.145 ;
      VIA 110 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 699.135 110.79 699.465 ;
      VIA 110 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 699.115 110.77 699.485 ;
      VIA 110 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 692.475 110.79 692.805 ;
      VIA 110 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 692.455 110.77 692.825 ;
      VIA 110 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 685.815 110.79 686.145 ;
      VIA 110 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 685.795 110.77 686.165 ;
      VIA 110 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 679.155 110.79 679.485 ;
      VIA 110 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 679.135 110.77 679.505 ;
      VIA 110 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 672.495 110.79 672.825 ;
      VIA 110 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 672.475 110.77 672.845 ;
      VIA 110 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 665.835 110.79 666.165 ;
      VIA 110 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 665.815 110.77 666.185 ;
      VIA 110 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 659.175 110.79 659.505 ;
      VIA 110 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 659.155 110.77 659.525 ;
      VIA 110 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 652.515 110.79 652.845 ;
      VIA 110 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 652.495 110.77 652.865 ;
      VIA 110 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 645.855 110.79 646.185 ;
      VIA 110 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 645.835 110.77 646.205 ;
      VIA 110 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 639.195 110.79 639.525 ;
      VIA 110 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 639.175 110.77 639.545 ;
      VIA 110 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 632.535 110.79 632.865 ;
      VIA 110 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 632.515 110.77 632.885 ;
      VIA 110 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 625.875 110.79 626.205 ;
      VIA 110 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 625.855 110.77 626.225 ;
      VIA 110 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 619.215 110.79 619.545 ;
      VIA 110 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 619.195 110.77 619.565 ;
      VIA 110 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 612.555 110.79 612.885 ;
      VIA 110 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 612.535 110.77 612.905 ;
      VIA 110 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 605.895 110.79 606.225 ;
      VIA 110 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 605.875 110.77 606.245 ;
      VIA 110 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 599.235 110.79 599.565 ;
      VIA 110 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 599.215 110.77 599.585 ;
      VIA 110 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 592.575 110.79 592.905 ;
      VIA 110 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 592.555 110.77 592.925 ;
      VIA 110 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 585.915 110.79 586.245 ;
      VIA 110 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 585.895 110.77 586.265 ;
      VIA 110 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 579.255 110.79 579.585 ;
      VIA 110 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 579.235 110.77 579.605 ;
      VIA 110 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 572.595 110.79 572.925 ;
      VIA 110 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 572.575 110.77 572.945 ;
      VIA 110 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 565.935 110.79 566.265 ;
      VIA 110 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 565.915 110.77 566.285 ;
      VIA 110 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 559.275 110.79 559.605 ;
      VIA 110 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 559.255 110.77 559.625 ;
      VIA 110 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 552.615 110.79 552.945 ;
      VIA 110 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 552.595 110.77 552.965 ;
      VIA 110 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 545.955 110.79 546.285 ;
      VIA 110 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 545.935 110.77 546.305 ;
      VIA 110 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 539.295 110.79 539.625 ;
      VIA 110 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 539.275 110.77 539.645 ;
      VIA 110 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 532.635 110.79 532.965 ;
      VIA 110 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 532.615 110.77 532.985 ;
      VIA 110 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 525.975 110.79 526.305 ;
      VIA 110 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 525.955 110.77 526.325 ;
      VIA 110 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 519.315 110.79 519.645 ;
      VIA 110 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 519.295 110.77 519.665 ;
      VIA 110 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 512.655 110.79 512.985 ;
      VIA 110 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 512.635 110.77 513.005 ;
      VIA 110 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 505.995 110.79 506.325 ;
      VIA 110 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 505.975 110.77 506.345 ;
      VIA 110 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 499.335 110.79 499.665 ;
      VIA 110 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 499.315 110.77 499.685 ;
      VIA 110 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 492.675 110.79 493.005 ;
      VIA 110 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 492.655 110.77 493.025 ;
      VIA 110 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 486.015 110.79 486.345 ;
      VIA 110 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 485.995 110.77 486.365 ;
      VIA 110 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 479.355 110.79 479.685 ;
      VIA 110 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 479.335 110.77 479.705 ;
      VIA 110 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 472.695 110.79 473.025 ;
      VIA 110 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 472.675 110.77 473.045 ;
      VIA 110 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 466.035 110.79 466.365 ;
      VIA 110 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 466.015 110.77 466.385 ;
      VIA 110 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 459.375 110.79 459.705 ;
      VIA 110 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 459.355 110.77 459.725 ;
      VIA 110 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 452.715 110.79 453.045 ;
      VIA 110 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 452.695 110.77 453.065 ;
      VIA 110 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 446.055 110.79 446.385 ;
      VIA 110 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 446.035 110.77 446.405 ;
      VIA 110 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 439.395 110.79 439.725 ;
      VIA 110 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 439.375 110.77 439.745 ;
      VIA 110 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 432.735 110.79 433.065 ;
      VIA 110 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 432.715 110.77 433.085 ;
      VIA 110 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 426.075 110.79 426.405 ;
      VIA 110 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 426.055 110.77 426.425 ;
      VIA 110 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 419.415 110.79 419.745 ;
      VIA 110 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 419.395 110.77 419.765 ;
      VIA 110 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 412.755 110.79 413.085 ;
      VIA 110 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 412.735 110.77 413.105 ;
      VIA 110 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 406.095 110.79 406.425 ;
      VIA 110 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 406.075 110.77 406.445 ;
      VIA 110 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 399.435 110.79 399.765 ;
      VIA 110 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 399.415 110.77 399.785 ;
      VIA 110 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 392.775 110.79 393.105 ;
      VIA 110 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 392.755 110.77 393.125 ;
      VIA 110 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 386.115 110.79 386.445 ;
      VIA 110 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 386.095 110.77 386.465 ;
      VIA 110 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 379.455 110.79 379.785 ;
      VIA 110 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 379.435 110.77 379.805 ;
      VIA 110 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 372.795 110.79 373.125 ;
      VIA 110 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 372.775 110.77 373.145 ;
      VIA 110 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 366.135 110.79 366.465 ;
      VIA 110 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 366.115 110.77 366.485 ;
      VIA 110 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 359.475 110.79 359.805 ;
      VIA 110 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 359.455 110.77 359.825 ;
      VIA 110 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 352.815 110.79 353.145 ;
      VIA 110 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 352.795 110.77 353.165 ;
      VIA 110 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 346.155 110.79 346.485 ;
      VIA 110 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 346.135 110.77 346.505 ;
      VIA 110 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 339.495 110.79 339.825 ;
      VIA 110 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 339.475 110.77 339.845 ;
      VIA 110 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 332.835 110.79 333.165 ;
      VIA 110 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 332.815 110.77 333.185 ;
      VIA 110 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 326.175 110.79 326.505 ;
      VIA 110 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 326.155 110.77 326.525 ;
      VIA 110 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 319.515 110.79 319.845 ;
      VIA 110 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 319.495 110.77 319.865 ;
      VIA 110 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 312.855 110.79 313.185 ;
      VIA 110 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 312.835 110.77 313.205 ;
      VIA 110 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 306.195 110.79 306.525 ;
      VIA 110 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 306.175 110.77 306.545 ;
      VIA 110 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 299.535 110.79 299.865 ;
      VIA 110 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 299.515 110.77 299.885 ;
      VIA 110 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 292.875 110.79 293.205 ;
      VIA 110 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 292.855 110.77 293.225 ;
      VIA 110 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 286.215 110.79 286.545 ;
      VIA 110 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 286.195 110.77 286.565 ;
      VIA 110 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 279.555 110.79 279.885 ;
      VIA 110 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 279.535 110.77 279.905 ;
      VIA 110 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 272.895 110.79 273.225 ;
      VIA 110 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 272.875 110.77 273.245 ;
      VIA 110 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 266.235 110.79 266.565 ;
      VIA 110 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 266.215 110.77 266.585 ;
      VIA 110 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 259.575 110.79 259.905 ;
      VIA 110 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 259.555 110.77 259.925 ;
      VIA 110 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 252.915 110.79 253.245 ;
      VIA 110 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 252.895 110.77 253.265 ;
      VIA 110 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 246.255 110.79 246.585 ;
      VIA 110 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 246.235 110.77 246.605 ;
      VIA 110 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 239.595 110.79 239.925 ;
      VIA 110 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 239.575 110.77 239.945 ;
      VIA 110 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 232.935 110.79 233.265 ;
      VIA 110 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 232.915 110.77 233.285 ;
      VIA 110 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 226.275 110.79 226.605 ;
      VIA 110 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 226.255 110.77 226.625 ;
      VIA 110 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 219.615 110.79 219.945 ;
      VIA 110 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 219.595 110.77 219.965 ;
      VIA 110 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 212.955 110.79 213.285 ;
      VIA 110 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 212.935 110.77 213.305 ;
      VIA 110 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 206.295 110.79 206.625 ;
      VIA 110 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 206.275 110.77 206.645 ;
      VIA 110 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 199.635 110.79 199.965 ;
      VIA 110 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 199.615 110.77 199.985 ;
      VIA 110 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 192.975 110.79 193.305 ;
      VIA 110 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 192.955 110.77 193.325 ;
      VIA 110 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 186.315 110.79 186.645 ;
      VIA 110 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 186.295 110.77 186.665 ;
      VIA 110 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 179.655 110.79 179.985 ;
      VIA 110 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 179.635 110.77 180.005 ;
      VIA 110 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 172.995 110.79 173.325 ;
      VIA 110 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 172.975 110.77 173.345 ;
      VIA 110 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 166.335 110.79 166.665 ;
      VIA 110 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 166.315 110.77 166.685 ;
      VIA 110 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 159.675 110.79 160.005 ;
      VIA 110 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 159.655 110.77 160.025 ;
      VIA 110 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 153.015 110.79 153.345 ;
      VIA 110 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 152.995 110.77 153.365 ;
      VIA 110 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 146.355 110.79 146.685 ;
      VIA 110 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 146.335 110.77 146.705 ;
      VIA 110 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 139.695 110.79 140.025 ;
      VIA 110 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 139.675 110.77 140.045 ;
      VIA 110 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 133.035 110.79 133.365 ;
      VIA 110 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 133.015 110.77 133.385 ;
      VIA 110 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 126.375 110.79 126.705 ;
      VIA 110 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 126.355 110.77 126.725 ;
      VIA 110 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 119.715 110.79 120.045 ;
      VIA 110 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 119.695 110.77 120.065 ;
      VIA 110 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 113.055 110.79 113.385 ;
      VIA 110 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 113.035 110.77 113.405 ;
      VIA 110 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 106.395 110.79 106.725 ;
      VIA 110 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 106.375 110.77 106.745 ;
      VIA 110 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 99.735 110.79 100.065 ;
      VIA 110 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 99.715 110.77 100.085 ;
      VIA 110 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 93.075 110.79 93.405 ;
      VIA 110 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 93.055 110.77 93.425 ;
      VIA 110 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 86.415 110.79 86.745 ;
      VIA 110 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 86.395 110.77 86.765 ;
      VIA 110 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 79.755 110.79 80.085 ;
      VIA 110 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 79.735 110.77 80.105 ;
      VIA 110 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 73.095 110.79 73.425 ;
      VIA 110 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 73.075 110.77 73.445 ;
      VIA 110 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 66.435 110.79 66.765 ;
      VIA 110 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 66.415 110.77 66.785 ;
      VIA 110 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 59.775 110.79 60.105 ;
      VIA 110 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 59.755 110.77 60.125 ;
      VIA 110 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 53.115 110.79 53.445 ;
      VIA 110 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 53.095 110.77 53.465 ;
      VIA 110 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 46.455 110.79 46.785 ;
      VIA 110 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 46.435 110.77 46.805 ;
      VIA 110 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 39.795 110.79 40.125 ;
      VIA 110 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 39.775 110.77 40.145 ;
      VIA 110 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 33.135 110.79 33.465 ;
      VIA 110 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 33.115 110.77 33.485 ;
      VIA 110 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 26.475 110.79 26.805 ;
      VIA 110 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 26.455 110.77 26.825 ;
      VIA 110 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 19.815 110.79 20.145 ;
      VIA 110 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 19.795 110.77 20.165 ;
      VIA 110 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 13.155 110.79 13.485 ;
      VIA 110 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 13.135 110.77 13.505 ;
      VIA 110 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.21 6.495 110.79 6.825 ;
      VIA 110 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.23 6.475 110.77 6.845 ;
      VIA 110 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 110 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 779.055 83.65 779.385 ;
      VIA 82.86 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 779.035 83.63 779.405 ;
      VIA 82.86 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 772.395 83.65 772.725 ;
      VIA 82.86 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 772.375 83.63 772.745 ;
      VIA 82.86 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 765.735 83.65 766.065 ;
      VIA 82.86 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 765.715 83.63 766.085 ;
      VIA 82.86 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 759.075 83.65 759.405 ;
      VIA 82.86 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 759.055 83.63 759.425 ;
      VIA 82.86 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 752.415 83.65 752.745 ;
      VIA 82.86 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 752.395 83.63 752.765 ;
      VIA 82.86 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 745.755 83.65 746.085 ;
      VIA 82.86 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 745.735 83.63 746.105 ;
      VIA 82.86 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 739.095 83.65 739.425 ;
      VIA 82.86 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 739.075 83.63 739.445 ;
      VIA 82.86 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 732.435 83.65 732.765 ;
      VIA 82.86 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 732.415 83.63 732.785 ;
      VIA 82.86 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 725.775 83.65 726.105 ;
      VIA 82.86 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 725.755 83.63 726.125 ;
      VIA 82.86 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 719.115 83.65 719.445 ;
      VIA 82.86 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 719.095 83.63 719.465 ;
      VIA 82.86 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 712.455 83.65 712.785 ;
      VIA 82.86 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 712.435 83.63 712.805 ;
      VIA 82.86 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 705.795 83.65 706.125 ;
      VIA 82.86 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 705.775 83.63 706.145 ;
      VIA 82.86 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 699.135 83.65 699.465 ;
      VIA 82.86 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 699.115 83.63 699.485 ;
      VIA 82.86 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 692.475 83.65 692.805 ;
      VIA 82.86 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 692.455 83.63 692.825 ;
      VIA 82.86 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 685.815 83.65 686.145 ;
      VIA 82.86 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 685.795 83.63 686.165 ;
      VIA 82.86 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 679.155 83.65 679.485 ;
      VIA 82.86 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 679.135 83.63 679.505 ;
      VIA 82.86 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 672.495 83.65 672.825 ;
      VIA 82.86 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 672.475 83.63 672.845 ;
      VIA 82.86 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 665.835 83.65 666.165 ;
      VIA 82.86 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 665.815 83.63 666.185 ;
      VIA 82.86 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 659.175 83.65 659.505 ;
      VIA 82.86 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 659.155 83.63 659.525 ;
      VIA 82.86 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 652.515 83.65 652.845 ;
      VIA 82.86 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 652.495 83.63 652.865 ;
      VIA 82.86 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 645.855 83.65 646.185 ;
      VIA 82.86 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 645.835 83.63 646.205 ;
      VIA 82.86 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 639.195 83.65 639.525 ;
      VIA 82.86 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 639.175 83.63 639.545 ;
      VIA 82.86 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 632.535 83.65 632.865 ;
      VIA 82.86 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 632.515 83.63 632.885 ;
      VIA 82.86 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 625.875 83.65 626.205 ;
      VIA 82.86 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 625.855 83.63 626.225 ;
      VIA 82.86 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 619.215 83.65 619.545 ;
      VIA 82.86 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 619.195 83.63 619.565 ;
      VIA 82.86 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 612.555 83.65 612.885 ;
      VIA 82.86 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 612.535 83.63 612.905 ;
      VIA 82.86 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 605.895 83.65 606.225 ;
      VIA 82.86 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 605.875 83.63 606.245 ;
      VIA 82.86 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 599.235 83.65 599.565 ;
      VIA 82.86 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 599.215 83.63 599.585 ;
      VIA 82.86 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 592.575 83.65 592.905 ;
      VIA 82.86 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 592.555 83.63 592.925 ;
      VIA 82.86 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 585.915 83.65 586.245 ;
      VIA 82.86 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 585.895 83.63 586.265 ;
      VIA 82.86 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 579.255 83.65 579.585 ;
      VIA 82.86 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 579.235 83.63 579.605 ;
      VIA 82.86 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 572.595 83.65 572.925 ;
      VIA 82.86 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 572.575 83.63 572.945 ;
      VIA 82.86 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 565.935 83.65 566.265 ;
      VIA 82.86 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 565.915 83.63 566.285 ;
      VIA 82.86 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 559.275 83.65 559.605 ;
      VIA 82.86 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 559.255 83.63 559.625 ;
      VIA 82.86 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 552.615 83.65 552.945 ;
      VIA 82.86 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 552.595 83.63 552.965 ;
      VIA 82.86 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 545.955 83.65 546.285 ;
      VIA 82.86 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 545.935 83.63 546.305 ;
      VIA 82.86 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 539.295 83.65 539.625 ;
      VIA 82.86 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 539.275 83.63 539.645 ;
      VIA 82.86 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 532.635 83.65 532.965 ;
      VIA 82.86 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 532.615 83.63 532.985 ;
      VIA 82.86 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 525.975 83.65 526.305 ;
      VIA 82.86 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 525.955 83.63 526.325 ;
      VIA 82.86 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 519.315 83.65 519.645 ;
      VIA 82.86 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 519.295 83.63 519.665 ;
      VIA 82.86 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 512.655 83.65 512.985 ;
      VIA 82.86 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 512.635 83.63 513.005 ;
      VIA 82.86 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 505.995 83.65 506.325 ;
      VIA 82.86 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 505.975 83.63 506.345 ;
      VIA 82.86 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 499.335 83.65 499.665 ;
      VIA 82.86 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 499.315 83.63 499.685 ;
      VIA 82.86 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 492.675 83.65 493.005 ;
      VIA 82.86 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 492.655 83.63 493.025 ;
      VIA 82.86 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 486.015 83.65 486.345 ;
      VIA 82.86 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 485.995 83.63 486.365 ;
      VIA 82.86 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 479.355 83.65 479.685 ;
      VIA 82.86 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 479.335 83.63 479.705 ;
      VIA 82.86 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 472.695 83.65 473.025 ;
      VIA 82.86 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 472.675 83.63 473.045 ;
      VIA 82.86 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 466.035 83.65 466.365 ;
      VIA 82.86 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 466.015 83.63 466.385 ;
      VIA 82.86 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 459.375 83.65 459.705 ;
      VIA 82.86 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 459.355 83.63 459.725 ;
      VIA 82.86 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 452.715 83.65 453.045 ;
      VIA 82.86 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 452.695 83.63 453.065 ;
      VIA 82.86 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 446.055 83.65 446.385 ;
      VIA 82.86 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 446.035 83.63 446.405 ;
      VIA 82.86 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 439.395 83.65 439.725 ;
      VIA 82.86 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 439.375 83.63 439.745 ;
      VIA 82.86 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 432.735 83.65 433.065 ;
      VIA 82.86 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 432.715 83.63 433.085 ;
      VIA 82.86 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 426.075 83.65 426.405 ;
      VIA 82.86 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 426.055 83.63 426.425 ;
      VIA 82.86 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 419.415 83.65 419.745 ;
      VIA 82.86 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 419.395 83.63 419.765 ;
      VIA 82.86 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 412.755 83.65 413.085 ;
      VIA 82.86 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 412.735 83.63 413.105 ;
      VIA 82.86 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 406.095 83.65 406.425 ;
      VIA 82.86 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 406.075 83.63 406.445 ;
      VIA 82.86 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 399.435 83.65 399.765 ;
      VIA 82.86 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 399.415 83.63 399.785 ;
      VIA 82.86 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 392.775 83.65 393.105 ;
      VIA 82.86 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 392.755 83.63 393.125 ;
      VIA 82.86 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 386.115 83.65 386.445 ;
      VIA 82.86 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 386.095 83.63 386.465 ;
      VIA 82.86 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 379.455 83.65 379.785 ;
      VIA 82.86 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 379.435 83.63 379.805 ;
      VIA 82.86 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 372.795 83.65 373.125 ;
      VIA 82.86 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 372.775 83.63 373.145 ;
      VIA 82.86 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 366.135 83.65 366.465 ;
      VIA 82.86 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 366.115 83.63 366.485 ;
      VIA 82.86 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 359.475 83.65 359.805 ;
      VIA 82.86 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 359.455 83.63 359.825 ;
      VIA 82.86 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 352.815 83.65 353.145 ;
      VIA 82.86 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 352.795 83.63 353.165 ;
      VIA 82.86 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 346.155 83.65 346.485 ;
      VIA 82.86 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 346.135 83.63 346.505 ;
      VIA 82.86 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 339.495 83.65 339.825 ;
      VIA 82.86 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 339.475 83.63 339.845 ;
      VIA 82.86 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 332.835 83.65 333.165 ;
      VIA 82.86 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 332.815 83.63 333.185 ;
      VIA 82.86 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 326.175 83.65 326.505 ;
      VIA 82.86 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 326.155 83.63 326.525 ;
      VIA 82.86 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 319.515 83.65 319.845 ;
      VIA 82.86 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 319.495 83.63 319.865 ;
      VIA 82.86 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 312.855 83.65 313.185 ;
      VIA 82.86 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 312.835 83.63 313.205 ;
      VIA 82.86 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 306.195 83.65 306.525 ;
      VIA 82.86 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 306.175 83.63 306.545 ;
      VIA 82.86 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 299.535 83.65 299.865 ;
      VIA 82.86 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 299.515 83.63 299.885 ;
      VIA 82.86 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 292.875 83.65 293.205 ;
      VIA 82.86 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 292.855 83.63 293.225 ;
      VIA 82.86 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 286.215 83.65 286.545 ;
      VIA 82.86 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 286.195 83.63 286.565 ;
      VIA 82.86 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 279.555 83.65 279.885 ;
      VIA 82.86 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 279.535 83.63 279.905 ;
      VIA 82.86 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 272.895 83.65 273.225 ;
      VIA 82.86 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 272.875 83.63 273.245 ;
      VIA 82.86 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 266.235 83.65 266.565 ;
      VIA 82.86 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 266.215 83.63 266.585 ;
      VIA 82.86 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 259.575 83.65 259.905 ;
      VIA 82.86 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 259.555 83.63 259.925 ;
      VIA 82.86 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 252.915 83.65 253.245 ;
      VIA 82.86 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 252.895 83.63 253.265 ;
      VIA 82.86 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 246.255 83.65 246.585 ;
      VIA 82.86 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 246.235 83.63 246.605 ;
      VIA 82.86 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 239.595 83.65 239.925 ;
      VIA 82.86 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 239.575 83.63 239.945 ;
      VIA 82.86 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 232.935 83.65 233.265 ;
      VIA 82.86 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 232.915 83.63 233.285 ;
      VIA 82.86 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 226.275 83.65 226.605 ;
      VIA 82.86 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 226.255 83.63 226.625 ;
      VIA 82.86 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 219.615 83.65 219.945 ;
      VIA 82.86 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 219.595 83.63 219.965 ;
      VIA 82.86 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 212.955 83.65 213.285 ;
      VIA 82.86 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 212.935 83.63 213.305 ;
      VIA 82.86 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 206.295 83.65 206.625 ;
      VIA 82.86 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 206.275 83.63 206.645 ;
      VIA 82.86 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 199.635 83.65 199.965 ;
      VIA 82.86 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 199.615 83.63 199.985 ;
      VIA 82.86 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 192.975 83.65 193.305 ;
      VIA 82.86 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 192.955 83.63 193.325 ;
      VIA 82.86 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 186.315 83.65 186.645 ;
      VIA 82.86 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 186.295 83.63 186.665 ;
      VIA 82.86 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 179.655 83.65 179.985 ;
      VIA 82.86 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 179.635 83.63 180.005 ;
      VIA 82.86 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 172.995 83.65 173.325 ;
      VIA 82.86 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 172.975 83.63 173.345 ;
      VIA 82.86 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 166.335 83.65 166.665 ;
      VIA 82.86 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 166.315 83.63 166.685 ;
      VIA 82.86 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 159.675 83.65 160.005 ;
      VIA 82.86 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 159.655 83.63 160.025 ;
      VIA 82.86 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 153.015 83.65 153.345 ;
      VIA 82.86 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 152.995 83.63 153.365 ;
      VIA 82.86 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 146.355 83.65 146.685 ;
      VIA 82.86 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 146.335 83.63 146.705 ;
      VIA 82.86 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 139.695 83.65 140.025 ;
      VIA 82.86 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 139.675 83.63 140.045 ;
      VIA 82.86 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 133.035 83.65 133.365 ;
      VIA 82.86 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 133.015 83.63 133.385 ;
      VIA 82.86 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 126.375 83.65 126.705 ;
      VIA 82.86 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 126.355 83.63 126.725 ;
      VIA 82.86 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 119.715 83.65 120.045 ;
      VIA 82.86 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 119.695 83.63 120.065 ;
      VIA 82.86 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 113.055 83.65 113.385 ;
      VIA 82.86 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 113.035 83.63 113.405 ;
      VIA 82.86 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 106.395 83.65 106.725 ;
      VIA 82.86 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 106.375 83.63 106.745 ;
      VIA 82.86 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 99.735 83.65 100.065 ;
      VIA 82.86 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 99.715 83.63 100.085 ;
      VIA 82.86 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 93.075 83.65 93.405 ;
      VIA 82.86 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 93.055 83.63 93.425 ;
      VIA 82.86 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 86.415 83.65 86.745 ;
      VIA 82.86 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 86.395 83.63 86.765 ;
      VIA 82.86 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 79.755 83.65 80.085 ;
      VIA 82.86 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 79.735 83.63 80.105 ;
      VIA 82.86 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 73.095 83.65 73.425 ;
      VIA 82.86 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 73.075 83.63 73.445 ;
      VIA 82.86 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 66.435 83.65 66.765 ;
      VIA 82.86 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 66.415 83.63 66.785 ;
      VIA 82.86 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 59.775 83.65 60.105 ;
      VIA 82.86 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 59.755 83.63 60.125 ;
      VIA 82.86 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 53.115 83.65 53.445 ;
      VIA 82.86 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 53.095 83.63 53.465 ;
      VIA 82.86 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 46.455 83.65 46.785 ;
      VIA 82.86 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 46.435 83.63 46.805 ;
      VIA 82.86 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 39.795 83.65 40.125 ;
      VIA 82.86 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 39.775 83.63 40.145 ;
      VIA 82.86 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 33.135 83.65 33.465 ;
      VIA 82.86 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 33.115 83.63 33.485 ;
      VIA 82.86 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 26.475 83.65 26.805 ;
      VIA 82.86 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 26.455 83.63 26.825 ;
      VIA 82.86 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 19.815 83.65 20.145 ;
      VIA 82.86 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 19.795 83.63 20.165 ;
      VIA 82.86 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 13.155 83.65 13.485 ;
      VIA 82.86 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 13.135 83.63 13.505 ;
      VIA 82.86 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.07 6.495 83.65 6.825 ;
      VIA 82.86 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.09 6.475 83.63 6.845 ;
      VIA 82.86 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 82.86 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 779.055 56.51 779.385 ;
      VIA 55.72 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 779.035 56.49 779.405 ;
      VIA 55.72 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 772.395 56.51 772.725 ;
      VIA 55.72 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 772.375 56.49 772.745 ;
      VIA 55.72 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 765.735 56.51 766.065 ;
      VIA 55.72 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 765.715 56.49 766.085 ;
      VIA 55.72 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 759.075 56.51 759.405 ;
      VIA 55.72 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 759.055 56.49 759.425 ;
      VIA 55.72 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 752.415 56.51 752.745 ;
      VIA 55.72 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 752.395 56.49 752.765 ;
      VIA 55.72 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 745.755 56.51 746.085 ;
      VIA 55.72 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 745.735 56.49 746.105 ;
      VIA 55.72 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 739.095 56.51 739.425 ;
      VIA 55.72 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 739.075 56.49 739.445 ;
      VIA 55.72 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 732.435 56.51 732.765 ;
      VIA 55.72 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 732.415 56.49 732.785 ;
      VIA 55.72 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 725.775 56.51 726.105 ;
      VIA 55.72 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 725.755 56.49 726.125 ;
      VIA 55.72 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 719.115 56.51 719.445 ;
      VIA 55.72 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 719.095 56.49 719.465 ;
      VIA 55.72 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 712.455 56.51 712.785 ;
      VIA 55.72 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 712.435 56.49 712.805 ;
      VIA 55.72 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 705.795 56.51 706.125 ;
      VIA 55.72 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 705.775 56.49 706.145 ;
      VIA 55.72 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 699.135 56.51 699.465 ;
      VIA 55.72 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 699.115 56.49 699.485 ;
      VIA 55.72 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 692.475 56.51 692.805 ;
      VIA 55.72 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 692.455 56.49 692.825 ;
      VIA 55.72 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 685.815 56.51 686.145 ;
      VIA 55.72 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 685.795 56.49 686.165 ;
      VIA 55.72 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 679.155 56.51 679.485 ;
      VIA 55.72 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 679.135 56.49 679.505 ;
      VIA 55.72 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 672.495 56.51 672.825 ;
      VIA 55.72 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 672.475 56.49 672.845 ;
      VIA 55.72 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 665.835 56.51 666.165 ;
      VIA 55.72 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 665.815 56.49 666.185 ;
      VIA 55.72 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 659.175 56.51 659.505 ;
      VIA 55.72 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 659.155 56.49 659.525 ;
      VIA 55.72 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 652.515 56.51 652.845 ;
      VIA 55.72 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 652.495 56.49 652.865 ;
      VIA 55.72 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 645.855 56.51 646.185 ;
      VIA 55.72 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 645.835 56.49 646.205 ;
      VIA 55.72 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 639.195 56.51 639.525 ;
      VIA 55.72 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 639.175 56.49 639.545 ;
      VIA 55.72 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 632.535 56.51 632.865 ;
      VIA 55.72 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 632.515 56.49 632.885 ;
      VIA 55.72 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 625.875 56.51 626.205 ;
      VIA 55.72 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 625.855 56.49 626.225 ;
      VIA 55.72 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 619.215 56.51 619.545 ;
      VIA 55.72 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 619.195 56.49 619.565 ;
      VIA 55.72 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 612.555 56.51 612.885 ;
      VIA 55.72 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 612.535 56.49 612.905 ;
      VIA 55.72 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 605.895 56.51 606.225 ;
      VIA 55.72 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 605.875 56.49 606.245 ;
      VIA 55.72 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 599.235 56.51 599.565 ;
      VIA 55.72 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 599.215 56.49 599.585 ;
      VIA 55.72 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 592.575 56.51 592.905 ;
      VIA 55.72 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 592.555 56.49 592.925 ;
      VIA 55.72 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 585.915 56.51 586.245 ;
      VIA 55.72 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 585.895 56.49 586.265 ;
      VIA 55.72 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 579.255 56.51 579.585 ;
      VIA 55.72 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 579.235 56.49 579.605 ;
      VIA 55.72 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 572.595 56.51 572.925 ;
      VIA 55.72 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 572.575 56.49 572.945 ;
      VIA 55.72 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 565.935 56.51 566.265 ;
      VIA 55.72 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 565.915 56.49 566.285 ;
      VIA 55.72 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 559.275 56.51 559.605 ;
      VIA 55.72 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 559.255 56.49 559.625 ;
      VIA 55.72 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 552.615 56.51 552.945 ;
      VIA 55.72 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 552.595 56.49 552.965 ;
      VIA 55.72 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 545.955 56.51 546.285 ;
      VIA 55.72 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 545.935 56.49 546.305 ;
      VIA 55.72 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 539.295 56.51 539.625 ;
      VIA 55.72 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 539.275 56.49 539.645 ;
      VIA 55.72 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 532.635 56.51 532.965 ;
      VIA 55.72 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 532.615 56.49 532.985 ;
      VIA 55.72 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 525.975 56.51 526.305 ;
      VIA 55.72 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 525.955 56.49 526.325 ;
      VIA 55.72 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 519.315 56.51 519.645 ;
      VIA 55.72 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 519.295 56.49 519.665 ;
      VIA 55.72 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 512.655 56.51 512.985 ;
      VIA 55.72 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 512.635 56.49 513.005 ;
      VIA 55.72 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 505.995 56.51 506.325 ;
      VIA 55.72 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 505.975 56.49 506.345 ;
      VIA 55.72 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 499.335 56.51 499.665 ;
      VIA 55.72 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 499.315 56.49 499.685 ;
      VIA 55.72 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 492.675 56.51 493.005 ;
      VIA 55.72 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 492.655 56.49 493.025 ;
      VIA 55.72 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 486.015 56.51 486.345 ;
      VIA 55.72 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 485.995 56.49 486.365 ;
      VIA 55.72 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 479.355 56.51 479.685 ;
      VIA 55.72 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 479.335 56.49 479.705 ;
      VIA 55.72 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 472.695 56.51 473.025 ;
      VIA 55.72 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 472.675 56.49 473.045 ;
      VIA 55.72 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 466.035 56.51 466.365 ;
      VIA 55.72 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 466.015 56.49 466.385 ;
      VIA 55.72 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 459.375 56.51 459.705 ;
      VIA 55.72 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 459.355 56.49 459.725 ;
      VIA 55.72 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 452.715 56.51 453.045 ;
      VIA 55.72 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 452.695 56.49 453.065 ;
      VIA 55.72 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 446.055 56.51 446.385 ;
      VIA 55.72 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 446.035 56.49 446.405 ;
      VIA 55.72 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 439.395 56.51 439.725 ;
      VIA 55.72 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 439.375 56.49 439.745 ;
      VIA 55.72 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 432.735 56.51 433.065 ;
      VIA 55.72 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 432.715 56.49 433.085 ;
      VIA 55.72 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 426.075 56.51 426.405 ;
      VIA 55.72 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 426.055 56.49 426.425 ;
      VIA 55.72 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 419.415 56.51 419.745 ;
      VIA 55.72 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 419.395 56.49 419.765 ;
      VIA 55.72 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 412.755 56.51 413.085 ;
      VIA 55.72 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 412.735 56.49 413.105 ;
      VIA 55.72 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 406.095 56.51 406.425 ;
      VIA 55.72 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 406.075 56.49 406.445 ;
      VIA 55.72 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 399.435 56.51 399.765 ;
      VIA 55.72 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 399.415 56.49 399.785 ;
      VIA 55.72 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 392.775 56.51 393.105 ;
      VIA 55.72 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 392.755 56.49 393.125 ;
      VIA 55.72 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 386.115 56.51 386.445 ;
      VIA 55.72 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 386.095 56.49 386.465 ;
      VIA 55.72 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 379.455 56.51 379.785 ;
      VIA 55.72 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 379.435 56.49 379.805 ;
      VIA 55.72 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 372.795 56.51 373.125 ;
      VIA 55.72 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 372.775 56.49 373.145 ;
      VIA 55.72 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 366.135 56.51 366.465 ;
      VIA 55.72 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 366.115 56.49 366.485 ;
      VIA 55.72 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 359.475 56.51 359.805 ;
      VIA 55.72 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 359.455 56.49 359.825 ;
      VIA 55.72 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 352.815 56.51 353.145 ;
      VIA 55.72 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 352.795 56.49 353.165 ;
      VIA 55.72 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 346.155 56.51 346.485 ;
      VIA 55.72 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 346.135 56.49 346.505 ;
      VIA 55.72 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 339.495 56.51 339.825 ;
      VIA 55.72 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 339.475 56.49 339.845 ;
      VIA 55.72 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 332.835 56.51 333.165 ;
      VIA 55.72 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 332.815 56.49 333.185 ;
      VIA 55.72 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 326.175 56.51 326.505 ;
      VIA 55.72 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 326.155 56.49 326.525 ;
      VIA 55.72 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 319.515 56.51 319.845 ;
      VIA 55.72 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 319.495 56.49 319.865 ;
      VIA 55.72 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 312.855 56.51 313.185 ;
      VIA 55.72 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 312.835 56.49 313.205 ;
      VIA 55.72 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 306.195 56.51 306.525 ;
      VIA 55.72 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 306.175 56.49 306.545 ;
      VIA 55.72 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 299.535 56.51 299.865 ;
      VIA 55.72 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 299.515 56.49 299.885 ;
      VIA 55.72 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 292.875 56.51 293.205 ;
      VIA 55.72 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 292.855 56.49 293.225 ;
      VIA 55.72 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 286.215 56.51 286.545 ;
      VIA 55.72 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 286.195 56.49 286.565 ;
      VIA 55.72 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 279.555 56.51 279.885 ;
      VIA 55.72 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 279.535 56.49 279.905 ;
      VIA 55.72 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 272.895 56.51 273.225 ;
      VIA 55.72 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 272.875 56.49 273.245 ;
      VIA 55.72 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 266.235 56.51 266.565 ;
      VIA 55.72 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 266.215 56.49 266.585 ;
      VIA 55.72 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 259.575 56.51 259.905 ;
      VIA 55.72 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 259.555 56.49 259.925 ;
      VIA 55.72 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 252.915 56.51 253.245 ;
      VIA 55.72 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 252.895 56.49 253.265 ;
      VIA 55.72 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 246.255 56.51 246.585 ;
      VIA 55.72 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 246.235 56.49 246.605 ;
      VIA 55.72 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 239.595 56.51 239.925 ;
      VIA 55.72 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 239.575 56.49 239.945 ;
      VIA 55.72 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 232.935 56.51 233.265 ;
      VIA 55.72 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 232.915 56.49 233.285 ;
      VIA 55.72 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 226.275 56.51 226.605 ;
      VIA 55.72 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 226.255 56.49 226.625 ;
      VIA 55.72 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 219.615 56.51 219.945 ;
      VIA 55.72 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 219.595 56.49 219.965 ;
      VIA 55.72 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 212.955 56.51 213.285 ;
      VIA 55.72 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 212.935 56.49 213.305 ;
      VIA 55.72 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 206.295 56.51 206.625 ;
      VIA 55.72 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 206.275 56.49 206.645 ;
      VIA 55.72 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 199.635 56.51 199.965 ;
      VIA 55.72 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 199.615 56.49 199.985 ;
      VIA 55.72 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 192.975 56.51 193.305 ;
      VIA 55.72 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 192.955 56.49 193.325 ;
      VIA 55.72 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 186.315 56.51 186.645 ;
      VIA 55.72 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 186.295 56.49 186.665 ;
      VIA 55.72 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 179.655 56.51 179.985 ;
      VIA 55.72 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 179.635 56.49 180.005 ;
      VIA 55.72 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 172.995 56.51 173.325 ;
      VIA 55.72 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 172.975 56.49 173.345 ;
      VIA 55.72 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 166.335 56.51 166.665 ;
      VIA 55.72 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 166.315 56.49 166.685 ;
      VIA 55.72 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 159.675 56.51 160.005 ;
      VIA 55.72 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 159.655 56.49 160.025 ;
      VIA 55.72 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 153.015 56.51 153.345 ;
      VIA 55.72 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 152.995 56.49 153.365 ;
      VIA 55.72 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 146.355 56.51 146.685 ;
      VIA 55.72 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 146.335 56.49 146.705 ;
      VIA 55.72 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 139.695 56.51 140.025 ;
      VIA 55.72 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 139.675 56.49 140.045 ;
      VIA 55.72 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 133.035 56.51 133.365 ;
      VIA 55.72 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 133.015 56.49 133.385 ;
      VIA 55.72 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 126.375 56.51 126.705 ;
      VIA 55.72 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 126.355 56.49 126.725 ;
      VIA 55.72 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 119.715 56.51 120.045 ;
      VIA 55.72 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 119.695 56.49 120.065 ;
      VIA 55.72 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 113.055 56.51 113.385 ;
      VIA 55.72 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 113.035 56.49 113.405 ;
      VIA 55.72 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 106.395 56.51 106.725 ;
      VIA 55.72 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 106.375 56.49 106.745 ;
      VIA 55.72 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 99.735 56.51 100.065 ;
      VIA 55.72 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 99.715 56.49 100.085 ;
      VIA 55.72 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 93.075 56.51 93.405 ;
      VIA 55.72 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 93.055 56.49 93.425 ;
      VIA 55.72 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 86.415 56.51 86.745 ;
      VIA 55.72 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 86.395 56.49 86.765 ;
      VIA 55.72 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 79.755 56.51 80.085 ;
      VIA 55.72 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 79.735 56.49 80.105 ;
      VIA 55.72 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 73.095 56.51 73.425 ;
      VIA 55.72 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 73.075 56.49 73.445 ;
      VIA 55.72 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 66.435 56.51 66.765 ;
      VIA 55.72 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 66.415 56.49 66.785 ;
      VIA 55.72 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 59.775 56.51 60.105 ;
      VIA 55.72 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 59.755 56.49 60.125 ;
      VIA 55.72 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 53.115 56.51 53.445 ;
      VIA 55.72 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 53.095 56.49 53.465 ;
      VIA 55.72 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 46.455 56.51 46.785 ;
      VIA 55.72 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 46.435 56.49 46.805 ;
      VIA 55.72 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 39.795 56.51 40.125 ;
      VIA 55.72 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 39.775 56.49 40.145 ;
      VIA 55.72 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 33.135 56.51 33.465 ;
      VIA 55.72 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 33.115 56.49 33.485 ;
      VIA 55.72 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 26.475 56.51 26.805 ;
      VIA 55.72 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 26.455 56.49 26.825 ;
      VIA 55.72 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 19.815 56.51 20.145 ;
      VIA 55.72 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 19.795 56.49 20.165 ;
      VIA 55.72 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 13.155 56.51 13.485 ;
      VIA 55.72 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 13.135 56.49 13.505 ;
      VIA 55.72 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.93 6.495 56.51 6.825 ;
      VIA 55.72 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.95 6.475 56.49 6.845 ;
      VIA 55.72 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 55.72 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 779.055 29.37 779.385 ;
      VIA 28.58 779.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 779.035 29.35 779.405 ;
      VIA 28.58 779.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 779.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 772.395 29.37 772.725 ;
      VIA 28.58 772.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 772.375 29.35 772.745 ;
      VIA 28.58 772.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 772.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 765.735 29.37 766.065 ;
      VIA 28.58 765.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 765.715 29.35 766.085 ;
      VIA 28.58 765.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 765.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 759.075 29.37 759.405 ;
      VIA 28.58 759.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 759.055 29.35 759.425 ;
      VIA 28.58 759.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 759.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 752.415 29.37 752.745 ;
      VIA 28.58 752.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 752.395 29.35 752.765 ;
      VIA 28.58 752.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 752.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 745.755 29.37 746.085 ;
      VIA 28.58 745.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 745.735 29.35 746.105 ;
      VIA 28.58 745.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 745.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 739.095 29.37 739.425 ;
      VIA 28.58 739.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 739.075 29.35 739.445 ;
      VIA 28.58 739.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 739.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 732.435 29.37 732.765 ;
      VIA 28.58 732.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 732.415 29.35 732.785 ;
      VIA 28.58 732.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 732.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 725.775 29.37 726.105 ;
      VIA 28.58 725.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 725.755 29.35 726.125 ;
      VIA 28.58 725.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 725.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 719.115 29.37 719.445 ;
      VIA 28.58 719.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 719.095 29.35 719.465 ;
      VIA 28.58 719.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 719.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 712.455 29.37 712.785 ;
      VIA 28.58 712.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 712.435 29.35 712.805 ;
      VIA 28.58 712.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 712.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 705.795 29.37 706.125 ;
      VIA 28.58 705.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 705.775 29.35 706.145 ;
      VIA 28.58 705.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 705.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 699.135 29.37 699.465 ;
      VIA 28.58 699.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 699.115 29.35 699.485 ;
      VIA 28.58 699.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 699.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 692.475 29.37 692.805 ;
      VIA 28.58 692.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 692.455 29.35 692.825 ;
      VIA 28.58 692.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 692.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 685.815 29.37 686.145 ;
      VIA 28.58 685.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 685.795 29.35 686.165 ;
      VIA 28.58 685.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 685.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 679.155 29.37 679.485 ;
      VIA 28.58 679.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 679.135 29.35 679.505 ;
      VIA 28.58 679.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 679.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 672.495 29.37 672.825 ;
      VIA 28.58 672.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 672.475 29.35 672.845 ;
      VIA 28.58 672.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 672.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 665.835 29.37 666.165 ;
      VIA 28.58 666 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 665.815 29.35 666.185 ;
      VIA 28.58 666 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 666 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 659.175 29.37 659.505 ;
      VIA 28.58 659.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 659.155 29.35 659.525 ;
      VIA 28.58 659.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 659.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 652.515 29.37 652.845 ;
      VIA 28.58 652.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 652.495 29.35 652.865 ;
      VIA 28.58 652.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 652.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 645.855 29.37 646.185 ;
      VIA 28.58 646.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 645.835 29.35 646.205 ;
      VIA 28.58 646.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 646.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 639.195 29.37 639.525 ;
      VIA 28.58 639.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 639.175 29.35 639.545 ;
      VIA 28.58 639.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 639.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 632.535 29.37 632.865 ;
      VIA 28.58 632.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 632.515 29.35 632.885 ;
      VIA 28.58 632.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 632.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 625.875 29.37 626.205 ;
      VIA 28.58 626.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 625.855 29.35 626.225 ;
      VIA 28.58 626.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 626.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 619.215 29.37 619.545 ;
      VIA 28.58 619.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 619.195 29.35 619.565 ;
      VIA 28.58 619.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 619.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 612.555 29.37 612.885 ;
      VIA 28.58 612.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 612.535 29.35 612.905 ;
      VIA 28.58 612.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 612.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 605.895 29.37 606.225 ;
      VIA 28.58 606.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 605.875 29.35 606.245 ;
      VIA 28.58 606.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 606.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 599.235 29.37 599.565 ;
      VIA 28.58 599.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 599.215 29.35 599.585 ;
      VIA 28.58 599.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 599.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 592.575 29.37 592.905 ;
      VIA 28.58 592.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 592.555 29.35 592.925 ;
      VIA 28.58 592.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 592.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 585.915 29.37 586.245 ;
      VIA 28.58 586.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 585.895 29.35 586.265 ;
      VIA 28.58 586.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 586.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 579.255 29.37 579.585 ;
      VIA 28.58 579.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 579.235 29.35 579.605 ;
      VIA 28.58 579.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 579.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 572.595 29.37 572.925 ;
      VIA 28.58 572.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 572.575 29.35 572.945 ;
      VIA 28.58 572.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 572.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 565.935 29.37 566.265 ;
      VIA 28.58 566.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 565.915 29.35 566.285 ;
      VIA 28.58 566.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 566.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 559.275 29.37 559.605 ;
      VIA 28.58 559.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 559.255 29.35 559.625 ;
      VIA 28.58 559.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 559.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 552.615 29.37 552.945 ;
      VIA 28.58 552.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 552.595 29.35 552.965 ;
      VIA 28.58 552.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 552.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 545.955 29.37 546.285 ;
      VIA 28.58 546.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 545.935 29.35 546.305 ;
      VIA 28.58 546.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 546.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 539.295 29.37 539.625 ;
      VIA 28.58 539.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 539.275 29.35 539.645 ;
      VIA 28.58 539.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 539.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 532.635 29.37 532.965 ;
      VIA 28.58 532.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 532.615 29.35 532.985 ;
      VIA 28.58 532.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 532.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 525.975 29.37 526.305 ;
      VIA 28.58 526.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 525.955 29.35 526.325 ;
      VIA 28.58 526.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 526.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 519.315 29.37 519.645 ;
      VIA 28.58 519.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 519.295 29.35 519.665 ;
      VIA 28.58 519.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 519.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 512.655 29.37 512.985 ;
      VIA 28.58 512.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 512.635 29.35 513.005 ;
      VIA 28.58 512.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 512.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 505.995 29.37 506.325 ;
      VIA 28.58 506.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 505.975 29.35 506.345 ;
      VIA 28.58 506.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 506.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 499.335 29.37 499.665 ;
      VIA 28.58 499.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 499.315 29.35 499.685 ;
      VIA 28.58 499.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 499.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 492.675 29.37 493.005 ;
      VIA 28.58 492.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 492.655 29.35 493.025 ;
      VIA 28.58 492.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 492.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 486.015 29.37 486.345 ;
      VIA 28.58 486.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 485.995 29.35 486.365 ;
      VIA 28.58 486.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 486.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 479.355 29.37 479.685 ;
      VIA 28.58 479.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 479.335 29.35 479.705 ;
      VIA 28.58 479.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 479.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 472.695 29.37 473.025 ;
      VIA 28.58 472.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 472.675 29.35 473.045 ;
      VIA 28.58 472.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 472.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 466.035 29.37 466.365 ;
      VIA 28.58 466.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 466.015 29.35 466.385 ;
      VIA 28.58 466.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 466.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 459.375 29.37 459.705 ;
      VIA 28.58 459.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 459.355 29.35 459.725 ;
      VIA 28.58 459.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 459.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 452.715 29.37 453.045 ;
      VIA 28.58 452.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 452.695 29.35 453.065 ;
      VIA 28.58 452.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 452.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 446.055 29.37 446.385 ;
      VIA 28.58 446.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 446.035 29.35 446.405 ;
      VIA 28.58 446.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 446.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 439.395 29.37 439.725 ;
      VIA 28.58 439.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 439.375 29.35 439.745 ;
      VIA 28.58 439.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 439.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 432.735 29.37 433.065 ;
      VIA 28.58 432.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 432.715 29.35 433.085 ;
      VIA 28.58 432.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 432.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 426.075 29.37 426.405 ;
      VIA 28.58 426.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 426.055 29.35 426.425 ;
      VIA 28.58 426.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 426.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 419.415 29.37 419.745 ;
      VIA 28.58 419.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 419.395 29.35 419.765 ;
      VIA 28.58 419.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 419.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 412.755 29.37 413.085 ;
      VIA 28.58 412.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 412.735 29.35 413.105 ;
      VIA 28.58 412.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 412.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 406.095 29.37 406.425 ;
      VIA 28.58 406.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 406.075 29.35 406.445 ;
      VIA 28.58 406.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 406.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 399.435 29.37 399.765 ;
      VIA 28.58 399.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 399.415 29.35 399.785 ;
      VIA 28.58 399.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 399.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 392.775 29.37 393.105 ;
      VIA 28.58 392.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 392.755 29.35 393.125 ;
      VIA 28.58 392.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 392.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 386.115 29.37 386.445 ;
      VIA 28.58 386.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 386.095 29.35 386.465 ;
      VIA 28.58 386.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 386.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 379.455 29.37 379.785 ;
      VIA 28.58 379.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 379.435 29.35 379.805 ;
      VIA 28.58 379.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 379.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 372.795 29.37 373.125 ;
      VIA 28.58 372.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 372.775 29.35 373.145 ;
      VIA 28.58 372.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 372.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 366.135 29.37 366.465 ;
      VIA 28.58 366.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 366.115 29.35 366.485 ;
      VIA 28.58 366.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 366.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 359.475 29.37 359.805 ;
      VIA 28.58 359.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 359.455 29.35 359.825 ;
      VIA 28.58 359.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 359.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 352.815 29.37 353.145 ;
      VIA 28.58 352.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 352.795 29.35 353.165 ;
      VIA 28.58 352.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 352.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 346.155 29.37 346.485 ;
      VIA 28.58 346.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 346.135 29.35 346.505 ;
      VIA 28.58 346.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 346.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 339.495 29.37 339.825 ;
      VIA 28.58 339.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 339.475 29.35 339.845 ;
      VIA 28.58 339.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 339.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 332.835 29.37 333.165 ;
      VIA 28.58 333 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 332.815 29.35 333.185 ;
      VIA 28.58 333 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 333 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 326.175 29.37 326.505 ;
      VIA 28.58 326.34 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 326.155 29.35 326.525 ;
      VIA 28.58 326.34 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 326.34 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 319.515 29.37 319.845 ;
      VIA 28.58 319.68 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 319.495 29.35 319.865 ;
      VIA 28.58 319.68 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 319.68 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 312.855 29.37 313.185 ;
      VIA 28.58 313.02 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 312.835 29.35 313.205 ;
      VIA 28.58 313.02 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 313.02 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 306.195 29.37 306.525 ;
      VIA 28.58 306.36 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 306.175 29.35 306.545 ;
      VIA 28.58 306.36 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 306.36 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 299.535 29.37 299.865 ;
      VIA 28.58 299.7 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 299.515 29.35 299.885 ;
      VIA 28.58 299.7 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 299.7 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 292.875 29.37 293.205 ;
      VIA 28.58 293.04 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 292.855 29.35 293.225 ;
      VIA 28.58 293.04 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 293.04 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 286.215 29.37 286.545 ;
      VIA 28.58 286.38 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 286.195 29.35 286.565 ;
      VIA 28.58 286.38 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 286.38 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 279.555 29.37 279.885 ;
      VIA 28.58 279.72 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 279.535 29.35 279.905 ;
      VIA 28.58 279.72 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 279.72 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 272.895 29.37 273.225 ;
      VIA 28.58 273.06 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 272.875 29.35 273.245 ;
      VIA 28.58 273.06 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 273.06 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 266.235 29.37 266.565 ;
      VIA 28.58 266.4 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 266.215 29.35 266.585 ;
      VIA 28.58 266.4 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 266.4 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 259.575 29.37 259.905 ;
      VIA 28.58 259.74 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 259.555 29.35 259.925 ;
      VIA 28.58 259.74 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 259.74 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 252.915 29.37 253.245 ;
      VIA 28.58 253.08 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 252.895 29.35 253.265 ;
      VIA 28.58 253.08 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 253.08 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 246.255 29.37 246.585 ;
      VIA 28.58 246.42 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 246.235 29.35 246.605 ;
      VIA 28.58 246.42 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 246.42 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 239.595 29.37 239.925 ;
      VIA 28.58 239.76 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 239.575 29.35 239.945 ;
      VIA 28.58 239.76 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 239.76 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 232.935 29.37 233.265 ;
      VIA 28.58 233.1 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 232.915 29.35 233.285 ;
      VIA 28.58 233.1 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 233.1 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 226.275 29.37 226.605 ;
      VIA 28.58 226.44 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 226.255 29.35 226.625 ;
      VIA 28.58 226.44 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 226.44 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 219.615 29.37 219.945 ;
      VIA 28.58 219.78 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 219.595 29.35 219.965 ;
      VIA 28.58 219.78 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 219.78 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 212.955 29.37 213.285 ;
      VIA 28.58 213.12 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 212.935 29.35 213.305 ;
      VIA 28.58 213.12 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 213.12 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 206.295 29.37 206.625 ;
      VIA 28.58 206.46 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 206.275 29.35 206.645 ;
      VIA 28.58 206.46 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 206.46 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 199.635 29.37 199.965 ;
      VIA 28.58 199.8 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 199.615 29.35 199.985 ;
      VIA 28.58 199.8 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 199.8 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 192.975 29.37 193.305 ;
      VIA 28.58 193.14 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 192.955 29.35 193.325 ;
      VIA 28.58 193.14 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 193.14 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 186.315 29.37 186.645 ;
      VIA 28.58 186.48 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 186.295 29.35 186.665 ;
      VIA 28.58 186.48 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 186.48 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 179.655 29.37 179.985 ;
      VIA 28.58 179.82 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 179.635 29.35 180.005 ;
      VIA 28.58 179.82 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 179.82 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 172.995 29.37 173.325 ;
      VIA 28.58 173.16 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 172.975 29.35 173.345 ;
      VIA 28.58 173.16 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 173.16 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 166.335 29.37 166.665 ;
      VIA 28.58 166.5 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 166.315 29.35 166.685 ;
      VIA 28.58 166.5 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 166.5 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 159.675 29.37 160.005 ;
      VIA 28.58 159.84 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 159.655 29.35 160.025 ;
      VIA 28.58 159.84 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 159.84 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 153.015 29.37 153.345 ;
      VIA 28.58 153.18 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 152.995 29.35 153.365 ;
      VIA 28.58 153.18 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 153.18 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 146.355 29.37 146.685 ;
      VIA 28.58 146.52 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 146.335 29.35 146.705 ;
      VIA 28.58 146.52 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 146.52 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 139.695 29.37 140.025 ;
      VIA 28.58 139.86 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 139.675 29.35 140.045 ;
      VIA 28.58 139.86 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 139.86 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 133.035 29.37 133.365 ;
      VIA 28.58 133.2 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 133.015 29.35 133.385 ;
      VIA 28.58 133.2 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 133.2 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 126.375 29.37 126.705 ;
      VIA 28.58 126.54 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 126.355 29.35 126.725 ;
      VIA 28.58 126.54 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 126.54 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 119.715 29.37 120.045 ;
      VIA 28.58 119.88 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 119.695 29.35 120.065 ;
      VIA 28.58 119.88 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 119.88 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 113.055 29.37 113.385 ;
      VIA 28.58 113.22 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 113.035 29.35 113.405 ;
      VIA 28.58 113.22 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 113.22 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 106.395 29.37 106.725 ;
      VIA 28.58 106.56 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 106.375 29.35 106.745 ;
      VIA 28.58 106.56 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 106.56 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 99.735 29.37 100.065 ;
      VIA 28.58 99.9 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 99.715 29.35 100.085 ;
      VIA 28.58 99.9 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 99.9 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 93.075 29.37 93.405 ;
      VIA 28.58 93.24 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 93.055 29.35 93.425 ;
      VIA 28.58 93.24 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 93.24 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 86.415 29.37 86.745 ;
      VIA 28.58 86.58 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 86.395 29.35 86.765 ;
      VIA 28.58 86.58 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 86.58 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 79.755 29.37 80.085 ;
      VIA 28.58 79.92 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 79.735 29.35 80.105 ;
      VIA 28.58 79.92 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 79.92 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 73.095 29.37 73.425 ;
      VIA 28.58 73.26 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 73.075 29.35 73.445 ;
      VIA 28.58 73.26 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 73.26 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 66.435 29.37 66.765 ;
      VIA 28.58 66.6 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 66.415 29.35 66.785 ;
      VIA 28.58 66.6 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 66.6 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 59.775 29.37 60.105 ;
      VIA 28.58 59.94 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 59.755 29.35 60.125 ;
      VIA 28.58 59.94 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 59.94 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 53.115 29.37 53.445 ;
      VIA 28.58 53.28 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 53.095 29.35 53.465 ;
      VIA 28.58 53.28 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 53.28 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 46.455 29.37 46.785 ;
      VIA 28.58 46.62 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 46.435 29.35 46.805 ;
      VIA 28.58 46.62 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 46.62 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 39.795 29.37 40.125 ;
      VIA 28.58 39.96 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 39.775 29.35 40.145 ;
      VIA 28.58 39.96 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 39.96 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 33.135 29.37 33.465 ;
      VIA 28.58 33.3 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 33.115 29.35 33.485 ;
      VIA 28.58 33.3 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 33.3 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 26.475 29.37 26.805 ;
      VIA 28.58 26.64 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 26.455 29.35 26.825 ;
      VIA 28.58 26.64 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 26.64 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 19.815 29.37 20.145 ;
      VIA 28.58 19.98 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 19.795 29.35 20.165 ;
      VIA 28.58 19.98 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 19.98 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 13.155 29.37 13.485 ;
      VIA 28.58 13.32 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 13.135 29.35 13.505 ;
      VIA 28.58 13.32 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 13.32 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.79 6.495 29.37 6.825 ;
      VIA 28.58 6.66 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.81 6.475 29.35 6.845 ;
      VIA 28.58 6.66 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 28.58 6.66 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  14.21 777.73 260.07 779.33 ;
        RECT  14.21 750.53 260.07 752.13 ;
        RECT  14.21 723.33 260.07 724.93 ;
        RECT  14.21 696.13 260.07 697.73 ;
        RECT  14.21 668.93 260.07 670.53 ;
        RECT  14.21 641.73 260.07 643.33 ;
        RECT  14.21 614.53 260.07 616.13 ;
        RECT  14.21 587.33 260.07 588.93 ;
        RECT  14.21 560.13 260.07 561.73 ;
        RECT  14.21 532.93 260.07 534.53 ;
        RECT  14.21 505.73 260.07 507.33 ;
        RECT  14.21 478.53 260.07 480.13 ;
        RECT  14.21 451.33 260.07 452.93 ;
        RECT  14.21 424.13 260.07 425.73 ;
        RECT  14.21 396.93 260.07 398.53 ;
        RECT  14.21 369.73 260.07 371.33 ;
        RECT  14.21 342.53 260.07 344.13 ;
        RECT  14.21 315.33 260.07 316.93 ;
        RECT  14.21 288.13 260.07 289.73 ;
        RECT  14.21 260.93 260.07 262.53 ;
        RECT  14.21 233.73 260.07 235.33 ;
        RECT  14.21 206.53 260.07 208.13 ;
        RECT  14.21 179.33 260.07 180.93 ;
        RECT  14.21 152.13 260.07 153.73 ;
        RECT  14.21 124.93 260.07 126.53 ;
        RECT  14.21 97.73 260.07 99.33 ;
        RECT  14.21 70.53 260.07 72.13 ;
        RECT  14.21 43.33 260.07 44.93 ;
        RECT  14.21 16.13 260.07 17.73 ;
      LAYER met4 ;
        RECT  258.47 3.09 260.07 779.33 ;
        RECT  231.33 3.09 232.93 779.33 ;
        RECT  204.19 3.09 205.79 779.33 ;
        RECT  177.05 3.09 178.65 779.33 ;
        RECT  149.91 3.09 151.51 779.33 ;
        RECT  122.77 3.09 124.37 779.33 ;
        RECT  95.63 3.09 97.23 779.33 ;
        RECT  68.49 3.09 70.09 779.33 ;
        RECT  41.35 3.09 42.95 779.33 ;
        RECT  14.21 3.09 15.81 779.33 ;
      LAYER met1 ;
        RECT  1.44 775.65 260.64 776.13 ;
        RECT  1.44 768.99 260.64 769.47 ;
        RECT  1.44 762.33 260.64 762.81 ;
        RECT  1.44 755.67 260.64 756.15 ;
        RECT  1.44 749.01 260.64 749.49 ;
        RECT  1.44 742.35 260.64 742.83 ;
        RECT  1.44 735.69 260.64 736.17 ;
        RECT  1.44 729.03 260.64 729.51 ;
        RECT  1.44 722.37 260.64 722.85 ;
        RECT  1.44 715.71 260.64 716.19 ;
        RECT  1.44 709.05 260.64 709.53 ;
        RECT  1.44 702.39 260.64 702.87 ;
        RECT  1.44 695.73 260.64 696.21 ;
        RECT  1.44 689.07 260.64 689.55 ;
        RECT  1.44 682.41 260.64 682.89 ;
        RECT  1.44 675.75 260.64 676.23 ;
        RECT  1.44 669.09 260.64 669.57 ;
        RECT  1.44 662.43 260.64 662.91 ;
        RECT  1.44 655.77 260.64 656.25 ;
        RECT  1.44 649.11 260.64 649.59 ;
        RECT  1.44 642.45 260.64 642.93 ;
        RECT  1.44 635.79 260.64 636.27 ;
        RECT  1.44 629.13 260.64 629.61 ;
        RECT  1.44 622.47 260.64 622.95 ;
        RECT  1.44 615.81 260.64 616.29 ;
        RECT  1.44 609.15 260.64 609.63 ;
        RECT  1.44 602.49 260.64 602.97 ;
        RECT  1.44 595.83 260.64 596.31 ;
        RECT  1.44 589.17 260.64 589.65 ;
        RECT  1.44 582.51 260.64 582.99 ;
        RECT  1.44 575.85 260.64 576.33 ;
        RECT  1.44 569.19 260.64 569.67 ;
        RECT  1.44 562.53 260.64 563.01 ;
        RECT  1.44 555.87 260.64 556.35 ;
        RECT  1.44 549.21 260.64 549.69 ;
        RECT  1.44 542.55 260.64 543.03 ;
        RECT  1.44 535.89 260.64 536.37 ;
        RECT  1.44 529.23 260.64 529.71 ;
        RECT  1.44 522.57 260.64 523.05 ;
        RECT  1.44 515.91 260.64 516.39 ;
        RECT  1.44 509.25 260.64 509.73 ;
        RECT  1.44 502.59 260.64 503.07 ;
        RECT  1.44 495.93 260.64 496.41 ;
        RECT  1.44 489.27 260.64 489.75 ;
        RECT  1.44 482.61 260.64 483.09 ;
        RECT  1.44 475.95 260.64 476.43 ;
        RECT  1.44 469.29 260.64 469.77 ;
        RECT  1.44 462.63 260.64 463.11 ;
        RECT  1.44 455.97 260.64 456.45 ;
        RECT  1.44 449.31 260.64 449.79 ;
        RECT  1.44 442.65 260.64 443.13 ;
        RECT  1.44 435.99 260.64 436.47 ;
        RECT  1.44 429.33 260.64 429.81 ;
        RECT  1.44 422.67 260.64 423.15 ;
        RECT  1.44 416.01 260.64 416.49 ;
        RECT  1.44 409.35 260.64 409.83 ;
        RECT  1.44 402.69 260.64 403.17 ;
        RECT  1.44 396.03 260.64 396.51 ;
        RECT  1.44 389.37 260.64 389.85 ;
        RECT  1.44 382.71 260.64 383.19 ;
        RECT  1.44 376.05 260.64 376.53 ;
        RECT  1.44 369.39 260.64 369.87 ;
        RECT  1.44 362.73 260.64 363.21 ;
        RECT  1.44 356.07 260.64 356.55 ;
        RECT  1.44 349.41 260.64 349.89 ;
        RECT  1.44 342.75 260.64 343.23 ;
        RECT  1.44 336.09 260.64 336.57 ;
        RECT  1.44 329.43 260.64 329.91 ;
        RECT  1.44 322.77 260.64 323.25 ;
        RECT  1.44 316.11 260.64 316.59 ;
        RECT  1.44 309.45 260.64 309.93 ;
        RECT  1.44 302.79 260.64 303.27 ;
        RECT  1.44 296.13 260.64 296.61 ;
        RECT  1.44 289.47 260.64 289.95 ;
        RECT  1.44 282.81 260.64 283.29 ;
        RECT  1.44 276.15 260.64 276.63 ;
        RECT  1.44 269.49 260.64 269.97 ;
        RECT  1.44 262.83 260.64 263.31 ;
        RECT  1.44 256.17 260.64 256.65 ;
        RECT  1.44 249.51 260.64 249.99 ;
        RECT  1.44 242.85 260.64 243.33 ;
        RECT  1.44 236.19 260.64 236.67 ;
        RECT  1.44 229.53 260.64 230.01 ;
        RECT  1.44 222.87 260.64 223.35 ;
        RECT  1.44 216.21 260.64 216.69 ;
        RECT  1.44 209.55 260.64 210.03 ;
        RECT  1.44 202.89 260.64 203.37 ;
        RECT  1.44 196.23 260.64 196.71 ;
        RECT  1.44 189.57 260.64 190.05 ;
        RECT  1.44 182.91 260.64 183.39 ;
        RECT  1.44 176.25 260.64 176.73 ;
        RECT  1.44 169.59 260.64 170.07 ;
        RECT  1.44 162.93 260.64 163.41 ;
        RECT  1.44 156.27 260.64 156.75 ;
        RECT  1.44 149.61 260.64 150.09 ;
        RECT  1.44 142.95 260.64 143.43 ;
        RECT  1.44 136.29 260.64 136.77 ;
        RECT  1.44 129.63 260.64 130.11 ;
        RECT  1.44 122.97 260.64 123.45 ;
        RECT  1.44 116.31 260.64 116.79 ;
        RECT  1.44 109.65 260.64 110.13 ;
        RECT  1.44 102.99 260.64 103.47 ;
        RECT  1.44 96.33 260.64 96.81 ;
        RECT  1.44 89.67 260.64 90.15 ;
        RECT  1.44 83.01 260.64 83.49 ;
        RECT  1.44 76.35 260.64 76.83 ;
        RECT  1.44 69.69 260.64 70.17 ;
        RECT  1.44 63.03 260.64 63.51 ;
        RECT  1.44 56.37 260.64 56.85 ;
        RECT  1.44 49.71 260.64 50.19 ;
        RECT  1.44 43.05 260.64 43.53 ;
        RECT  1.44 36.39 260.64 36.87 ;
        RECT  1.44 29.73 260.64 30.21 ;
        RECT  1.44 23.07 260.64 23.55 ;
        RECT  1.44 16.41 260.64 16.89 ;
        RECT  1.44 9.75 260.64 10.23 ;
        RECT  1.44 3.09 260.64 3.57 ;
      VIA 259.27 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 259.27 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 232.13 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 204.99 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 177.85 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.71 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.57 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.43 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.29 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.15 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 778.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 751.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 724.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 696.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 669.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 642.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 615.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 588.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 560.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 533.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 506.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 479.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 452.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 424.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 397.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 370.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 343.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 316.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 288.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 261.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 234.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 207.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 180.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 152.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 125.73 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 98.53 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 71.33 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 44.13 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 15.01 16.93 ibex_ex_block_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  258.48 775.725 260.06 776.055 ;
      VIA 259.27 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 775.705 260.04 776.075 ;
      VIA 259.27 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 769.065 260.06 769.395 ;
      VIA 259.27 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 769.045 260.04 769.415 ;
      VIA 259.27 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 762.405 260.06 762.735 ;
      VIA 259.27 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 762.385 260.04 762.755 ;
      VIA 259.27 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 755.745 260.06 756.075 ;
      VIA 259.27 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 755.725 260.04 756.095 ;
      VIA 259.27 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 749.085 260.06 749.415 ;
      VIA 259.27 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 749.065 260.04 749.435 ;
      VIA 259.27 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 742.425 260.06 742.755 ;
      VIA 259.27 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 742.405 260.04 742.775 ;
      VIA 259.27 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 735.765 260.06 736.095 ;
      VIA 259.27 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 735.745 260.04 736.115 ;
      VIA 259.27 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 729.105 260.06 729.435 ;
      VIA 259.27 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 729.085 260.04 729.455 ;
      VIA 259.27 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 722.445 260.06 722.775 ;
      VIA 259.27 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 722.425 260.04 722.795 ;
      VIA 259.27 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 715.785 260.06 716.115 ;
      VIA 259.27 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 715.765 260.04 716.135 ;
      VIA 259.27 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 709.125 260.06 709.455 ;
      VIA 259.27 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 709.105 260.04 709.475 ;
      VIA 259.27 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 702.465 260.06 702.795 ;
      VIA 259.27 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 702.445 260.04 702.815 ;
      VIA 259.27 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 695.805 260.06 696.135 ;
      VIA 259.27 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 695.785 260.04 696.155 ;
      VIA 259.27 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 689.145 260.06 689.475 ;
      VIA 259.27 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 689.125 260.04 689.495 ;
      VIA 259.27 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 682.485 260.06 682.815 ;
      VIA 259.27 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 682.465 260.04 682.835 ;
      VIA 259.27 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 675.825 260.06 676.155 ;
      VIA 259.27 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 675.805 260.04 676.175 ;
      VIA 259.27 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 669.165 260.06 669.495 ;
      VIA 259.27 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 669.145 260.04 669.515 ;
      VIA 259.27 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 662.505 260.06 662.835 ;
      VIA 259.27 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 662.485 260.04 662.855 ;
      VIA 259.27 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 655.845 260.06 656.175 ;
      VIA 259.27 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 655.825 260.04 656.195 ;
      VIA 259.27 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 649.185 260.06 649.515 ;
      VIA 259.27 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 649.165 260.04 649.535 ;
      VIA 259.27 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 642.525 260.06 642.855 ;
      VIA 259.27 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 642.505 260.04 642.875 ;
      VIA 259.27 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 635.865 260.06 636.195 ;
      VIA 259.27 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 635.845 260.04 636.215 ;
      VIA 259.27 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 629.205 260.06 629.535 ;
      VIA 259.27 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 629.185 260.04 629.555 ;
      VIA 259.27 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 622.545 260.06 622.875 ;
      VIA 259.27 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 622.525 260.04 622.895 ;
      VIA 259.27 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 615.885 260.06 616.215 ;
      VIA 259.27 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 615.865 260.04 616.235 ;
      VIA 259.27 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 609.225 260.06 609.555 ;
      VIA 259.27 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 609.205 260.04 609.575 ;
      VIA 259.27 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 602.565 260.06 602.895 ;
      VIA 259.27 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 602.545 260.04 602.915 ;
      VIA 259.27 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 595.905 260.06 596.235 ;
      VIA 259.27 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 595.885 260.04 596.255 ;
      VIA 259.27 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 589.245 260.06 589.575 ;
      VIA 259.27 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 589.225 260.04 589.595 ;
      VIA 259.27 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 582.585 260.06 582.915 ;
      VIA 259.27 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 582.565 260.04 582.935 ;
      VIA 259.27 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 575.925 260.06 576.255 ;
      VIA 259.27 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 575.905 260.04 576.275 ;
      VIA 259.27 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 569.265 260.06 569.595 ;
      VIA 259.27 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 569.245 260.04 569.615 ;
      VIA 259.27 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 562.605 260.06 562.935 ;
      VIA 259.27 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 562.585 260.04 562.955 ;
      VIA 259.27 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 555.945 260.06 556.275 ;
      VIA 259.27 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 555.925 260.04 556.295 ;
      VIA 259.27 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 549.285 260.06 549.615 ;
      VIA 259.27 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 549.265 260.04 549.635 ;
      VIA 259.27 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 542.625 260.06 542.955 ;
      VIA 259.27 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 542.605 260.04 542.975 ;
      VIA 259.27 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 535.965 260.06 536.295 ;
      VIA 259.27 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 535.945 260.04 536.315 ;
      VIA 259.27 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 529.305 260.06 529.635 ;
      VIA 259.27 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 529.285 260.04 529.655 ;
      VIA 259.27 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 522.645 260.06 522.975 ;
      VIA 259.27 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 522.625 260.04 522.995 ;
      VIA 259.27 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 515.985 260.06 516.315 ;
      VIA 259.27 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 515.965 260.04 516.335 ;
      VIA 259.27 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 509.325 260.06 509.655 ;
      VIA 259.27 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 509.305 260.04 509.675 ;
      VIA 259.27 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 502.665 260.06 502.995 ;
      VIA 259.27 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 502.645 260.04 503.015 ;
      VIA 259.27 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 496.005 260.06 496.335 ;
      VIA 259.27 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 495.985 260.04 496.355 ;
      VIA 259.27 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 489.345 260.06 489.675 ;
      VIA 259.27 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 489.325 260.04 489.695 ;
      VIA 259.27 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 482.685 260.06 483.015 ;
      VIA 259.27 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 482.665 260.04 483.035 ;
      VIA 259.27 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 476.025 260.06 476.355 ;
      VIA 259.27 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 476.005 260.04 476.375 ;
      VIA 259.27 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 469.365 260.06 469.695 ;
      VIA 259.27 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 469.345 260.04 469.715 ;
      VIA 259.27 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 462.705 260.06 463.035 ;
      VIA 259.27 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 462.685 260.04 463.055 ;
      VIA 259.27 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 456.045 260.06 456.375 ;
      VIA 259.27 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 456.025 260.04 456.395 ;
      VIA 259.27 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 449.385 260.06 449.715 ;
      VIA 259.27 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 449.365 260.04 449.735 ;
      VIA 259.27 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 442.725 260.06 443.055 ;
      VIA 259.27 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 442.705 260.04 443.075 ;
      VIA 259.27 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 436.065 260.06 436.395 ;
      VIA 259.27 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 436.045 260.04 436.415 ;
      VIA 259.27 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 429.405 260.06 429.735 ;
      VIA 259.27 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 429.385 260.04 429.755 ;
      VIA 259.27 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 422.745 260.06 423.075 ;
      VIA 259.27 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 422.725 260.04 423.095 ;
      VIA 259.27 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 416.085 260.06 416.415 ;
      VIA 259.27 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 416.065 260.04 416.435 ;
      VIA 259.27 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 409.425 260.06 409.755 ;
      VIA 259.27 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 409.405 260.04 409.775 ;
      VIA 259.27 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 402.765 260.06 403.095 ;
      VIA 259.27 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 402.745 260.04 403.115 ;
      VIA 259.27 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 396.105 260.06 396.435 ;
      VIA 259.27 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 396.085 260.04 396.455 ;
      VIA 259.27 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 389.445 260.06 389.775 ;
      VIA 259.27 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 389.425 260.04 389.795 ;
      VIA 259.27 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 382.785 260.06 383.115 ;
      VIA 259.27 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 382.765 260.04 383.135 ;
      VIA 259.27 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 376.125 260.06 376.455 ;
      VIA 259.27 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 376.105 260.04 376.475 ;
      VIA 259.27 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 369.465 260.06 369.795 ;
      VIA 259.27 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 369.445 260.04 369.815 ;
      VIA 259.27 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 362.805 260.06 363.135 ;
      VIA 259.27 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 362.785 260.04 363.155 ;
      VIA 259.27 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 356.145 260.06 356.475 ;
      VIA 259.27 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 356.125 260.04 356.495 ;
      VIA 259.27 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 349.485 260.06 349.815 ;
      VIA 259.27 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 349.465 260.04 349.835 ;
      VIA 259.27 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 342.825 260.06 343.155 ;
      VIA 259.27 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 342.805 260.04 343.175 ;
      VIA 259.27 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 336.165 260.06 336.495 ;
      VIA 259.27 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 336.145 260.04 336.515 ;
      VIA 259.27 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 329.505 260.06 329.835 ;
      VIA 259.27 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 329.485 260.04 329.855 ;
      VIA 259.27 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 322.845 260.06 323.175 ;
      VIA 259.27 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 322.825 260.04 323.195 ;
      VIA 259.27 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 316.185 260.06 316.515 ;
      VIA 259.27 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 316.165 260.04 316.535 ;
      VIA 259.27 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 309.525 260.06 309.855 ;
      VIA 259.27 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 309.505 260.04 309.875 ;
      VIA 259.27 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 302.865 260.06 303.195 ;
      VIA 259.27 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 302.845 260.04 303.215 ;
      VIA 259.27 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 296.205 260.06 296.535 ;
      VIA 259.27 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 296.185 260.04 296.555 ;
      VIA 259.27 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 289.545 260.06 289.875 ;
      VIA 259.27 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 289.525 260.04 289.895 ;
      VIA 259.27 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 282.885 260.06 283.215 ;
      VIA 259.27 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 282.865 260.04 283.235 ;
      VIA 259.27 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 276.225 260.06 276.555 ;
      VIA 259.27 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 276.205 260.04 276.575 ;
      VIA 259.27 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 269.565 260.06 269.895 ;
      VIA 259.27 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 269.545 260.04 269.915 ;
      VIA 259.27 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 262.905 260.06 263.235 ;
      VIA 259.27 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 262.885 260.04 263.255 ;
      VIA 259.27 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 256.245 260.06 256.575 ;
      VIA 259.27 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 256.225 260.04 256.595 ;
      VIA 259.27 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 249.585 260.06 249.915 ;
      VIA 259.27 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 249.565 260.04 249.935 ;
      VIA 259.27 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 242.925 260.06 243.255 ;
      VIA 259.27 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 242.905 260.04 243.275 ;
      VIA 259.27 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 236.265 260.06 236.595 ;
      VIA 259.27 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 236.245 260.04 236.615 ;
      VIA 259.27 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 229.605 260.06 229.935 ;
      VIA 259.27 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 229.585 260.04 229.955 ;
      VIA 259.27 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 222.945 260.06 223.275 ;
      VIA 259.27 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 222.925 260.04 223.295 ;
      VIA 259.27 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 216.285 260.06 216.615 ;
      VIA 259.27 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 216.265 260.04 216.635 ;
      VIA 259.27 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 209.625 260.06 209.955 ;
      VIA 259.27 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 209.605 260.04 209.975 ;
      VIA 259.27 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 202.965 260.06 203.295 ;
      VIA 259.27 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 202.945 260.04 203.315 ;
      VIA 259.27 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 196.305 260.06 196.635 ;
      VIA 259.27 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 196.285 260.04 196.655 ;
      VIA 259.27 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 189.645 260.06 189.975 ;
      VIA 259.27 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 189.625 260.04 189.995 ;
      VIA 259.27 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 182.985 260.06 183.315 ;
      VIA 259.27 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 182.965 260.04 183.335 ;
      VIA 259.27 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 176.325 260.06 176.655 ;
      VIA 259.27 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 176.305 260.04 176.675 ;
      VIA 259.27 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 169.665 260.06 169.995 ;
      VIA 259.27 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 169.645 260.04 170.015 ;
      VIA 259.27 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 163.005 260.06 163.335 ;
      VIA 259.27 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 162.985 260.04 163.355 ;
      VIA 259.27 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 156.345 260.06 156.675 ;
      VIA 259.27 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 156.325 260.04 156.695 ;
      VIA 259.27 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 149.685 260.06 150.015 ;
      VIA 259.27 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 149.665 260.04 150.035 ;
      VIA 259.27 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 143.025 260.06 143.355 ;
      VIA 259.27 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 143.005 260.04 143.375 ;
      VIA 259.27 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 136.365 260.06 136.695 ;
      VIA 259.27 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 136.345 260.04 136.715 ;
      VIA 259.27 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 129.705 260.06 130.035 ;
      VIA 259.27 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 129.685 260.04 130.055 ;
      VIA 259.27 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 123.045 260.06 123.375 ;
      VIA 259.27 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 123.025 260.04 123.395 ;
      VIA 259.27 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 116.385 260.06 116.715 ;
      VIA 259.27 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 116.365 260.04 116.735 ;
      VIA 259.27 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 109.725 260.06 110.055 ;
      VIA 259.27 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 109.705 260.04 110.075 ;
      VIA 259.27 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 103.065 260.06 103.395 ;
      VIA 259.27 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 103.045 260.04 103.415 ;
      VIA 259.27 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 96.405 260.06 96.735 ;
      VIA 259.27 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 96.385 260.04 96.755 ;
      VIA 259.27 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 89.745 260.06 90.075 ;
      VIA 259.27 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 89.725 260.04 90.095 ;
      VIA 259.27 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 83.085 260.06 83.415 ;
      VIA 259.27 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 83.065 260.04 83.435 ;
      VIA 259.27 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 76.425 260.06 76.755 ;
      VIA 259.27 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 76.405 260.04 76.775 ;
      VIA 259.27 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 69.765 260.06 70.095 ;
      VIA 259.27 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 69.745 260.04 70.115 ;
      VIA 259.27 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 63.105 260.06 63.435 ;
      VIA 259.27 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 63.085 260.04 63.455 ;
      VIA 259.27 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 56.445 260.06 56.775 ;
      VIA 259.27 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 56.425 260.04 56.795 ;
      VIA 259.27 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 49.785 260.06 50.115 ;
      VIA 259.27 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 49.765 260.04 50.135 ;
      VIA 259.27 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 43.125 260.06 43.455 ;
      VIA 259.27 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 43.105 260.04 43.475 ;
      VIA 259.27 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 36.465 260.06 36.795 ;
      VIA 259.27 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 36.445 260.04 36.815 ;
      VIA 259.27 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 29.805 260.06 30.135 ;
      VIA 259.27 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 29.785 260.04 30.155 ;
      VIA 259.27 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 23.145 260.06 23.475 ;
      VIA 259.27 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 23.125 260.04 23.495 ;
      VIA 259.27 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 16.485 260.06 16.815 ;
      VIA 259.27 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 16.465 260.04 16.835 ;
      VIA 259.27 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 9.825 260.06 10.155 ;
      VIA 259.27 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 9.805 260.04 10.175 ;
      VIA 259.27 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  258.48 3.165 260.06 3.495 ;
      VIA 259.27 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  258.5 3.145 260.04 3.515 ;
      VIA 259.27 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 259.27 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 775.725 232.92 776.055 ;
      VIA 232.13 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 775.705 232.9 776.075 ;
      VIA 232.13 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 769.065 232.92 769.395 ;
      VIA 232.13 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 769.045 232.9 769.415 ;
      VIA 232.13 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 762.405 232.92 762.735 ;
      VIA 232.13 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 762.385 232.9 762.755 ;
      VIA 232.13 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 755.745 232.92 756.075 ;
      VIA 232.13 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 755.725 232.9 756.095 ;
      VIA 232.13 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 749.085 232.92 749.415 ;
      VIA 232.13 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 749.065 232.9 749.435 ;
      VIA 232.13 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 742.425 232.92 742.755 ;
      VIA 232.13 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 742.405 232.9 742.775 ;
      VIA 232.13 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 735.765 232.92 736.095 ;
      VIA 232.13 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 735.745 232.9 736.115 ;
      VIA 232.13 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 729.105 232.92 729.435 ;
      VIA 232.13 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 729.085 232.9 729.455 ;
      VIA 232.13 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 722.445 232.92 722.775 ;
      VIA 232.13 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 722.425 232.9 722.795 ;
      VIA 232.13 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 715.785 232.92 716.115 ;
      VIA 232.13 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 715.765 232.9 716.135 ;
      VIA 232.13 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 709.125 232.92 709.455 ;
      VIA 232.13 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 709.105 232.9 709.475 ;
      VIA 232.13 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 702.465 232.92 702.795 ;
      VIA 232.13 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 702.445 232.9 702.815 ;
      VIA 232.13 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 695.805 232.92 696.135 ;
      VIA 232.13 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 695.785 232.9 696.155 ;
      VIA 232.13 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 689.145 232.92 689.475 ;
      VIA 232.13 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 689.125 232.9 689.495 ;
      VIA 232.13 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 682.485 232.92 682.815 ;
      VIA 232.13 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 682.465 232.9 682.835 ;
      VIA 232.13 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 675.825 232.92 676.155 ;
      VIA 232.13 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 675.805 232.9 676.175 ;
      VIA 232.13 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 669.165 232.92 669.495 ;
      VIA 232.13 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 669.145 232.9 669.515 ;
      VIA 232.13 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 662.505 232.92 662.835 ;
      VIA 232.13 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 662.485 232.9 662.855 ;
      VIA 232.13 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 655.845 232.92 656.175 ;
      VIA 232.13 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 655.825 232.9 656.195 ;
      VIA 232.13 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 649.185 232.92 649.515 ;
      VIA 232.13 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 649.165 232.9 649.535 ;
      VIA 232.13 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 642.525 232.92 642.855 ;
      VIA 232.13 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 642.505 232.9 642.875 ;
      VIA 232.13 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 635.865 232.92 636.195 ;
      VIA 232.13 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 635.845 232.9 636.215 ;
      VIA 232.13 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 629.205 232.92 629.535 ;
      VIA 232.13 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 629.185 232.9 629.555 ;
      VIA 232.13 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 622.545 232.92 622.875 ;
      VIA 232.13 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 622.525 232.9 622.895 ;
      VIA 232.13 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 615.885 232.92 616.215 ;
      VIA 232.13 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 615.865 232.9 616.235 ;
      VIA 232.13 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 609.225 232.92 609.555 ;
      VIA 232.13 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 609.205 232.9 609.575 ;
      VIA 232.13 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 602.565 232.92 602.895 ;
      VIA 232.13 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 602.545 232.9 602.915 ;
      VIA 232.13 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 595.905 232.92 596.235 ;
      VIA 232.13 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 595.885 232.9 596.255 ;
      VIA 232.13 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 589.245 232.92 589.575 ;
      VIA 232.13 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 589.225 232.9 589.595 ;
      VIA 232.13 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 582.585 232.92 582.915 ;
      VIA 232.13 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 582.565 232.9 582.935 ;
      VIA 232.13 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 575.925 232.92 576.255 ;
      VIA 232.13 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 575.905 232.9 576.275 ;
      VIA 232.13 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 569.265 232.92 569.595 ;
      VIA 232.13 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 569.245 232.9 569.615 ;
      VIA 232.13 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 562.605 232.92 562.935 ;
      VIA 232.13 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 562.585 232.9 562.955 ;
      VIA 232.13 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 555.945 232.92 556.275 ;
      VIA 232.13 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 555.925 232.9 556.295 ;
      VIA 232.13 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 549.285 232.92 549.615 ;
      VIA 232.13 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 549.265 232.9 549.635 ;
      VIA 232.13 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 542.625 232.92 542.955 ;
      VIA 232.13 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 542.605 232.9 542.975 ;
      VIA 232.13 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 535.965 232.92 536.295 ;
      VIA 232.13 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 535.945 232.9 536.315 ;
      VIA 232.13 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 529.305 232.92 529.635 ;
      VIA 232.13 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 529.285 232.9 529.655 ;
      VIA 232.13 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 522.645 232.92 522.975 ;
      VIA 232.13 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 522.625 232.9 522.995 ;
      VIA 232.13 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 515.985 232.92 516.315 ;
      VIA 232.13 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 515.965 232.9 516.335 ;
      VIA 232.13 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 509.325 232.92 509.655 ;
      VIA 232.13 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 509.305 232.9 509.675 ;
      VIA 232.13 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 502.665 232.92 502.995 ;
      VIA 232.13 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 502.645 232.9 503.015 ;
      VIA 232.13 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 496.005 232.92 496.335 ;
      VIA 232.13 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 495.985 232.9 496.355 ;
      VIA 232.13 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 489.345 232.92 489.675 ;
      VIA 232.13 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 489.325 232.9 489.695 ;
      VIA 232.13 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 482.685 232.92 483.015 ;
      VIA 232.13 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 482.665 232.9 483.035 ;
      VIA 232.13 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 476.025 232.92 476.355 ;
      VIA 232.13 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 476.005 232.9 476.375 ;
      VIA 232.13 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 469.365 232.92 469.695 ;
      VIA 232.13 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 469.345 232.9 469.715 ;
      VIA 232.13 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 462.705 232.92 463.035 ;
      VIA 232.13 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 462.685 232.9 463.055 ;
      VIA 232.13 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 456.045 232.92 456.375 ;
      VIA 232.13 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 456.025 232.9 456.395 ;
      VIA 232.13 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 449.385 232.92 449.715 ;
      VIA 232.13 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 449.365 232.9 449.735 ;
      VIA 232.13 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 442.725 232.92 443.055 ;
      VIA 232.13 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 442.705 232.9 443.075 ;
      VIA 232.13 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 436.065 232.92 436.395 ;
      VIA 232.13 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 436.045 232.9 436.415 ;
      VIA 232.13 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 429.405 232.92 429.735 ;
      VIA 232.13 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 429.385 232.9 429.755 ;
      VIA 232.13 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 422.745 232.92 423.075 ;
      VIA 232.13 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 422.725 232.9 423.095 ;
      VIA 232.13 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 416.085 232.92 416.415 ;
      VIA 232.13 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 416.065 232.9 416.435 ;
      VIA 232.13 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 409.425 232.92 409.755 ;
      VIA 232.13 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 409.405 232.9 409.775 ;
      VIA 232.13 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 402.765 232.92 403.095 ;
      VIA 232.13 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 402.745 232.9 403.115 ;
      VIA 232.13 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 396.105 232.92 396.435 ;
      VIA 232.13 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 396.085 232.9 396.455 ;
      VIA 232.13 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 389.445 232.92 389.775 ;
      VIA 232.13 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 389.425 232.9 389.795 ;
      VIA 232.13 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 382.785 232.92 383.115 ;
      VIA 232.13 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 382.765 232.9 383.135 ;
      VIA 232.13 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 376.125 232.92 376.455 ;
      VIA 232.13 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 376.105 232.9 376.475 ;
      VIA 232.13 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 369.465 232.92 369.795 ;
      VIA 232.13 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 369.445 232.9 369.815 ;
      VIA 232.13 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 362.805 232.92 363.135 ;
      VIA 232.13 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 362.785 232.9 363.155 ;
      VIA 232.13 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 356.145 232.92 356.475 ;
      VIA 232.13 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 356.125 232.9 356.495 ;
      VIA 232.13 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 349.485 232.92 349.815 ;
      VIA 232.13 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 349.465 232.9 349.835 ;
      VIA 232.13 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 342.825 232.92 343.155 ;
      VIA 232.13 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 342.805 232.9 343.175 ;
      VIA 232.13 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 336.165 232.92 336.495 ;
      VIA 232.13 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 336.145 232.9 336.515 ;
      VIA 232.13 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 329.505 232.92 329.835 ;
      VIA 232.13 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 329.485 232.9 329.855 ;
      VIA 232.13 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 322.845 232.92 323.175 ;
      VIA 232.13 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 322.825 232.9 323.195 ;
      VIA 232.13 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 316.185 232.92 316.515 ;
      VIA 232.13 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 316.165 232.9 316.535 ;
      VIA 232.13 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 309.525 232.92 309.855 ;
      VIA 232.13 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 309.505 232.9 309.875 ;
      VIA 232.13 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 302.865 232.92 303.195 ;
      VIA 232.13 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 302.845 232.9 303.215 ;
      VIA 232.13 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 296.205 232.92 296.535 ;
      VIA 232.13 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 296.185 232.9 296.555 ;
      VIA 232.13 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 289.545 232.92 289.875 ;
      VIA 232.13 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 289.525 232.9 289.895 ;
      VIA 232.13 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 282.885 232.92 283.215 ;
      VIA 232.13 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 282.865 232.9 283.235 ;
      VIA 232.13 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 276.225 232.92 276.555 ;
      VIA 232.13 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 276.205 232.9 276.575 ;
      VIA 232.13 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 269.565 232.92 269.895 ;
      VIA 232.13 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 269.545 232.9 269.915 ;
      VIA 232.13 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 262.905 232.92 263.235 ;
      VIA 232.13 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 262.885 232.9 263.255 ;
      VIA 232.13 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 256.245 232.92 256.575 ;
      VIA 232.13 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 256.225 232.9 256.595 ;
      VIA 232.13 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 249.585 232.92 249.915 ;
      VIA 232.13 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 249.565 232.9 249.935 ;
      VIA 232.13 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 242.925 232.92 243.255 ;
      VIA 232.13 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 242.905 232.9 243.275 ;
      VIA 232.13 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 236.265 232.92 236.595 ;
      VIA 232.13 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 236.245 232.9 236.615 ;
      VIA 232.13 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 229.605 232.92 229.935 ;
      VIA 232.13 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 229.585 232.9 229.955 ;
      VIA 232.13 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 222.945 232.92 223.275 ;
      VIA 232.13 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 222.925 232.9 223.295 ;
      VIA 232.13 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 216.285 232.92 216.615 ;
      VIA 232.13 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 216.265 232.9 216.635 ;
      VIA 232.13 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 209.625 232.92 209.955 ;
      VIA 232.13 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 209.605 232.9 209.975 ;
      VIA 232.13 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 202.965 232.92 203.295 ;
      VIA 232.13 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 202.945 232.9 203.315 ;
      VIA 232.13 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 196.305 232.92 196.635 ;
      VIA 232.13 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 196.285 232.9 196.655 ;
      VIA 232.13 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 189.645 232.92 189.975 ;
      VIA 232.13 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 189.625 232.9 189.995 ;
      VIA 232.13 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 182.985 232.92 183.315 ;
      VIA 232.13 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 182.965 232.9 183.335 ;
      VIA 232.13 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 176.325 232.92 176.655 ;
      VIA 232.13 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 176.305 232.9 176.675 ;
      VIA 232.13 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 169.665 232.92 169.995 ;
      VIA 232.13 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 169.645 232.9 170.015 ;
      VIA 232.13 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 163.005 232.92 163.335 ;
      VIA 232.13 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 162.985 232.9 163.355 ;
      VIA 232.13 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 156.345 232.92 156.675 ;
      VIA 232.13 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 156.325 232.9 156.695 ;
      VIA 232.13 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 149.685 232.92 150.015 ;
      VIA 232.13 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 149.665 232.9 150.035 ;
      VIA 232.13 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 143.025 232.92 143.355 ;
      VIA 232.13 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 143.005 232.9 143.375 ;
      VIA 232.13 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 136.365 232.92 136.695 ;
      VIA 232.13 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 136.345 232.9 136.715 ;
      VIA 232.13 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 129.705 232.92 130.035 ;
      VIA 232.13 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 129.685 232.9 130.055 ;
      VIA 232.13 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 123.045 232.92 123.375 ;
      VIA 232.13 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 123.025 232.9 123.395 ;
      VIA 232.13 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 116.385 232.92 116.715 ;
      VIA 232.13 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 116.365 232.9 116.735 ;
      VIA 232.13 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 109.725 232.92 110.055 ;
      VIA 232.13 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 109.705 232.9 110.075 ;
      VIA 232.13 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 103.065 232.92 103.395 ;
      VIA 232.13 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 103.045 232.9 103.415 ;
      VIA 232.13 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 96.405 232.92 96.735 ;
      VIA 232.13 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 96.385 232.9 96.755 ;
      VIA 232.13 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 89.745 232.92 90.075 ;
      VIA 232.13 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 89.725 232.9 90.095 ;
      VIA 232.13 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 83.085 232.92 83.415 ;
      VIA 232.13 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 83.065 232.9 83.435 ;
      VIA 232.13 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 76.425 232.92 76.755 ;
      VIA 232.13 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 76.405 232.9 76.775 ;
      VIA 232.13 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 69.765 232.92 70.095 ;
      VIA 232.13 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 69.745 232.9 70.115 ;
      VIA 232.13 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 63.105 232.92 63.435 ;
      VIA 232.13 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 63.085 232.9 63.455 ;
      VIA 232.13 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 56.445 232.92 56.775 ;
      VIA 232.13 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 56.425 232.9 56.795 ;
      VIA 232.13 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 49.785 232.92 50.115 ;
      VIA 232.13 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 49.765 232.9 50.135 ;
      VIA 232.13 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 43.125 232.92 43.455 ;
      VIA 232.13 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 43.105 232.9 43.475 ;
      VIA 232.13 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 36.465 232.92 36.795 ;
      VIA 232.13 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 36.445 232.9 36.815 ;
      VIA 232.13 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 29.805 232.92 30.135 ;
      VIA 232.13 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 29.785 232.9 30.155 ;
      VIA 232.13 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 23.145 232.92 23.475 ;
      VIA 232.13 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 23.125 232.9 23.495 ;
      VIA 232.13 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 16.485 232.92 16.815 ;
      VIA 232.13 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 16.465 232.9 16.835 ;
      VIA 232.13 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 9.825 232.92 10.155 ;
      VIA 232.13 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 9.805 232.9 10.175 ;
      VIA 232.13 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  231.34 3.165 232.92 3.495 ;
      VIA 232.13 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  231.36 3.145 232.9 3.515 ;
      VIA 232.13 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 232.13 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 775.725 205.78 776.055 ;
      VIA 204.99 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 775.705 205.76 776.075 ;
      VIA 204.99 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 769.065 205.78 769.395 ;
      VIA 204.99 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 769.045 205.76 769.415 ;
      VIA 204.99 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 762.405 205.78 762.735 ;
      VIA 204.99 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 762.385 205.76 762.755 ;
      VIA 204.99 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 755.745 205.78 756.075 ;
      VIA 204.99 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 755.725 205.76 756.095 ;
      VIA 204.99 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 749.085 205.78 749.415 ;
      VIA 204.99 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 749.065 205.76 749.435 ;
      VIA 204.99 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 742.425 205.78 742.755 ;
      VIA 204.99 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 742.405 205.76 742.775 ;
      VIA 204.99 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 735.765 205.78 736.095 ;
      VIA 204.99 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 735.745 205.76 736.115 ;
      VIA 204.99 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 729.105 205.78 729.435 ;
      VIA 204.99 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 729.085 205.76 729.455 ;
      VIA 204.99 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 722.445 205.78 722.775 ;
      VIA 204.99 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 722.425 205.76 722.795 ;
      VIA 204.99 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 715.785 205.78 716.115 ;
      VIA 204.99 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 715.765 205.76 716.135 ;
      VIA 204.99 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 709.125 205.78 709.455 ;
      VIA 204.99 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 709.105 205.76 709.475 ;
      VIA 204.99 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 702.465 205.78 702.795 ;
      VIA 204.99 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 702.445 205.76 702.815 ;
      VIA 204.99 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 695.805 205.78 696.135 ;
      VIA 204.99 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 695.785 205.76 696.155 ;
      VIA 204.99 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 689.145 205.78 689.475 ;
      VIA 204.99 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 689.125 205.76 689.495 ;
      VIA 204.99 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 682.485 205.78 682.815 ;
      VIA 204.99 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 682.465 205.76 682.835 ;
      VIA 204.99 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 675.825 205.78 676.155 ;
      VIA 204.99 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 675.805 205.76 676.175 ;
      VIA 204.99 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 669.165 205.78 669.495 ;
      VIA 204.99 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 669.145 205.76 669.515 ;
      VIA 204.99 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 662.505 205.78 662.835 ;
      VIA 204.99 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 662.485 205.76 662.855 ;
      VIA 204.99 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 655.845 205.78 656.175 ;
      VIA 204.99 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 655.825 205.76 656.195 ;
      VIA 204.99 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 649.185 205.78 649.515 ;
      VIA 204.99 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 649.165 205.76 649.535 ;
      VIA 204.99 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 642.525 205.78 642.855 ;
      VIA 204.99 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 642.505 205.76 642.875 ;
      VIA 204.99 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 635.865 205.78 636.195 ;
      VIA 204.99 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 635.845 205.76 636.215 ;
      VIA 204.99 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 629.205 205.78 629.535 ;
      VIA 204.99 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 629.185 205.76 629.555 ;
      VIA 204.99 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 622.545 205.78 622.875 ;
      VIA 204.99 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 622.525 205.76 622.895 ;
      VIA 204.99 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 615.885 205.78 616.215 ;
      VIA 204.99 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 615.865 205.76 616.235 ;
      VIA 204.99 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 609.225 205.78 609.555 ;
      VIA 204.99 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 609.205 205.76 609.575 ;
      VIA 204.99 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 602.565 205.78 602.895 ;
      VIA 204.99 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 602.545 205.76 602.915 ;
      VIA 204.99 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 595.905 205.78 596.235 ;
      VIA 204.99 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 595.885 205.76 596.255 ;
      VIA 204.99 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 589.245 205.78 589.575 ;
      VIA 204.99 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 589.225 205.76 589.595 ;
      VIA 204.99 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 582.585 205.78 582.915 ;
      VIA 204.99 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 582.565 205.76 582.935 ;
      VIA 204.99 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 575.925 205.78 576.255 ;
      VIA 204.99 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 575.905 205.76 576.275 ;
      VIA 204.99 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 569.265 205.78 569.595 ;
      VIA 204.99 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 569.245 205.76 569.615 ;
      VIA 204.99 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 562.605 205.78 562.935 ;
      VIA 204.99 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 562.585 205.76 562.955 ;
      VIA 204.99 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 555.945 205.78 556.275 ;
      VIA 204.99 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 555.925 205.76 556.295 ;
      VIA 204.99 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 549.285 205.78 549.615 ;
      VIA 204.99 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 549.265 205.76 549.635 ;
      VIA 204.99 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 542.625 205.78 542.955 ;
      VIA 204.99 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 542.605 205.76 542.975 ;
      VIA 204.99 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 535.965 205.78 536.295 ;
      VIA 204.99 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 535.945 205.76 536.315 ;
      VIA 204.99 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 529.305 205.78 529.635 ;
      VIA 204.99 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 529.285 205.76 529.655 ;
      VIA 204.99 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 522.645 205.78 522.975 ;
      VIA 204.99 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 522.625 205.76 522.995 ;
      VIA 204.99 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 515.985 205.78 516.315 ;
      VIA 204.99 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 515.965 205.76 516.335 ;
      VIA 204.99 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 509.325 205.78 509.655 ;
      VIA 204.99 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 509.305 205.76 509.675 ;
      VIA 204.99 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 502.665 205.78 502.995 ;
      VIA 204.99 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 502.645 205.76 503.015 ;
      VIA 204.99 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 496.005 205.78 496.335 ;
      VIA 204.99 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 495.985 205.76 496.355 ;
      VIA 204.99 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 489.345 205.78 489.675 ;
      VIA 204.99 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 489.325 205.76 489.695 ;
      VIA 204.99 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 482.685 205.78 483.015 ;
      VIA 204.99 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 482.665 205.76 483.035 ;
      VIA 204.99 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 476.025 205.78 476.355 ;
      VIA 204.99 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 476.005 205.76 476.375 ;
      VIA 204.99 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 469.365 205.78 469.695 ;
      VIA 204.99 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 469.345 205.76 469.715 ;
      VIA 204.99 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 462.705 205.78 463.035 ;
      VIA 204.99 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 462.685 205.76 463.055 ;
      VIA 204.99 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 456.045 205.78 456.375 ;
      VIA 204.99 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 456.025 205.76 456.395 ;
      VIA 204.99 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 449.385 205.78 449.715 ;
      VIA 204.99 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 449.365 205.76 449.735 ;
      VIA 204.99 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 442.725 205.78 443.055 ;
      VIA 204.99 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 442.705 205.76 443.075 ;
      VIA 204.99 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 436.065 205.78 436.395 ;
      VIA 204.99 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 436.045 205.76 436.415 ;
      VIA 204.99 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 429.405 205.78 429.735 ;
      VIA 204.99 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 429.385 205.76 429.755 ;
      VIA 204.99 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 422.745 205.78 423.075 ;
      VIA 204.99 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 422.725 205.76 423.095 ;
      VIA 204.99 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 416.085 205.78 416.415 ;
      VIA 204.99 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 416.065 205.76 416.435 ;
      VIA 204.99 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 409.425 205.78 409.755 ;
      VIA 204.99 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 409.405 205.76 409.775 ;
      VIA 204.99 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 402.765 205.78 403.095 ;
      VIA 204.99 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 402.745 205.76 403.115 ;
      VIA 204.99 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 396.105 205.78 396.435 ;
      VIA 204.99 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 396.085 205.76 396.455 ;
      VIA 204.99 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 389.445 205.78 389.775 ;
      VIA 204.99 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 389.425 205.76 389.795 ;
      VIA 204.99 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 382.785 205.78 383.115 ;
      VIA 204.99 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 382.765 205.76 383.135 ;
      VIA 204.99 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 376.125 205.78 376.455 ;
      VIA 204.99 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 376.105 205.76 376.475 ;
      VIA 204.99 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 369.465 205.78 369.795 ;
      VIA 204.99 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 369.445 205.76 369.815 ;
      VIA 204.99 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 362.805 205.78 363.135 ;
      VIA 204.99 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 362.785 205.76 363.155 ;
      VIA 204.99 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 356.145 205.78 356.475 ;
      VIA 204.99 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 356.125 205.76 356.495 ;
      VIA 204.99 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 349.485 205.78 349.815 ;
      VIA 204.99 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 349.465 205.76 349.835 ;
      VIA 204.99 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 342.825 205.78 343.155 ;
      VIA 204.99 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 342.805 205.76 343.175 ;
      VIA 204.99 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 336.165 205.78 336.495 ;
      VIA 204.99 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 336.145 205.76 336.515 ;
      VIA 204.99 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 329.505 205.78 329.835 ;
      VIA 204.99 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 329.485 205.76 329.855 ;
      VIA 204.99 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 322.845 205.78 323.175 ;
      VIA 204.99 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 322.825 205.76 323.195 ;
      VIA 204.99 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 316.185 205.78 316.515 ;
      VIA 204.99 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 316.165 205.76 316.535 ;
      VIA 204.99 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 309.525 205.78 309.855 ;
      VIA 204.99 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 309.505 205.76 309.875 ;
      VIA 204.99 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 302.865 205.78 303.195 ;
      VIA 204.99 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 302.845 205.76 303.215 ;
      VIA 204.99 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 296.205 205.78 296.535 ;
      VIA 204.99 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 296.185 205.76 296.555 ;
      VIA 204.99 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 289.545 205.78 289.875 ;
      VIA 204.99 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 289.525 205.76 289.895 ;
      VIA 204.99 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 282.885 205.78 283.215 ;
      VIA 204.99 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 282.865 205.76 283.235 ;
      VIA 204.99 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 276.225 205.78 276.555 ;
      VIA 204.99 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 276.205 205.76 276.575 ;
      VIA 204.99 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 269.565 205.78 269.895 ;
      VIA 204.99 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 269.545 205.76 269.915 ;
      VIA 204.99 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 262.905 205.78 263.235 ;
      VIA 204.99 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 262.885 205.76 263.255 ;
      VIA 204.99 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 256.245 205.78 256.575 ;
      VIA 204.99 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 256.225 205.76 256.595 ;
      VIA 204.99 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 249.585 205.78 249.915 ;
      VIA 204.99 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 249.565 205.76 249.935 ;
      VIA 204.99 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 242.925 205.78 243.255 ;
      VIA 204.99 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 242.905 205.76 243.275 ;
      VIA 204.99 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 236.265 205.78 236.595 ;
      VIA 204.99 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 236.245 205.76 236.615 ;
      VIA 204.99 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 229.605 205.78 229.935 ;
      VIA 204.99 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 229.585 205.76 229.955 ;
      VIA 204.99 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 222.945 205.78 223.275 ;
      VIA 204.99 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 222.925 205.76 223.295 ;
      VIA 204.99 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 216.285 205.78 216.615 ;
      VIA 204.99 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 216.265 205.76 216.635 ;
      VIA 204.99 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 209.625 205.78 209.955 ;
      VIA 204.99 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 209.605 205.76 209.975 ;
      VIA 204.99 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 202.965 205.78 203.295 ;
      VIA 204.99 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 202.945 205.76 203.315 ;
      VIA 204.99 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 196.305 205.78 196.635 ;
      VIA 204.99 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 196.285 205.76 196.655 ;
      VIA 204.99 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 189.645 205.78 189.975 ;
      VIA 204.99 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 189.625 205.76 189.995 ;
      VIA 204.99 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 182.985 205.78 183.315 ;
      VIA 204.99 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 182.965 205.76 183.335 ;
      VIA 204.99 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 176.325 205.78 176.655 ;
      VIA 204.99 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 176.305 205.76 176.675 ;
      VIA 204.99 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 169.665 205.78 169.995 ;
      VIA 204.99 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 169.645 205.76 170.015 ;
      VIA 204.99 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 163.005 205.78 163.335 ;
      VIA 204.99 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 162.985 205.76 163.355 ;
      VIA 204.99 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 156.345 205.78 156.675 ;
      VIA 204.99 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 156.325 205.76 156.695 ;
      VIA 204.99 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 149.685 205.78 150.015 ;
      VIA 204.99 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 149.665 205.76 150.035 ;
      VIA 204.99 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 143.025 205.78 143.355 ;
      VIA 204.99 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 143.005 205.76 143.375 ;
      VIA 204.99 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 136.365 205.78 136.695 ;
      VIA 204.99 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 136.345 205.76 136.715 ;
      VIA 204.99 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 129.705 205.78 130.035 ;
      VIA 204.99 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 129.685 205.76 130.055 ;
      VIA 204.99 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 123.045 205.78 123.375 ;
      VIA 204.99 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 123.025 205.76 123.395 ;
      VIA 204.99 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 116.385 205.78 116.715 ;
      VIA 204.99 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 116.365 205.76 116.735 ;
      VIA 204.99 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 109.725 205.78 110.055 ;
      VIA 204.99 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 109.705 205.76 110.075 ;
      VIA 204.99 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 103.065 205.78 103.395 ;
      VIA 204.99 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 103.045 205.76 103.415 ;
      VIA 204.99 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 96.405 205.78 96.735 ;
      VIA 204.99 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 96.385 205.76 96.755 ;
      VIA 204.99 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 89.745 205.78 90.075 ;
      VIA 204.99 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 89.725 205.76 90.095 ;
      VIA 204.99 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 83.085 205.78 83.415 ;
      VIA 204.99 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 83.065 205.76 83.435 ;
      VIA 204.99 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 76.425 205.78 76.755 ;
      VIA 204.99 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 76.405 205.76 76.775 ;
      VIA 204.99 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 69.765 205.78 70.095 ;
      VIA 204.99 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 69.745 205.76 70.115 ;
      VIA 204.99 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 63.105 205.78 63.435 ;
      VIA 204.99 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 63.085 205.76 63.455 ;
      VIA 204.99 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 56.445 205.78 56.775 ;
      VIA 204.99 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 56.425 205.76 56.795 ;
      VIA 204.99 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 49.785 205.78 50.115 ;
      VIA 204.99 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 49.765 205.76 50.135 ;
      VIA 204.99 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 43.125 205.78 43.455 ;
      VIA 204.99 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 43.105 205.76 43.475 ;
      VIA 204.99 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 36.465 205.78 36.795 ;
      VIA 204.99 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 36.445 205.76 36.815 ;
      VIA 204.99 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 29.805 205.78 30.135 ;
      VIA 204.99 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 29.785 205.76 30.155 ;
      VIA 204.99 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 23.145 205.78 23.475 ;
      VIA 204.99 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 23.125 205.76 23.495 ;
      VIA 204.99 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 16.485 205.78 16.815 ;
      VIA 204.99 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 16.465 205.76 16.835 ;
      VIA 204.99 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 9.825 205.78 10.155 ;
      VIA 204.99 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 9.805 205.76 10.175 ;
      VIA 204.99 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  204.2 3.165 205.78 3.495 ;
      VIA 204.99 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  204.22 3.145 205.76 3.515 ;
      VIA 204.99 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 204.99 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 775.725 178.64 776.055 ;
      VIA 177.85 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 775.705 178.62 776.075 ;
      VIA 177.85 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 769.065 178.64 769.395 ;
      VIA 177.85 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 769.045 178.62 769.415 ;
      VIA 177.85 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 762.405 178.64 762.735 ;
      VIA 177.85 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 762.385 178.62 762.755 ;
      VIA 177.85 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 755.745 178.64 756.075 ;
      VIA 177.85 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 755.725 178.62 756.095 ;
      VIA 177.85 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 749.085 178.64 749.415 ;
      VIA 177.85 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 749.065 178.62 749.435 ;
      VIA 177.85 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 742.425 178.64 742.755 ;
      VIA 177.85 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 742.405 178.62 742.775 ;
      VIA 177.85 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 735.765 178.64 736.095 ;
      VIA 177.85 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 735.745 178.62 736.115 ;
      VIA 177.85 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 729.105 178.64 729.435 ;
      VIA 177.85 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 729.085 178.62 729.455 ;
      VIA 177.85 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 722.445 178.64 722.775 ;
      VIA 177.85 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 722.425 178.62 722.795 ;
      VIA 177.85 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 715.785 178.64 716.115 ;
      VIA 177.85 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 715.765 178.62 716.135 ;
      VIA 177.85 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 709.125 178.64 709.455 ;
      VIA 177.85 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 709.105 178.62 709.475 ;
      VIA 177.85 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 702.465 178.64 702.795 ;
      VIA 177.85 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 702.445 178.62 702.815 ;
      VIA 177.85 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 695.805 178.64 696.135 ;
      VIA 177.85 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 695.785 178.62 696.155 ;
      VIA 177.85 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 689.145 178.64 689.475 ;
      VIA 177.85 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 689.125 178.62 689.495 ;
      VIA 177.85 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 682.485 178.64 682.815 ;
      VIA 177.85 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 682.465 178.62 682.835 ;
      VIA 177.85 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 675.825 178.64 676.155 ;
      VIA 177.85 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 675.805 178.62 676.175 ;
      VIA 177.85 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 669.165 178.64 669.495 ;
      VIA 177.85 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 669.145 178.62 669.515 ;
      VIA 177.85 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 662.505 178.64 662.835 ;
      VIA 177.85 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 662.485 178.62 662.855 ;
      VIA 177.85 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 655.845 178.64 656.175 ;
      VIA 177.85 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 655.825 178.62 656.195 ;
      VIA 177.85 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 649.185 178.64 649.515 ;
      VIA 177.85 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 649.165 178.62 649.535 ;
      VIA 177.85 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 642.525 178.64 642.855 ;
      VIA 177.85 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 642.505 178.62 642.875 ;
      VIA 177.85 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 635.865 178.64 636.195 ;
      VIA 177.85 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 635.845 178.62 636.215 ;
      VIA 177.85 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 629.205 178.64 629.535 ;
      VIA 177.85 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 629.185 178.62 629.555 ;
      VIA 177.85 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 622.545 178.64 622.875 ;
      VIA 177.85 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 622.525 178.62 622.895 ;
      VIA 177.85 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 615.885 178.64 616.215 ;
      VIA 177.85 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 615.865 178.62 616.235 ;
      VIA 177.85 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 609.225 178.64 609.555 ;
      VIA 177.85 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 609.205 178.62 609.575 ;
      VIA 177.85 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 602.565 178.64 602.895 ;
      VIA 177.85 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 602.545 178.62 602.915 ;
      VIA 177.85 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 595.905 178.64 596.235 ;
      VIA 177.85 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 595.885 178.62 596.255 ;
      VIA 177.85 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 589.245 178.64 589.575 ;
      VIA 177.85 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 589.225 178.62 589.595 ;
      VIA 177.85 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 582.585 178.64 582.915 ;
      VIA 177.85 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 582.565 178.62 582.935 ;
      VIA 177.85 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 575.925 178.64 576.255 ;
      VIA 177.85 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 575.905 178.62 576.275 ;
      VIA 177.85 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 569.265 178.64 569.595 ;
      VIA 177.85 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 569.245 178.62 569.615 ;
      VIA 177.85 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 562.605 178.64 562.935 ;
      VIA 177.85 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 562.585 178.62 562.955 ;
      VIA 177.85 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 555.945 178.64 556.275 ;
      VIA 177.85 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 555.925 178.62 556.295 ;
      VIA 177.85 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 549.285 178.64 549.615 ;
      VIA 177.85 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 549.265 178.62 549.635 ;
      VIA 177.85 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 542.625 178.64 542.955 ;
      VIA 177.85 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 542.605 178.62 542.975 ;
      VIA 177.85 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 535.965 178.64 536.295 ;
      VIA 177.85 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 535.945 178.62 536.315 ;
      VIA 177.85 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 529.305 178.64 529.635 ;
      VIA 177.85 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 529.285 178.62 529.655 ;
      VIA 177.85 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 522.645 178.64 522.975 ;
      VIA 177.85 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 522.625 178.62 522.995 ;
      VIA 177.85 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 515.985 178.64 516.315 ;
      VIA 177.85 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 515.965 178.62 516.335 ;
      VIA 177.85 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 509.325 178.64 509.655 ;
      VIA 177.85 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 509.305 178.62 509.675 ;
      VIA 177.85 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 502.665 178.64 502.995 ;
      VIA 177.85 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 502.645 178.62 503.015 ;
      VIA 177.85 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 496.005 178.64 496.335 ;
      VIA 177.85 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 495.985 178.62 496.355 ;
      VIA 177.85 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 489.345 178.64 489.675 ;
      VIA 177.85 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 489.325 178.62 489.695 ;
      VIA 177.85 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 482.685 178.64 483.015 ;
      VIA 177.85 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 482.665 178.62 483.035 ;
      VIA 177.85 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 476.025 178.64 476.355 ;
      VIA 177.85 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 476.005 178.62 476.375 ;
      VIA 177.85 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 469.365 178.64 469.695 ;
      VIA 177.85 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 469.345 178.62 469.715 ;
      VIA 177.85 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 462.705 178.64 463.035 ;
      VIA 177.85 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 462.685 178.62 463.055 ;
      VIA 177.85 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 456.045 178.64 456.375 ;
      VIA 177.85 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 456.025 178.62 456.395 ;
      VIA 177.85 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 449.385 178.64 449.715 ;
      VIA 177.85 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 449.365 178.62 449.735 ;
      VIA 177.85 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 442.725 178.64 443.055 ;
      VIA 177.85 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 442.705 178.62 443.075 ;
      VIA 177.85 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 436.065 178.64 436.395 ;
      VIA 177.85 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 436.045 178.62 436.415 ;
      VIA 177.85 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 429.405 178.64 429.735 ;
      VIA 177.85 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 429.385 178.62 429.755 ;
      VIA 177.85 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 422.745 178.64 423.075 ;
      VIA 177.85 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 422.725 178.62 423.095 ;
      VIA 177.85 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 416.085 178.64 416.415 ;
      VIA 177.85 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 416.065 178.62 416.435 ;
      VIA 177.85 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 409.425 178.64 409.755 ;
      VIA 177.85 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 409.405 178.62 409.775 ;
      VIA 177.85 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 402.765 178.64 403.095 ;
      VIA 177.85 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 402.745 178.62 403.115 ;
      VIA 177.85 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 396.105 178.64 396.435 ;
      VIA 177.85 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 396.085 178.62 396.455 ;
      VIA 177.85 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 389.445 178.64 389.775 ;
      VIA 177.85 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 389.425 178.62 389.795 ;
      VIA 177.85 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 382.785 178.64 383.115 ;
      VIA 177.85 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 382.765 178.62 383.135 ;
      VIA 177.85 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 376.125 178.64 376.455 ;
      VIA 177.85 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 376.105 178.62 376.475 ;
      VIA 177.85 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 369.465 178.64 369.795 ;
      VIA 177.85 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 369.445 178.62 369.815 ;
      VIA 177.85 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 362.805 178.64 363.135 ;
      VIA 177.85 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 362.785 178.62 363.155 ;
      VIA 177.85 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 356.145 178.64 356.475 ;
      VIA 177.85 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 356.125 178.62 356.495 ;
      VIA 177.85 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 349.485 178.64 349.815 ;
      VIA 177.85 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 349.465 178.62 349.835 ;
      VIA 177.85 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 342.825 178.64 343.155 ;
      VIA 177.85 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 342.805 178.62 343.175 ;
      VIA 177.85 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 336.165 178.64 336.495 ;
      VIA 177.85 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 336.145 178.62 336.515 ;
      VIA 177.85 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 329.505 178.64 329.835 ;
      VIA 177.85 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 329.485 178.62 329.855 ;
      VIA 177.85 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 322.845 178.64 323.175 ;
      VIA 177.85 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 322.825 178.62 323.195 ;
      VIA 177.85 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 316.185 178.64 316.515 ;
      VIA 177.85 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 316.165 178.62 316.535 ;
      VIA 177.85 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 309.525 178.64 309.855 ;
      VIA 177.85 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 309.505 178.62 309.875 ;
      VIA 177.85 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 302.865 178.64 303.195 ;
      VIA 177.85 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 302.845 178.62 303.215 ;
      VIA 177.85 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 296.205 178.64 296.535 ;
      VIA 177.85 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 296.185 178.62 296.555 ;
      VIA 177.85 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 289.545 178.64 289.875 ;
      VIA 177.85 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 289.525 178.62 289.895 ;
      VIA 177.85 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 282.885 178.64 283.215 ;
      VIA 177.85 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 282.865 178.62 283.235 ;
      VIA 177.85 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 276.225 178.64 276.555 ;
      VIA 177.85 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 276.205 178.62 276.575 ;
      VIA 177.85 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 269.565 178.64 269.895 ;
      VIA 177.85 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 269.545 178.62 269.915 ;
      VIA 177.85 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 262.905 178.64 263.235 ;
      VIA 177.85 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 262.885 178.62 263.255 ;
      VIA 177.85 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 256.245 178.64 256.575 ;
      VIA 177.85 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 256.225 178.62 256.595 ;
      VIA 177.85 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 249.585 178.64 249.915 ;
      VIA 177.85 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 249.565 178.62 249.935 ;
      VIA 177.85 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 242.925 178.64 243.255 ;
      VIA 177.85 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 242.905 178.62 243.275 ;
      VIA 177.85 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 236.265 178.64 236.595 ;
      VIA 177.85 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 236.245 178.62 236.615 ;
      VIA 177.85 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 229.605 178.64 229.935 ;
      VIA 177.85 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 229.585 178.62 229.955 ;
      VIA 177.85 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 222.945 178.64 223.275 ;
      VIA 177.85 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 222.925 178.62 223.295 ;
      VIA 177.85 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 216.285 178.64 216.615 ;
      VIA 177.85 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 216.265 178.62 216.635 ;
      VIA 177.85 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 209.625 178.64 209.955 ;
      VIA 177.85 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 209.605 178.62 209.975 ;
      VIA 177.85 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 202.965 178.64 203.295 ;
      VIA 177.85 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 202.945 178.62 203.315 ;
      VIA 177.85 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 196.305 178.64 196.635 ;
      VIA 177.85 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 196.285 178.62 196.655 ;
      VIA 177.85 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 189.645 178.64 189.975 ;
      VIA 177.85 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 189.625 178.62 189.995 ;
      VIA 177.85 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 182.985 178.64 183.315 ;
      VIA 177.85 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 182.965 178.62 183.335 ;
      VIA 177.85 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 176.325 178.64 176.655 ;
      VIA 177.85 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 176.305 178.62 176.675 ;
      VIA 177.85 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 169.665 178.64 169.995 ;
      VIA 177.85 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 169.645 178.62 170.015 ;
      VIA 177.85 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 163.005 178.64 163.335 ;
      VIA 177.85 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 162.985 178.62 163.355 ;
      VIA 177.85 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 156.345 178.64 156.675 ;
      VIA 177.85 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 156.325 178.62 156.695 ;
      VIA 177.85 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 149.685 178.64 150.015 ;
      VIA 177.85 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 149.665 178.62 150.035 ;
      VIA 177.85 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 143.025 178.64 143.355 ;
      VIA 177.85 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 143.005 178.62 143.375 ;
      VIA 177.85 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 136.365 178.64 136.695 ;
      VIA 177.85 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 136.345 178.62 136.715 ;
      VIA 177.85 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 129.705 178.64 130.035 ;
      VIA 177.85 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 129.685 178.62 130.055 ;
      VIA 177.85 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 123.045 178.64 123.375 ;
      VIA 177.85 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 123.025 178.62 123.395 ;
      VIA 177.85 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 116.385 178.64 116.715 ;
      VIA 177.85 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 116.365 178.62 116.735 ;
      VIA 177.85 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 109.725 178.64 110.055 ;
      VIA 177.85 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 109.705 178.62 110.075 ;
      VIA 177.85 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 103.065 178.64 103.395 ;
      VIA 177.85 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 103.045 178.62 103.415 ;
      VIA 177.85 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 96.405 178.64 96.735 ;
      VIA 177.85 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 96.385 178.62 96.755 ;
      VIA 177.85 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 89.745 178.64 90.075 ;
      VIA 177.85 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 89.725 178.62 90.095 ;
      VIA 177.85 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 83.085 178.64 83.415 ;
      VIA 177.85 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 83.065 178.62 83.435 ;
      VIA 177.85 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 76.425 178.64 76.755 ;
      VIA 177.85 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 76.405 178.62 76.775 ;
      VIA 177.85 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 69.765 178.64 70.095 ;
      VIA 177.85 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 69.745 178.62 70.115 ;
      VIA 177.85 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 63.105 178.64 63.435 ;
      VIA 177.85 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 63.085 178.62 63.455 ;
      VIA 177.85 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 56.445 178.64 56.775 ;
      VIA 177.85 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 56.425 178.62 56.795 ;
      VIA 177.85 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 49.785 178.64 50.115 ;
      VIA 177.85 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 49.765 178.62 50.135 ;
      VIA 177.85 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 43.125 178.64 43.455 ;
      VIA 177.85 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 43.105 178.62 43.475 ;
      VIA 177.85 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 36.465 178.64 36.795 ;
      VIA 177.85 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 36.445 178.62 36.815 ;
      VIA 177.85 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 29.805 178.64 30.135 ;
      VIA 177.85 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 29.785 178.62 30.155 ;
      VIA 177.85 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 23.145 178.64 23.475 ;
      VIA 177.85 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 23.125 178.62 23.495 ;
      VIA 177.85 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 16.485 178.64 16.815 ;
      VIA 177.85 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 16.465 178.62 16.835 ;
      VIA 177.85 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 9.825 178.64 10.155 ;
      VIA 177.85 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 9.805 178.62 10.175 ;
      VIA 177.85 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  177.06 3.165 178.64 3.495 ;
      VIA 177.85 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  177.08 3.145 178.62 3.515 ;
      VIA 177.85 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 177.85 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 775.725 151.5 776.055 ;
      VIA 150.71 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 775.705 151.48 776.075 ;
      VIA 150.71 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 769.065 151.5 769.395 ;
      VIA 150.71 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 769.045 151.48 769.415 ;
      VIA 150.71 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 762.405 151.5 762.735 ;
      VIA 150.71 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 762.385 151.48 762.755 ;
      VIA 150.71 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 755.745 151.5 756.075 ;
      VIA 150.71 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 755.725 151.48 756.095 ;
      VIA 150.71 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 749.085 151.5 749.415 ;
      VIA 150.71 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 749.065 151.48 749.435 ;
      VIA 150.71 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 742.425 151.5 742.755 ;
      VIA 150.71 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 742.405 151.48 742.775 ;
      VIA 150.71 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 735.765 151.5 736.095 ;
      VIA 150.71 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 735.745 151.48 736.115 ;
      VIA 150.71 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 729.105 151.5 729.435 ;
      VIA 150.71 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 729.085 151.48 729.455 ;
      VIA 150.71 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 722.445 151.5 722.775 ;
      VIA 150.71 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 722.425 151.48 722.795 ;
      VIA 150.71 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 715.785 151.5 716.115 ;
      VIA 150.71 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 715.765 151.48 716.135 ;
      VIA 150.71 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 709.125 151.5 709.455 ;
      VIA 150.71 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 709.105 151.48 709.475 ;
      VIA 150.71 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 702.465 151.5 702.795 ;
      VIA 150.71 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 702.445 151.48 702.815 ;
      VIA 150.71 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 695.805 151.5 696.135 ;
      VIA 150.71 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 695.785 151.48 696.155 ;
      VIA 150.71 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 689.145 151.5 689.475 ;
      VIA 150.71 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 689.125 151.48 689.495 ;
      VIA 150.71 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 682.485 151.5 682.815 ;
      VIA 150.71 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 682.465 151.48 682.835 ;
      VIA 150.71 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 675.825 151.5 676.155 ;
      VIA 150.71 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 675.805 151.48 676.175 ;
      VIA 150.71 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 669.165 151.5 669.495 ;
      VIA 150.71 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 669.145 151.48 669.515 ;
      VIA 150.71 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 662.505 151.5 662.835 ;
      VIA 150.71 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 662.485 151.48 662.855 ;
      VIA 150.71 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 655.845 151.5 656.175 ;
      VIA 150.71 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 655.825 151.48 656.195 ;
      VIA 150.71 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 649.185 151.5 649.515 ;
      VIA 150.71 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 649.165 151.48 649.535 ;
      VIA 150.71 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 642.525 151.5 642.855 ;
      VIA 150.71 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 642.505 151.48 642.875 ;
      VIA 150.71 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 635.865 151.5 636.195 ;
      VIA 150.71 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 635.845 151.48 636.215 ;
      VIA 150.71 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 629.205 151.5 629.535 ;
      VIA 150.71 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 629.185 151.48 629.555 ;
      VIA 150.71 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 622.545 151.5 622.875 ;
      VIA 150.71 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 622.525 151.48 622.895 ;
      VIA 150.71 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 615.885 151.5 616.215 ;
      VIA 150.71 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 615.865 151.48 616.235 ;
      VIA 150.71 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 609.225 151.5 609.555 ;
      VIA 150.71 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 609.205 151.48 609.575 ;
      VIA 150.71 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 602.565 151.5 602.895 ;
      VIA 150.71 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 602.545 151.48 602.915 ;
      VIA 150.71 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 595.905 151.5 596.235 ;
      VIA 150.71 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 595.885 151.48 596.255 ;
      VIA 150.71 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 589.245 151.5 589.575 ;
      VIA 150.71 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 589.225 151.48 589.595 ;
      VIA 150.71 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 582.585 151.5 582.915 ;
      VIA 150.71 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 582.565 151.48 582.935 ;
      VIA 150.71 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 575.925 151.5 576.255 ;
      VIA 150.71 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 575.905 151.48 576.275 ;
      VIA 150.71 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 569.265 151.5 569.595 ;
      VIA 150.71 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 569.245 151.48 569.615 ;
      VIA 150.71 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 562.605 151.5 562.935 ;
      VIA 150.71 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 562.585 151.48 562.955 ;
      VIA 150.71 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 555.945 151.5 556.275 ;
      VIA 150.71 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 555.925 151.48 556.295 ;
      VIA 150.71 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 549.285 151.5 549.615 ;
      VIA 150.71 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 549.265 151.48 549.635 ;
      VIA 150.71 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 542.625 151.5 542.955 ;
      VIA 150.71 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 542.605 151.48 542.975 ;
      VIA 150.71 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 535.965 151.5 536.295 ;
      VIA 150.71 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 535.945 151.48 536.315 ;
      VIA 150.71 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 529.305 151.5 529.635 ;
      VIA 150.71 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 529.285 151.48 529.655 ;
      VIA 150.71 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 522.645 151.5 522.975 ;
      VIA 150.71 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 522.625 151.48 522.995 ;
      VIA 150.71 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 515.985 151.5 516.315 ;
      VIA 150.71 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 515.965 151.48 516.335 ;
      VIA 150.71 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 509.325 151.5 509.655 ;
      VIA 150.71 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 509.305 151.48 509.675 ;
      VIA 150.71 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 502.665 151.5 502.995 ;
      VIA 150.71 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 502.645 151.48 503.015 ;
      VIA 150.71 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 496.005 151.5 496.335 ;
      VIA 150.71 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 495.985 151.48 496.355 ;
      VIA 150.71 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 489.345 151.5 489.675 ;
      VIA 150.71 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 489.325 151.48 489.695 ;
      VIA 150.71 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 482.685 151.5 483.015 ;
      VIA 150.71 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 482.665 151.48 483.035 ;
      VIA 150.71 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 476.025 151.5 476.355 ;
      VIA 150.71 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 476.005 151.48 476.375 ;
      VIA 150.71 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 469.365 151.5 469.695 ;
      VIA 150.71 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 469.345 151.48 469.715 ;
      VIA 150.71 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 462.705 151.5 463.035 ;
      VIA 150.71 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 462.685 151.48 463.055 ;
      VIA 150.71 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 456.045 151.5 456.375 ;
      VIA 150.71 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 456.025 151.48 456.395 ;
      VIA 150.71 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 449.385 151.5 449.715 ;
      VIA 150.71 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 449.365 151.48 449.735 ;
      VIA 150.71 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 442.725 151.5 443.055 ;
      VIA 150.71 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 442.705 151.48 443.075 ;
      VIA 150.71 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 436.065 151.5 436.395 ;
      VIA 150.71 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 436.045 151.48 436.415 ;
      VIA 150.71 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 429.405 151.5 429.735 ;
      VIA 150.71 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 429.385 151.48 429.755 ;
      VIA 150.71 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 422.745 151.5 423.075 ;
      VIA 150.71 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 422.725 151.48 423.095 ;
      VIA 150.71 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 416.085 151.5 416.415 ;
      VIA 150.71 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 416.065 151.48 416.435 ;
      VIA 150.71 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 409.425 151.5 409.755 ;
      VIA 150.71 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 409.405 151.48 409.775 ;
      VIA 150.71 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 402.765 151.5 403.095 ;
      VIA 150.71 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 402.745 151.48 403.115 ;
      VIA 150.71 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 396.105 151.5 396.435 ;
      VIA 150.71 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 396.085 151.48 396.455 ;
      VIA 150.71 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 389.445 151.5 389.775 ;
      VIA 150.71 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 389.425 151.48 389.795 ;
      VIA 150.71 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 382.785 151.5 383.115 ;
      VIA 150.71 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 382.765 151.48 383.135 ;
      VIA 150.71 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 376.125 151.5 376.455 ;
      VIA 150.71 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 376.105 151.48 376.475 ;
      VIA 150.71 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 369.465 151.5 369.795 ;
      VIA 150.71 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 369.445 151.48 369.815 ;
      VIA 150.71 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 362.805 151.5 363.135 ;
      VIA 150.71 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 362.785 151.48 363.155 ;
      VIA 150.71 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 356.145 151.5 356.475 ;
      VIA 150.71 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 356.125 151.48 356.495 ;
      VIA 150.71 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 349.485 151.5 349.815 ;
      VIA 150.71 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 349.465 151.48 349.835 ;
      VIA 150.71 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 342.825 151.5 343.155 ;
      VIA 150.71 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 342.805 151.48 343.175 ;
      VIA 150.71 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 336.165 151.5 336.495 ;
      VIA 150.71 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 336.145 151.48 336.515 ;
      VIA 150.71 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 329.505 151.5 329.835 ;
      VIA 150.71 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 329.485 151.48 329.855 ;
      VIA 150.71 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 322.845 151.5 323.175 ;
      VIA 150.71 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 322.825 151.48 323.195 ;
      VIA 150.71 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 316.185 151.5 316.515 ;
      VIA 150.71 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 316.165 151.48 316.535 ;
      VIA 150.71 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 309.525 151.5 309.855 ;
      VIA 150.71 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 309.505 151.48 309.875 ;
      VIA 150.71 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 302.865 151.5 303.195 ;
      VIA 150.71 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 302.845 151.48 303.215 ;
      VIA 150.71 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 296.205 151.5 296.535 ;
      VIA 150.71 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 296.185 151.48 296.555 ;
      VIA 150.71 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 289.545 151.5 289.875 ;
      VIA 150.71 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 289.525 151.48 289.895 ;
      VIA 150.71 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 282.885 151.5 283.215 ;
      VIA 150.71 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 282.865 151.48 283.235 ;
      VIA 150.71 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 276.225 151.5 276.555 ;
      VIA 150.71 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 276.205 151.48 276.575 ;
      VIA 150.71 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 269.565 151.5 269.895 ;
      VIA 150.71 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 269.545 151.48 269.915 ;
      VIA 150.71 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 262.905 151.5 263.235 ;
      VIA 150.71 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 262.885 151.48 263.255 ;
      VIA 150.71 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 256.245 151.5 256.575 ;
      VIA 150.71 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 256.225 151.48 256.595 ;
      VIA 150.71 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 249.585 151.5 249.915 ;
      VIA 150.71 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 249.565 151.48 249.935 ;
      VIA 150.71 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 242.925 151.5 243.255 ;
      VIA 150.71 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 242.905 151.48 243.275 ;
      VIA 150.71 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 236.265 151.5 236.595 ;
      VIA 150.71 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 236.245 151.48 236.615 ;
      VIA 150.71 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 229.605 151.5 229.935 ;
      VIA 150.71 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 229.585 151.48 229.955 ;
      VIA 150.71 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 222.945 151.5 223.275 ;
      VIA 150.71 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 222.925 151.48 223.295 ;
      VIA 150.71 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 216.285 151.5 216.615 ;
      VIA 150.71 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 216.265 151.48 216.635 ;
      VIA 150.71 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 209.625 151.5 209.955 ;
      VIA 150.71 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 209.605 151.48 209.975 ;
      VIA 150.71 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 202.965 151.5 203.295 ;
      VIA 150.71 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 202.945 151.48 203.315 ;
      VIA 150.71 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 196.305 151.5 196.635 ;
      VIA 150.71 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 196.285 151.48 196.655 ;
      VIA 150.71 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 189.645 151.5 189.975 ;
      VIA 150.71 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 189.625 151.48 189.995 ;
      VIA 150.71 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 182.985 151.5 183.315 ;
      VIA 150.71 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 182.965 151.48 183.335 ;
      VIA 150.71 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 176.325 151.5 176.655 ;
      VIA 150.71 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 176.305 151.48 176.675 ;
      VIA 150.71 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 169.665 151.5 169.995 ;
      VIA 150.71 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 169.645 151.48 170.015 ;
      VIA 150.71 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 163.005 151.5 163.335 ;
      VIA 150.71 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 162.985 151.48 163.355 ;
      VIA 150.71 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 156.345 151.5 156.675 ;
      VIA 150.71 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 156.325 151.48 156.695 ;
      VIA 150.71 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 149.685 151.5 150.015 ;
      VIA 150.71 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 149.665 151.48 150.035 ;
      VIA 150.71 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 143.025 151.5 143.355 ;
      VIA 150.71 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 143.005 151.48 143.375 ;
      VIA 150.71 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 136.365 151.5 136.695 ;
      VIA 150.71 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 136.345 151.48 136.715 ;
      VIA 150.71 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 129.705 151.5 130.035 ;
      VIA 150.71 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 129.685 151.48 130.055 ;
      VIA 150.71 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 123.045 151.5 123.375 ;
      VIA 150.71 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 123.025 151.48 123.395 ;
      VIA 150.71 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 116.385 151.5 116.715 ;
      VIA 150.71 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 116.365 151.48 116.735 ;
      VIA 150.71 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 109.725 151.5 110.055 ;
      VIA 150.71 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 109.705 151.48 110.075 ;
      VIA 150.71 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 103.065 151.5 103.395 ;
      VIA 150.71 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 103.045 151.48 103.415 ;
      VIA 150.71 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 96.405 151.5 96.735 ;
      VIA 150.71 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 96.385 151.48 96.755 ;
      VIA 150.71 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 89.745 151.5 90.075 ;
      VIA 150.71 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 89.725 151.48 90.095 ;
      VIA 150.71 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 83.085 151.5 83.415 ;
      VIA 150.71 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 83.065 151.48 83.435 ;
      VIA 150.71 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 76.425 151.5 76.755 ;
      VIA 150.71 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 76.405 151.48 76.775 ;
      VIA 150.71 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 69.765 151.5 70.095 ;
      VIA 150.71 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 69.745 151.48 70.115 ;
      VIA 150.71 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 63.105 151.5 63.435 ;
      VIA 150.71 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 63.085 151.48 63.455 ;
      VIA 150.71 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 56.445 151.5 56.775 ;
      VIA 150.71 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 56.425 151.48 56.795 ;
      VIA 150.71 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 49.785 151.5 50.115 ;
      VIA 150.71 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 49.765 151.48 50.135 ;
      VIA 150.71 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 43.125 151.5 43.455 ;
      VIA 150.71 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 43.105 151.48 43.475 ;
      VIA 150.71 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 36.465 151.5 36.795 ;
      VIA 150.71 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 36.445 151.48 36.815 ;
      VIA 150.71 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 29.805 151.5 30.135 ;
      VIA 150.71 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 29.785 151.48 30.155 ;
      VIA 150.71 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 23.145 151.5 23.475 ;
      VIA 150.71 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 23.125 151.48 23.495 ;
      VIA 150.71 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 16.485 151.5 16.815 ;
      VIA 150.71 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 16.465 151.48 16.835 ;
      VIA 150.71 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 9.825 151.5 10.155 ;
      VIA 150.71 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 9.805 151.48 10.175 ;
      VIA 150.71 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.92 3.165 151.5 3.495 ;
      VIA 150.71 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.94 3.145 151.48 3.515 ;
      VIA 150.71 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 150.71 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 775.725 124.36 776.055 ;
      VIA 123.57 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 775.705 124.34 776.075 ;
      VIA 123.57 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 769.065 124.36 769.395 ;
      VIA 123.57 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 769.045 124.34 769.415 ;
      VIA 123.57 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 762.405 124.36 762.735 ;
      VIA 123.57 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 762.385 124.34 762.755 ;
      VIA 123.57 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 755.745 124.36 756.075 ;
      VIA 123.57 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 755.725 124.34 756.095 ;
      VIA 123.57 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 749.085 124.36 749.415 ;
      VIA 123.57 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 749.065 124.34 749.435 ;
      VIA 123.57 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 742.425 124.36 742.755 ;
      VIA 123.57 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 742.405 124.34 742.775 ;
      VIA 123.57 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 735.765 124.36 736.095 ;
      VIA 123.57 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 735.745 124.34 736.115 ;
      VIA 123.57 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 729.105 124.36 729.435 ;
      VIA 123.57 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 729.085 124.34 729.455 ;
      VIA 123.57 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 722.445 124.36 722.775 ;
      VIA 123.57 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 722.425 124.34 722.795 ;
      VIA 123.57 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 715.785 124.36 716.115 ;
      VIA 123.57 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 715.765 124.34 716.135 ;
      VIA 123.57 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 709.125 124.36 709.455 ;
      VIA 123.57 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 709.105 124.34 709.475 ;
      VIA 123.57 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 702.465 124.36 702.795 ;
      VIA 123.57 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 702.445 124.34 702.815 ;
      VIA 123.57 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 695.805 124.36 696.135 ;
      VIA 123.57 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 695.785 124.34 696.155 ;
      VIA 123.57 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 689.145 124.36 689.475 ;
      VIA 123.57 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 689.125 124.34 689.495 ;
      VIA 123.57 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 682.485 124.36 682.815 ;
      VIA 123.57 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 682.465 124.34 682.835 ;
      VIA 123.57 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 675.825 124.36 676.155 ;
      VIA 123.57 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 675.805 124.34 676.175 ;
      VIA 123.57 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 669.165 124.36 669.495 ;
      VIA 123.57 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 669.145 124.34 669.515 ;
      VIA 123.57 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 662.505 124.36 662.835 ;
      VIA 123.57 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 662.485 124.34 662.855 ;
      VIA 123.57 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 655.845 124.36 656.175 ;
      VIA 123.57 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 655.825 124.34 656.195 ;
      VIA 123.57 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 649.185 124.36 649.515 ;
      VIA 123.57 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 649.165 124.34 649.535 ;
      VIA 123.57 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 642.525 124.36 642.855 ;
      VIA 123.57 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 642.505 124.34 642.875 ;
      VIA 123.57 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 635.865 124.36 636.195 ;
      VIA 123.57 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 635.845 124.34 636.215 ;
      VIA 123.57 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 629.205 124.36 629.535 ;
      VIA 123.57 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 629.185 124.34 629.555 ;
      VIA 123.57 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 622.545 124.36 622.875 ;
      VIA 123.57 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 622.525 124.34 622.895 ;
      VIA 123.57 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 615.885 124.36 616.215 ;
      VIA 123.57 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 615.865 124.34 616.235 ;
      VIA 123.57 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 609.225 124.36 609.555 ;
      VIA 123.57 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 609.205 124.34 609.575 ;
      VIA 123.57 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 602.565 124.36 602.895 ;
      VIA 123.57 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 602.545 124.34 602.915 ;
      VIA 123.57 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 595.905 124.36 596.235 ;
      VIA 123.57 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 595.885 124.34 596.255 ;
      VIA 123.57 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 589.245 124.36 589.575 ;
      VIA 123.57 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 589.225 124.34 589.595 ;
      VIA 123.57 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 582.585 124.36 582.915 ;
      VIA 123.57 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 582.565 124.34 582.935 ;
      VIA 123.57 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 575.925 124.36 576.255 ;
      VIA 123.57 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 575.905 124.34 576.275 ;
      VIA 123.57 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 569.265 124.36 569.595 ;
      VIA 123.57 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 569.245 124.34 569.615 ;
      VIA 123.57 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 562.605 124.36 562.935 ;
      VIA 123.57 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 562.585 124.34 562.955 ;
      VIA 123.57 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 555.945 124.36 556.275 ;
      VIA 123.57 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 555.925 124.34 556.295 ;
      VIA 123.57 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 549.285 124.36 549.615 ;
      VIA 123.57 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 549.265 124.34 549.635 ;
      VIA 123.57 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 542.625 124.36 542.955 ;
      VIA 123.57 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 542.605 124.34 542.975 ;
      VIA 123.57 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 535.965 124.36 536.295 ;
      VIA 123.57 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 535.945 124.34 536.315 ;
      VIA 123.57 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 529.305 124.36 529.635 ;
      VIA 123.57 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 529.285 124.34 529.655 ;
      VIA 123.57 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 522.645 124.36 522.975 ;
      VIA 123.57 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 522.625 124.34 522.995 ;
      VIA 123.57 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 515.985 124.36 516.315 ;
      VIA 123.57 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 515.965 124.34 516.335 ;
      VIA 123.57 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 509.325 124.36 509.655 ;
      VIA 123.57 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 509.305 124.34 509.675 ;
      VIA 123.57 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 502.665 124.36 502.995 ;
      VIA 123.57 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 502.645 124.34 503.015 ;
      VIA 123.57 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 496.005 124.36 496.335 ;
      VIA 123.57 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 495.985 124.34 496.355 ;
      VIA 123.57 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 489.345 124.36 489.675 ;
      VIA 123.57 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 489.325 124.34 489.695 ;
      VIA 123.57 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 482.685 124.36 483.015 ;
      VIA 123.57 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 482.665 124.34 483.035 ;
      VIA 123.57 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 476.025 124.36 476.355 ;
      VIA 123.57 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 476.005 124.34 476.375 ;
      VIA 123.57 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 469.365 124.36 469.695 ;
      VIA 123.57 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 469.345 124.34 469.715 ;
      VIA 123.57 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 462.705 124.36 463.035 ;
      VIA 123.57 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 462.685 124.34 463.055 ;
      VIA 123.57 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 456.045 124.36 456.375 ;
      VIA 123.57 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 456.025 124.34 456.395 ;
      VIA 123.57 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 449.385 124.36 449.715 ;
      VIA 123.57 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 449.365 124.34 449.735 ;
      VIA 123.57 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 442.725 124.36 443.055 ;
      VIA 123.57 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 442.705 124.34 443.075 ;
      VIA 123.57 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 436.065 124.36 436.395 ;
      VIA 123.57 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 436.045 124.34 436.415 ;
      VIA 123.57 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 429.405 124.36 429.735 ;
      VIA 123.57 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 429.385 124.34 429.755 ;
      VIA 123.57 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 422.745 124.36 423.075 ;
      VIA 123.57 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 422.725 124.34 423.095 ;
      VIA 123.57 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 416.085 124.36 416.415 ;
      VIA 123.57 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 416.065 124.34 416.435 ;
      VIA 123.57 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 409.425 124.36 409.755 ;
      VIA 123.57 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 409.405 124.34 409.775 ;
      VIA 123.57 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 402.765 124.36 403.095 ;
      VIA 123.57 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 402.745 124.34 403.115 ;
      VIA 123.57 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 396.105 124.36 396.435 ;
      VIA 123.57 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 396.085 124.34 396.455 ;
      VIA 123.57 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 389.445 124.36 389.775 ;
      VIA 123.57 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 389.425 124.34 389.795 ;
      VIA 123.57 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 382.785 124.36 383.115 ;
      VIA 123.57 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 382.765 124.34 383.135 ;
      VIA 123.57 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 376.125 124.36 376.455 ;
      VIA 123.57 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 376.105 124.34 376.475 ;
      VIA 123.57 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 369.465 124.36 369.795 ;
      VIA 123.57 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 369.445 124.34 369.815 ;
      VIA 123.57 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 362.805 124.36 363.135 ;
      VIA 123.57 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 362.785 124.34 363.155 ;
      VIA 123.57 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 356.145 124.36 356.475 ;
      VIA 123.57 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 356.125 124.34 356.495 ;
      VIA 123.57 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 349.485 124.36 349.815 ;
      VIA 123.57 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 349.465 124.34 349.835 ;
      VIA 123.57 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 342.825 124.36 343.155 ;
      VIA 123.57 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 342.805 124.34 343.175 ;
      VIA 123.57 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 336.165 124.36 336.495 ;
      VIA 123.57 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 336.145 124.34 336.515 ;
      VIA 123.57 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 329.505 124.36 329.835 ;
      VIA 123.57 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 329.485 124.34 329.855 ;
      VIA 123.57 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 322.845 124.36 323.175 ;
      VIA 123.57 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 322.825 124.34 323.195 ;
      VIA 123.57 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 316.185 124.36 316.515 ;
      VIA 123.57 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 316.165 124.34 316.535 ;
      VIA 123.57 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 309.525 124.36 309.855 ;
      VIA 123.57 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 309.505 124.34 309.875 ;
      VIA 123.57 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 302.865 124.36 303.195 ;
      VIA 123.57 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 302.845 124.34 303.215 ;
      VIA 123.57 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 296.205 124.36 296.535 ;
      VIA 123.57 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 296.185 124.34 296.555 ;
      VIA 123.57 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 289.545 124.36 289.875 ;
      VIA 123.57 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 289.525 124.34 289.895 ;
      VIA 123.57 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 282.885 124.36 283.215 ;
      VIA 123.57 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 282.865 124.34 283.235 ;
      VIA 123.57 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 276.225 124.36 276.555 ;
      VIA 123.57 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 276.205 124.34 276.575 ;
      VIA 123.57 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 269.565 124.36 269.895 ;
      VIA 123.57 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 269.545 124.34 269.915 ;
      VIA 123.57 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 262.905 124.36 263.235 ;
      VIA 123.57 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 262.885 124.34 263.255 ;
      VIA 123.57 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 256.245 124.36 256.575 ;
      VIA 123.57 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 256.225 124.34 256.595 ;
      VIA 123.57 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 249.585 124.36 249.915 ;
      VIA 123.57 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 249.565 124.34 249.935 ;
      VIA 123.57 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 242.925 124.36 243.255 ;
      VIA 123.57 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 242.905 124.34 243.275 ;
      VIA 123.57 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 236.265 124.36 236.595 ;
      VIA 123.57 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 236.245 124.34 236.615 ;
      VIA 123.57 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 229.605 124.36 229.935 ;
      VIA 123.57 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 229.585 124.34 229.955 ;
      VIA 123.57 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 222.945 124.36 223.275 ;
      VIA 123.57 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 222.925 124.34 223.295 ;
      VIA 123.57 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 216.285 124.36 216.615 ;
      VIA 123.57 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 216.265 124.34 216.635 ;
      VIA 123.57 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 209.625 124.36 209.955 ;
      VIA 123.57 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 209.605 124.34 209.975 ;
      VIA 123.57 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 202.965 124.36 203.295 ;
      VIA 123.57 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 202.945 124.34 203.315 ;
      VIA 123.57 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 196.305 124.36 196.635 ;
      VIA 123.57 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 196.285 124.34 196.655 ;
      VIA 123.57 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 189.645 124.36 189.975 ;
      VIA 123.57 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 189.625 124.34 189.995 ;
      VIA 123.57 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 182.985 124.36 183.315 ;
      VIA 123.57 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 182.965 124.34 183.335 ;
      VIA 123.57 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 176.325 124.36 176.655 ;
      VIA 123.57 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 176.305 124.34 176.675 ;
      VIA 123.57 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 169.665 124.36 169.995 ;
      VIA 123.57 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 169.645 124.34 170.015 ;
      VIA 123.57 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 163.005 124.36 163.335 ;
      VIA 123.57 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 162.985 124.34 163.355 ;
      VIA 123.57 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 156.345 124.36 156.675 ;
      VIA 123.57 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 156.325 124.34 156.695 ;
      VIA 123.57 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 149.685 124.36 150.015 ;
      VIA 123.57 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 149.665 124.34 150.035 ;
      VIA 123.57 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 143.025 124.36 143.355 ;
      VIA 123.57 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 143.005 124.34 143.375 ;
      VIA 123.57 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 136.365 124.36 136.695 ;
      VIA 123.57 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 136.345 124.34 136.715 ;
      VIA 123.57 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 129.705 124.36 130.035 ;
      VIA 123.57 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 129.685 124.34 130.055 ;
      VIA 123.57 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 123.045 124.36 123.375 ;
      VIA 123.57 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 123.025 124.34 123.395 ;
      VIA 123.57 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 116.385 124.36 116.715 ;
      VIA 123.57 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 116.365 124.34 116.735 ;
      VIA 123.57 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 109.725 124.36 110.055 ;
      VIA 123.57 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 109.705 124.34 110.075 ;
      VIA 123.57 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 103.065 124.36 103.395 ;
      VIA 123.57 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 103.045 124.34 103.415 ;
      VIA 123.57 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 96.405 124.36 96.735 ;
      VIA 123.57 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 96.385 124.34 96.755 ;
      VIA 123.57 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 89.745 124.36 90.075 ;
      VIA 123.57 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 89.725 124.34 90.095 ;
      VIA 123.57 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 83.085 124.36 83.415 ;
      VIA 123.57 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 83.065 124.34 83.435 ;
      VIA 123.57 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 76.425 124.36 76.755 ;
      VIA 123.57 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 76.405 124.34 76.775 ;
      VIA 123.57 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 69.765 124.36 70.095 ;
      VIA 123.57 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 69.745 124.34 70.115 ;
      VIA 123.57 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 63.105 124.36 63.435 ;
      VIA 123.57 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 63.085 124.34 63.455 ;
      VIA 123.57 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 56.445 124.36 56.775 ;
      VIA 123.57 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 56.425 124.34 56.795 ;
      VIA 123.57 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 49.785 124.36 50.115 ;
      VIA 123.57 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 49.765 124.34 50.135 ;
      VIA 123.57 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 43.125 124.36 43.455 ;
      VIA 123.57 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 43.105 124.34 43.475 ;
      VIA 123.57 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 36.465 124.36 36.795 ;
      VIA 123.57 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 36.445 124.34 36.815 ;
      VIA 123.57 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 29.805 124.36 30.135 ;
      VIA 123.57 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 29.785 124.34 30.155 ;
      VIA 123.57 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 23.145 124.36 23.475 ;
      VIA 123.57 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 23.125 124.34 23.495 ;
      VIA 123.57 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 16.485 124.36 16.815 ;
      VIA 123.57 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 16.465 124.34 16.835 ;
      VIA 123.57 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 9.825 124.36 10.155 ;
      VIA 123.57 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 9.805 124.34 10.175 ;
      VIA 123.57 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.78 3.165 124.36 3.495 ;
      VIA 123.57 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.8 3.145 124.34 3.515 ;
      VIA 123.57 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 123.57 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 775.725 97.22 776.055 ;
      VIA 96.43 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 775.705 97.2 776.075 ;
      VIA 96.43 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 769.065 97.22 769.395 ;
      VIA 96.43 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 769.045 97.2 769.415 ;
      VIA 96.43 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 762.405 97.22 762.735 ;
      VIA 96.43 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 762.385 97.2 762.755 ;
      VIA 96.43 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 755.745 97.22 756.075 ;
      VIA 96.43 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 755.725 97.2 756.095 ;
      VIA 96.43 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 749.085 97.22 749.415 ;
      VIA 96.43 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 749.065 97.2 749.435 ;
      VIA 96.43 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 742.425 97.22 742.755 ;
      VIA 96.43 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 742.405 97.2 742.775 ;
      VIA 96.43 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 735.765 97.22 736.095 ;
      VIA 96.43 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 735.745 97.2 736.115 ;
      VIA 96.43 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 729.105 97.22 729.435 ;
      VIA 96.43 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 729.085 97.2 729.455 ;
      VIA 96.43 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 722.445 97.22 722.775 ;
      VIA 96.43 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 722.425 97.2 722.795 ;
      VIA 96.43 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 715.785 97.22 716.115 ;
      VIA 96.43 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 715.765 97.2 716.135 ;
      VIA 96.43 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 709.125 97.22 709.455 ;
      VIA 96.43 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 709.105 97.2 709.475 ;
      VIA 96.43 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 702.465 97.22 702.795 ;
      VIA 96.43 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 702.445 97.2 702.815 ;
      VIA 96.43 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 695.805 97.22 696.135 ;
      VIA 96.43 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 695.785 97.2 696.155 ;
      VIA 96.43 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 689.145 97.22 689.475 ;
      VIA 96.43 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 689.125 97.2 689.495 ;
      VIA 96.43 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 682.485 97.22 682.815 ;
      VIA 96.43 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 682.465 97.2 682.835 ;
      VIA 96.43 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 675.825 97.22 676.155 ;
      VIA 96.43 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 675.805 97.2 676.175 ;
      VIA 96.43 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 669.165 97.22 669.495 ;
      VIA 96.43 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 669.145 97.2 669.515 ;
      VIA 96.43 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 662.505 97.22 662.835 ;
      VIA 96.43 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 662.485 97.2 662.855 ;
      VIA 96.43 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 655.845 97.22 656.175 ;
      VIA 96.43 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 655.825 97.2 656.195 ;
      VIA 96.43 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 649.185 97.22 649.515 ;
      VIA 96.43 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 649.165 97.2 649.535 ;
      VIA 96.43 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 642.525 97.22 642.855 ;
      VIA 96.43 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 642.505 97.2 642.875 ;
      VIA 96.43 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 635.865 97.22 636.195 ;
      VIA 96.43 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 635.845 97.2 636.215 ;
      VIA 96.43 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 629.205 97.22 629.535 ;
      VIA 96.43 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 629.185 97.2 629.555 ;
      VIA 96.43 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 622.545 97.22 622.875 ;
      VIA 96.43 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 622.525 97.2 622.895 ;
      VIA 96.43 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 615.885 97.22 616.215 ;
      VIA 96.43 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 615.865 97.2 616.235 ;
      VIA 96.43 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 609.225 97.22 609.555 ;
      VIA 96.43 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 609.205 97.2 609.575 ;
      VIA 96.43 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 602.565 97.22 602.895 ;
      VIA 96.43 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 602.545 97.2 602.915 ;
      VIA 96.43 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 595.905 97.22 596.235 ;
      VIA 96.43 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 595.885 97.2 596.255 ;
      VIA 96.43 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 589.245 97.22 589.575 ;
      VIA 96.43 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 589.225 97.2 589.595 ;
      VIA 96.43 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 582.585 97.22 582.915 ;
      VIA 96.43 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 582.565 97.2 582.935 ;
      VIA 96.43 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 575.925 97.22 576.255 ;
      VIA 96.43 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 575.905 97.2 576.275 ;
      VIA 96.43 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 569.265 97.22 569.595 ;
      VIA 96.43 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 569.245 97.2 569.615 ;
      VIA 96.43 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 562.605 97.22 562.935 ;
      VIA 96.43 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 562.585 97.2 562.955 ;
      VIA 96.43 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 555.945 97.22 556.275 ;
      VIA 96.43 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 555.925 97.2 556.295 ;
      VIA 96.43 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 549.285 97.22 549.615 ;
      VIA 96.43 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 549.265 97.2 549.635 ;
      VIA 96.43 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 542.625 97.22 542.955 ;
      VIA 96.43 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 542.605 97.2 542.975 ;
      VIA 96.43 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 535.965 97.22 536.295 ;
      VIA 96.43 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 535.945 97.2 536.315 ;
      VIA 96.43 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 529.305 97.22 529.635 ;
      VIA 96.43 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 529.285 97.2 529.655 ;
      VIA 96.43 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 522.645 97.22 522.975 ;
      VIA 96.43 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 522.625 97.2 522.995 ;
      VIA 96.43 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 515.985 97.22 516.315 ;
      VIA 96.43 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 515.965 97.2 516.335 ;
      VIA 96.43 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 509.325 97.22 509.655 ;
      VIA 96.43 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 509.305 97.2 509.675 ;
      VIA 96.43 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 502.665 97.22 502.995 ;
      VIA 96.43 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 502.645 97.2 503.015 ;
      VIA 96.43 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 496.005 97.22 496.335 ;
      VIA 96.43 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 495.985 97.2 496.355 ;
      VIA 96.43 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 489.345 97.22 489.675 ;
      VIA 96.43 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 489.325 97.2 489.695 ;
      VIA 96.43 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 482.685 97.22 483.015 ;
      VIA 96.43 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 482.665 97.2 483.035 ;
      VIA 96.43 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 476.025 97.22 476.355 ;
      VIA 96.43 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 476.005 97.2 476.375 ;
      VIA 96.43 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 469.365 97.22 469.695 ;
      VIA 96.43 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 469.345 97.2 469.715 ;
      VIA 96.43 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 462.705 97.22 463.035 ;
      VIA 96.43 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 462.685 97.2 463.055 ;
      VIA 96.43 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 456.045 97.22 456.375 ;
      VIA 96.43 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 456.025 97.2 456.395 ;
      VIA 96.43 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 449.385 97.22 449.715 ;
      VIA 96.43 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 449.365 97.2 449.735 ;
      VIA 96.43 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 442.725 97.22 443.055 ;
      VIA 96.43 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 442.705 97.2 443.075 ;
      VIA 96.43 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 436.065 97.22 436.395 ;
      VIA 96.43 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 436.045 97.2 436.415 ;
      VIA 96.43 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 429.405 97.22 429.735 ;
      VIA 96.43 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 429.385 97.2 429.755 ;
      VIA 96.43 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 422.745 97.22 423.075 ;
      VIA 96.43 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 422.725 97.2 423.095 ;
      VIA 96.43 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 416.085 97.22 416.415 ;
      VIA 96.43 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 416.065 97.2 416.435 ;
      VIA 96.43 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 409.425 97.22 409.755 ;
      VIA 96.43 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 409.405 97.2 409.775 ;
      VIA 96.43 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 402.765 97.22 403.095 ;
      VIA 96.43 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 402.745 97.2 403.115 ;
      VIA 96.43 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 396.105 97.22 396.435 ;
      VIA 96.43 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 396.085 97.2 396.455 ;
      VIA 96.43 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 389.445 97.22 389.775 ;
      VIA 96.43 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 389.425 97.2 389.795 ;
      VIA 96.43 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 382.785 97.22 383.115 ;
      VIA 96.43 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 382.765 97.2 383.135 ;
      VIA 96.43 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 376.125 97.22 376.455 ;
      VIA 96.43 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 376.105 97.2 376.475 ;
      VIA 96.43 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 369.465 97.22 369.795 ;
      VIA 96.43 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 369.445 97.2 369.815 ;
      VIA 96.43 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 362.805 97.22 363.135 ;
      VIA 96.43 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 362.785 97.2 363.155 ;
      VIA 96.43 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 356.145 97.22 356.475 ;
      VIA 96.43 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 356.125 97.2 356.495 ;
      VIA 96.43 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 349.485 97.22 349.815 ;
      VIA 96.43 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 349.465 97.2 349.835 ;
      VIA 96.43 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 342.825 97.22 343.155 ;
      VIA 96.43 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 342.805 97.2 343.175 ;
      VIA 96.43 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 336.165 97.22 336.495 ;
      VIA 96.43 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 336.145 97.2 336.515 ;
      VIA 96.43 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 329.505 97.22 329.835 ;
      VIA 96.43 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 329.485 97.2 329.855 ;
      VIA 96.43 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 322.845 97.22 323.175 ;
      VIA 96.43 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 322.825 97.2 323.195 ;
      VIA 96.43 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 316.185 97.22 316.515 ;
      VIA 96.43 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 316.165 97.2 316.535 ;
      VIA 96.43 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 309.525 97.22 309.855 ;
      VIA 96.43 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 309.505 97.2 309.875 ;
      VIA 96.43 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 302.865 97.22 303.195 ;
      VIA 96.43 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 302.845 97.2 303.215 ;
      VIA 96.43 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 296.205 97.22 296.535 ;
      VIA 96.43 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 296.185 97.2 296.555 ;
      VIA 96.43 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 289.545 97.22 289.875 ;
      VIA 96.43 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 289.525 97.2 289.895 ;
      VIA 96.43 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 282.885 97.22 283.215 ;
      VIA 96.43 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 282.865 97.2 283.235 ;
      VIA 96.43 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 276.225 97.22 276.555 ;
      VIA 96.43 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 276.205 97.2 276.575 ;
      VIA 96.43 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 269.565 97.22 269.895 ;
      VIA 96.43 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 269.545 97.2 269.915 ;
      VIA 96.43 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 262.905 97.22 263.235 ;
      VIA 96.43 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 262.885 97.2 263.255 ;
      VIA 96.43 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 256.245 97.22 256.575 ;
      VIA 96.43 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 256.225 97.2 256.595 ;
      VIA 96.43 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 249.585 97.22 249.915 ;
      VIA 96.43 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 249.565 97.2 249.935 ;
      VIA 96.43 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 242.925 97.22 243.255 ;
      VIA 96.43 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 242.905 97.2 243.275 ;
      VIA 96.43 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 236.265 97.22 236.595 ;
      VIA 96.43 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 236.245 97.2 236.615 ;
      VIA 96.43 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 229.605 97.22 229.935 ;
      VIA 96.43 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 229.585 97.2 229.955 ;
      VIA 96.43 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 222.945 97.22 223.275 ;
      VIA 96.43 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 222.925 97.2 223.295 ;
      VIA 96.43 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 216.285 97.22 216.615 ;
      VIA 96.43 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 216.265 97.2 216.635 ;
      VIA 96.43 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 209.625 97.22 209.955 ;
      VIA 96.43 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 209.605 97.2 209.975 ;
      VIA 96.43 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 202.965 97.22 203.295 ;
      VIA 96.43 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 202.945 97.2 203.315 ;
      VIA 96.43 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 196.305 97.22 196.635 ;
      VIA 96.43 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 196.285 97.2 196.655 ;
      VIA 96.43 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 189.645 97.22 189.975 ;
      VIA 96.43 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 189.625 97.2 189.995 ;
      VIA 96.43 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 182.985 97.22 183.315 ;
      VIA 96.43 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 182.965 97.2 183.335 ;
      VIA 96.43 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 176.325 97.22 176.655 ;
      VIA 96.43 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 176.305 97.2 176.675 ;
      VIA 96.43 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 169.665 97.22 169.995 ;
      VIA 96.43 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 169.645 97.2 170.015 ;
      VIA 96.43 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 163.005 97.22 163.335 ;
      VIA 96.43 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 162.985 97.2 163.355 ;
      VIA 96.43 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 156.345 97.22 156.675 ;
      VIA 96.43 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 156.325 97.2 156.695 ;
      VIA 96.43 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 149.685 97.22 150.015 ;
      VIA 96.43 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 149.665 97.2 150.035 ;
      VIA 96.43 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 143.025 97.22 143.355 ;
      VIA 96.43 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 143.005 97.2 143.375 ;
      VIA 96.43 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 136.365 97.22 136.695 ;
      VIA 96.43 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 136.345 97.2 136.715 ;
      VIA 96.43 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 129.705 97.22 130.035 ;
      VIA 96.43 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 129.685 97.2 130.055 ;
      VIA 96.43 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 123.045 97.22 123.375 ;
      VIA 96.43 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 123.025 97.2 123.395 ;
      VIA 96.43 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 116.385 97.22 116.715 ;
      VIA 96.43 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 116.365 97.2 116.735 ;
      VIA 96.43 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 109.725 97.22 110.055 ;
      VIA 96.43 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 109.705 97.2 110.075 ;
      VIA 96.43 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 103.065 97.22 103.395 ;
      VIA 96.43 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 103.045 97.2 103.415 ;
      VIA 96.43 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 96.405 97.22 96.735 ;
      VIA 96.43 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 96.385 97.2 96.755 ;
      VIA 96.43 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 89.745 97.22 90.075 ;
      VIA 96.43 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 89.725 97.2 90.095 ;
      VIA 96.43 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 83.085 97.22 83.415 ;
      VIA 96.43 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 83.065 97.2 83.435 ;
      VIA 96.43 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 76.425 97.22 76.755 ;
      VIA 96.43 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 76.405 97.2 76.775 ;
      VIA 96.43 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 69.765 97.22 70.095 ;
      VIA 96.43 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 69.745 97.2 70.115 ;
      VIA 96.43 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 63.105 97.22 63.435 ;
      VIA 96.43 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 63.085 97.2 63.455 ;
      VIA 96.43 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 56.445 97.22 56.775 ;
      VIA 96.43 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 56.425 97.2 56.795 ;
      VIA 96.43 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 49.785 97.22 50.115 ;
      VIA 96.43 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 49.765 97.2 50.135 ;
      VIA 96.43 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 43.125 97.22 43.455 ;
      VIA 96.43 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 43.105 97.2 43.475 ;
      VIA 96.43 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 36.465 97.22 36.795 ;
      VIA 96.43 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 36.445 97.2 36.815 ;
      VIA 96.43 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 29.805 97.22 30.135 ;
      VIA 96.43 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 29.785 97.2 30.155 ;
      VIA 96.43 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 23.145 97.22 23.475 ;
      VIA 96.43 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 23.125 97.2 23.495 ;
      VIA 96.43 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 16.485 97.22 16.815 ;
      VIA 96.43 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 16.465 97.2 16.835 ;
      VIA 96.43 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 9.825 97.22 10.155 ;
      VIA 96.43 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 9.805 97.2 10.175 ;
      VIA 96.43 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.64 3.165 97.22 3.495 ;
      VIA 96.43 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.66 3.145 97.2 3.515 ;
      VIA 96.43 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 96.43 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 775.725 70.08 776.055 ;
      VIA 69.29 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 775.705 70.06 776.075 ;
      VIA 69.29 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 769.065 70.08 769.395 ;
      VIA 69.29 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 769.045 70.06 769.415 ;
      VIA 69.29 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 762.405 70.08 762.735 ;
      VIA 69.29 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 762.385 70.06 762.755 ;
      VIA 69.29 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 755.745 70.08 756.075 ;
      VIA 69.29 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 755.725 70.06 756.095 ;
      VIA 69.29 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 749.085 70.08 749.415 ;
      VIA 69.29 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 749.065 70.06 749.435 ;
      VIA 69.29 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 742.425 70.08 742.755 ;
      VIA 69.29 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 742.405 70.06 742.775 ;
      VIA 69.29 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 735.765 70.08 736.095 ;
      VIA 69.29 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 735.745 70.06 736.115 ;
      VIA 69.29 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 729.105 70.08 729.435 ;
      VIA 69.29 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 729.085 70.06 729.455 ;
      VIA 69.29 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 722.445 70.08 722.775 ;
      VIA 69.29 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 722.425 70.06 722.795 ;
      VIA 69.29 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 715.785 70.08 716.115 ;
      VIA 69.29 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 715.765 70.06 716.135 ;
      VIA 69.29 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 709.125 70.08 709.455 ;
      VIA 69.29 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 709.105 70.06 709.475 ;
      VIA 69.29 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 702.465 70.08 702.795 ;
      VIA 69.29 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 702.445 70.06 702.815 ;
      VIA 69.29 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 695.805 70.08 696.135 ;
      VIA 69.29 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 695.785 70.06 696.155 ;
      VIA 69.29 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 689.145 70.08 689.475 ;
      VIA 69.29 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 689.125 70.06 689.495 ;
      VIA 69.29 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 682.485 70.08 682.815 ;
      VIA 69.29 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 682.465 70.06 682.835 ;
      VIA 69.29 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 675.825 70.08 676.155 ;
      VIA 69.29 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 675.805 70.06 676.175 ;
      VIA 69.29 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 669.165 70.08 669.495 ;
      VIA 69.29 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 669.145 70.06 669.515 ;
      VIA 69.29 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 662.505 70.08 662.835 ;
      VIA 69.29 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 662.485 70.06 662.855 ;
      VIA 69.29 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 655.845 70.08 656.175 ;
      VIA 69.29 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 655.825 70.06 656.195 ;
      VIA 69.29 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 649.185 70.08 649.515 ;
      VIA 69.29 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 649.165 70.06 649.535 ;
      VIA 69.29 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 642.525 70.08 642.855 ;
      VIA 69.29 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 642.505 70.06 642.875 ;
      VIA 69.29 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 635.865 70.08 636.195 ;
      VIA 69.29 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 635.845 70.06 636.215 ;
      VIA 69.29 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 629.205 70.08 629.535 ;
      VIA 69.29 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 629.185 70.06 629.555 ;
      VIA 69.29 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 622.545 70.08 622.875 ;
      VIA 69.29 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 622.525 70.06 622.895 ;
      VIA 69.29 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 615.885 70.08 616.215 ;
      VIA 69.29 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 615.865 70.06 616.235 ;
      VIA 69.29 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 609.225 70.08 609.555 ;
      VIA 69.29 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 609.205 70.06 609.575 ;
      VIA 69.29 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 602.565 70.08 602.895 ;
      VIA 69.29 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 602.545 70.06 602.915 ;
      VIA 69.29 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 595.905 70.08 596.235 ;
      VIA 69.29 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 595.885 70.06 596.255 ;
      VIA 69.29 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 589.245 70.08 589.575 ;
      VIA 69.29 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 589.225 70.06 589.595 ;
      VIA 69.29 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 582.585 70.08 582.915 ;
      VIA 69.29 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 582.565 70.06 582.935 ;
      VIA 69.29 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 575.925 70.08 576.255 ;
      VIA 69.29 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 575.905 70.06 576.275 ;
      VIA 69.29 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 569.265 70.08 569.595 ;
      VIA 69.29 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 569.245 70.06 569.615 ;
      VIA 69.29 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 562.605 70.08 562.935 ;
      VIA 69.29 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 562.585 70.06 562.955 ;
      VIA 69.29 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 555.945 70.08 556.275 ;
      VIA 69.29 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 555.925 70.06 556.295 ;
      VIA 69.29 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 549.285 70.08 549.615 ;
      VIA 69.29 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 549.265 70.06 549.635 ;
      VIA 69.29 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 542.625 70.08 542.955 ;
      VIA 69.29 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 542.605 70.06 542.975 ;
      VIA 69.29 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 535.965 70.08 536.295 ;
      VIA 69.29 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 535.945 70.06 536.315 ;
      VIA 69.29 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 529.305 70.08 529.635 ;
      VIA 69.29 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 529.285 70.06 529.655 ;
      VIA 69.29 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 522.645 70.08 522.975 ;
      VIA 69.29 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 522.625 70.06 522.995 ;
      VIA 69.29 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 515.985 70.08 516.315 ;
      VIA 69.29 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 515.965 70.06 516.335 ;
      VIA 69.29 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 509.325 70.08 509.655 ;
      VIA 69.29 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 509.305 70.06 509.675 ;
      VIA 69.29 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 502.665 70.08 502.995 ;
      VIA 69.29 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 502.645 70.06 503.015 ;
      VIA 69.29 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 496.005 70.08 496.335 ;
      VIA 69.29 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 495.985 70.06 496.355 ;
      VIA 69.29 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 489.345 70.08 489.675 ;
      VIA 69.29 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 489.325 70.06 489.695 ;
      VIA 69.29 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 482.685 70.08 483.015 ;
      VIA 69.29 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 482.665 70.06 483.035 ;
      VIA 69.29 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 476.025 70.08 476.355 ;
      VIA 69.29 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 476.005 70.06 476.375 ;
      VIA 69.29 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 469.365 70.08 469.695 ;
      VIA 69.29 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 469.345 70.06 469.715 ;
      VIA 69.29 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 462.705 70.08 463.035 ;
      VIA 69.29 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 462.685 70.06 463.055 ;
      VIA 69.29 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 456.045 70.08 456.375 ;
      VIA 69.29 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 456.025 70.06 456.395 ;
      VIA 69.29 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 449.385 70.08 449.715 ;
      VIA 69.29 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 449.365 70.06 449.735 ;
      VIA 69.29 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 442.725 70.08 443.055 ;
      VIA 69.29 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 442.705 70.06 443.075 ;
      VIA 69.29 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 436.065 70.08 436.395 ;
      VIA 69.29 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 436.045 70.06 436.415 ;
      VIA 69.29 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 429.405 70.08 429.735 ;
      VIA 69.29 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 429.385 70.06 429.755 ;
      VIA 69.29 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 422.745 70.08 423.075 ;
      VIA 69.29 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 422.725 70.06 423.095 ;
      VIA 69.29 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 416.085 70.08 416.415 ;
      VIA 69.29 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 416.065 70.06 416.435 ;
      VIA 69.29 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 409.425 70.08 409.755 ;
      VIA 69.29 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 409.405 70.06 409.775 ;
      VIA 69.29 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 402.765 70.08 403.095 ;
      VIA 69.29 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 402.745 70.06 403.115 ;
      VIA 69.29 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 396.105 70.08 396.435 ;
      VIA 69.29 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 396.085 70.06 396.455 ;
      VIA 69.29 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 389.445 70.08 389.775 ;
      VIA 69.29 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 389.425 70.06 389.795 ;
      VIA 69.29 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 382.785 70.08 383.115 ;
      VIA 69.29 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 382.765 70.06 383.135 ;
      VIA 69.29 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 376.125 70.08 376.455 ;
      VIA 69.29 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 376.105 70.06 376.475 ;
      VIA 69.29 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 369.465 70.08 369.795 ;
      VIA 69.29 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 369.445 70.06 369.815 ;
      VIA 69.29 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 362.805 70.08 363.135 ;
      VIA 69.29 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 362.785 70.06 363.155 ;
      VIA 69.29 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 356.145 70.08 356.475 ;
      VIA 69.29 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 356.125 70.06 356.495 ;
      VIA 69.29 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 349.485 70.08 349.815 ;
      VIA 69.29 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 349.465 70.06 349.835 ;
      VIA 69.29 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 342.825 70.08 343.155 ;
      VIA 69.29 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 342.805 70.06 343.175 ;
      VIA 69.29 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 336.165 70.08 336.495 ;
      VIA 69.29 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 336.145 70.06 336.515 ;
      VIA 69.29 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 329.505 70.08 329.835 ;
      VIA 69.29 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 329.485 70.06 329.855 ;
      VIA 69.29 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 322.845 70.08 323.175 ;
      VIA 69.29 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 322.825 70.06 323.195 ;
      VIA 69.29 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 316.185 70.08 316.515 ;
      VIA 69.29 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 316.165 70.06 316.535 ;
      VIA 69.29 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 309.525 70.08 309.855 ;
      VIA 69.29 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 309.505 70.06 309.875 ;
      VIA 69.29 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 302.865 70.08 303.195 ;
      VIA 69.29 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 302.845 70.06 303.215 ;
      VIA 69.29 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 296.205 70.08 296.535 ;
      VIA 69.29 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 296.185 70.06 296.555 ;
      VIA 69.29 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 289.545 70.08 289.875 ;
      VIA 69.29 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 289.525 70.06 289.895 ;
      VIA 69.29 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 282.885 70.08 283.215 ;
      VIA 69.29 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 282.865 70.06 283.235 ;
      VIA 69.29 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 276.225 70.08 276.555 ;
      VIA 69.29 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 276.205 70.06 276.575 ;
      VIA 69.29 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 269.565 70.08 269.895 ;
      VIA 69.29 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 269.545 70.06 269.915 ;
      VIA 69.29 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 262.905 70.08 263.235 ;
      VIA 69.29 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 262.885 70.06 263.255 ;
      VIA 69.29 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 256.245 70.08 256.575 ;
      VIA 69.29 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 256.225 70.06 256.595 ;
      VIA 69.29 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 249.585 70.08 249.915 ;
      VIA 69.29 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 249.565 70.06 249.935 ;
      VIA 69.29 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 242.925 70.08 243.255 ;
      VIA 69.29 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 242.905 70.06 243.275 ;
      VIA 69.29 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 236.265 70.08 236.595 ;
      VIA 69.29 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 236.245 70.06 236.615 ;
      VIA 69.29 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 229.605 70.08 229.935 ;
      VIA 69.29 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 229.585 70.06 229.955 ;
      VIA 69.29 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 222.945 70.08 223.275 ;
      VIA 69.29 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 222.925 70.06 223.295 ;
      VIA 69.29 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 216.285 70.08 216.615 ;
      VIA 69.29 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 216.265 70.06 216.635 ;
      VIA 69.29 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 209.625 70.08 209.955 ;
      VIA 69.29 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 209.605 70.06 209.975 ;
      VIA 69.29 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 202.965 70.08 203.295 ;
      VIA 69.29 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 202.945 70.06 203.315 ;
      VIA 69.29 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 196.305 70.08 196.635 ;
      VIA 69.29 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 196.285 70.06 196.655 ;
      VIA 69.29 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 189.645 70.08 189.975 ;
      VIA 69.29 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 189.625 70.06 189.995 ;
      VIA 69.29 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 182.985 70.08 183.315 ;
      VIA 69.29 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 182.965 70.06 183.335 ;
      VIA 69.29 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 176.325 70.08 176.655 ;
      VIA 69.29 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 176.305 70.06 176.675 ;
      VIA 69.29 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 169.665 70.08 169.995 ;
      VIA 69.29 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 169.645 70.06 170.015 ;
      VIA 69.29 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 163.005 70.08 163.335 ;
      VIA 69.29 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 162.985 70.06 163.355 ;
      VIA 69.29 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 156.345 70.08 156.675 ;
      VIA 69.29 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 156.325 70.06 156.695 ;
      VIA 69.29 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 149.685 70.08 150.015 ;
      VIA 69.29 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 149.665 70.06 150.035 ;
      VIA 69.29 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 143.025 70.08 143.355 ;
      VIA 69.29 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 143.005 70.06 143.375 ;
      VIA 69.29 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 136.365 70.08 136.695 ;
      VIA 69.29 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 136.345 70.06 136.715 ;
      VIA 69.29 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 129.705 70.08 130.035 ;
      VIA 69.29 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 129.685 70.06 130.055 ;
      VIA 69.29 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 123.045 70.08 123.375 ;
      VIA 69.29 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 123.025 70.06 123.395 ;
      VIA 69.29 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 116.385 70.08 116.715 ;
      VIA 69.29 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 116.365 70.06 116.735 ;
      VIA 69.29 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 109.725 70.08 110.055 ;
      VIA 69.29 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 109.705 70.06 110.075 ;
      VIA 69.29 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 103.065 70.08 103.395 ;
      VIA 69.29 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 103.045 70.06 103.415 ;
      VIA 69.29 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 96.405 70.08 96.735 ;
      VIA 69.29 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 96.385 70.06 96.755 ;
      VIA 69.29 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 89.745 70.08 90.075 ;
      VIA 69.29 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 89.725 70.06 90.095 ;
      VIA 69.29 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 83.085 70.08 83.415 ;
      VIA 69.29 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 83.065 70.06 83.435 ;
      VIA 69.29 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 76.425 70.08 76.755 ;
      VIA 69.29 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 76.405 70.06 76.775 ;
      VIA 69.29 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 69.765 70.08 70.095 ;
      VIA 69.29 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 69.745 70.06 70.115 ;
      VIA 69.29 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 63.105 70.08 63.435 ;
      VIA 69.29 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 63.085 70.06 63.455 ;
      VIA 69.29 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 56.445 70.08 56.775 ;
      VIA 69.29 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 56.425 70.06 56.795 ;
      VIA 69.29 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 49.785 70.08 50.115 ;
      VIA 69.29 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 49.765 70.06 50.135 ;
      VIA 69.29 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 43.125 70.08 43.455 ;
      VIA 69.29 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 43.105 70.06 43.475 ;
      VIA 69.29 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 36.465 70.08 36.795 ;
      VIA 69.29 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 36.445 70.06 36.815 ;
      VIA 69.29 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 29.805 70.08 30.135 ;
      VIA 69.29 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 29.785 70.06 30.155 ;
      VIA 69.29 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 23.145 70.08 23.475 ;
      VIA 69.29 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 23.125 70.06 23.495 ;
      VIA 69.29 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 16.485 70.08 16.815 ;
      VIA 69.29 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 16.465 70.06 16.835 ;
      VIA 69.29 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 9.825 70.08 10.155 ;
      VIA 69.29 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 9.805 70.06 10.175 ;
      VIA 69.29 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.5 3.165 70.08 3.495 ;
      VIA 69.29 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.52 3.145 70.06 3.515 ;
      VIA 69.29 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 69.29 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 775.725 42.94 776.055 ;
      VIA 42.15 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 775.705 42.92 776.075 ;
      VIA 42.15 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 769.065 42.94 769.395 ;
      VIA 42.15 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 769.045 42.92 769.415 ;
      VIA 42.15 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 762.405 42.94 762.735 ;
      VIA 42.15 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 762.385 42.92 762.755 ;
      VIA 42.15 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 755.745 42.94 756.075 ;
      VIA 42.15 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 755.725 42.92 756.095 ;
      VIA 42.15 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 749.085 42.94 749.415 ;
      VIA 42.15 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 749.065 42.92 749.435 ;
      VIA 42.15 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 742.425 42.94 742.755 ;
      VIA 42.15 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 742.405 42.92 742.775 ;
      VIA 42.15 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 735.765 42.94 736.095 ;
      VIA 42.15 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 735.745 42.92 736.115 ;
      VIA 42.15 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 729.105 42.94 729.435 ;
      VIA 42.15 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 729.085 42.92 729.455 ;
      VIA 42.15 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 722.445 42.94 722.775 ;
      VIA 42.15 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 722.425 42.92 722.795 ;
      VIA 42.15 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 715.785 42.94 716.115 ;
      VIA 42.15 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 715.765 42.92 716.135 ;
      VIA 42.15 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 709.125 42.94 709.455 ;
      VIA 42.15 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 709.105 42.92 709.475 ;
      VIA 42.15 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 702.465 42.94 702.795 ;
      VIA 42.15 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 702.445 42.92 702.815 ;
      VIA 42.15 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 695.805 42.94 696.135 ;
      VIA 42.15 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 695.785 42.92 696.155 ;
      VIA 42.15 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 689.145 42.94 689.475 ;
      VIA 42.15 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 689.125 42.92 689.495 ;
      VIA 42.15 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 682.485 42.94 682.815 ;
      VIA 42.15 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 682.465 42.92 682.835 ;
      VIA 42.15 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 675.825 42.94 676.155 ;
      VIA 42.15 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 675.805 42.92 676.175 ;
      VIA 42.15 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 669.165 42.94 669.495 ;
      VIA 42.15 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 669.145 42.92 669.515 ;
      VIA 42.15 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 662.505 42.94 662.835 ;
      VIA 42.15 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 662.485 42.92 662.855 ;
      VIA 42.15 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 655.845 42.94 656.175 ;
      VIA 42.15 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 655.825 42.92 656.195 ;
      VIA 42.15 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 649.185 42.94 649.515 ;
      VIA 42.15 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 649.165 42.92 649.535 ;
      VIA 42.15 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 642.525 42.94 642.855 ;
      VIA 42.15 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 642.505 42.92 642.875 ;
      VIA 42.15 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 635.865 42.94 636.195 ;
      VIA 42.15 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 635.845 42.92 636.215 ;
      VIA 42.15 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 629.205 42.94 629.535 ;
      VIA 42.15 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 629.185 42.92 629.555 ;
      VIA 42.15 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 622.545 42.94 622.875 ;
      VIA 42.15 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 622.525 42.92 622.895 ;
      VIA 42.15 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 615.885 42.94 616.215 ;
      VIA 42.15 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 615.865 42.92 616.235 ;
      VIA 42.15 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 609.225 42.94 609.555 ;
      VIA 42.15 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 609.205 42.92 609.575 ;
      VIA 42.15 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 602.565 42.94 602.895 ;
      VIA 42.15 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 602.545 42.92 602.915 ;
      VIA 42.15 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 595.905 42.94 596.235 ;
      VIA 42.15 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 595.885 42.92 596.255 ;
      VIA 42.15 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 589.245 42.94 589.575 ;
      VIA 42.15 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 589.225 42.92 589.595 ;
      VIA 42.15 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 582.585 42.94 582.915 ;
      VIA 42.15 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 582.565 42.92 582.935 ;
      VIA 42.15 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 575.925 42.94 576.255 ;
      VIA 42.15 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 575.905 42.92 576.275 ;
      VIA 42.15 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 569.265 42.94 569.595 ;
      VIA 42.15 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 569.245 42.92 569.615 ;
      VIA 42.15 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 562.605 42.94 562.935 ;
      VIA 42.15 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 562.585 42.92 562.955 ;
      VIA 42.15 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 555.945 42.94 556.275 ;
      VIA 42.15 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 555.925 42.92 556.295 ;
      VIA 42.15 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 549.285 42.94 549.615 ;
      VIA 42.15 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 549.265 42.92 549.635 ;
      VIA 42.15 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 542.625 42.94 542.955 ;
      VIA 42.15 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 542.605 42.92 542.975 ;
      VIA 42.15 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 535.965 42.94 536.295 ;
      VIA 42.15 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 535.945 42.92 536.315 ;
      VIA 42.15 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 529.305 42.94 529.635 ;
      VIA 42.15 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 529.285 42.92 529.655 ;
      VIA 42.15 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 522.645 42.94 522.975 ;
      VIA 42.15 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 522.625 42.92 522.995 ;
      VIA 42.15 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 515.985 42.94 516.315 ;
      VIA 42.15 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 515.965 42.92 516.335 ;
      VIA 42.15 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 509.325 42.94 509.655 ;
      VIA 42.15 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 509.305 42.92 509.675 ;
      VIA 42.15 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 502.665 42.94 502.995 ;
      VIA 42.15 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 502.645 42.92 503.015 ;
      VIA 42.15 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 496.005 42.94 496.335 ;
      VIA 42.15 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 495.985 42.92 496.355 ;
      VIA 42.15 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 489.345 42.94 489.675 ;
      VIA 42.15 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 489.325 42.92 489.695 ;
      VIA 42.15 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 482.685 42.94 483.015 ;
      VIA 42.15 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 482.665 42.92 483.035 ;
      VIA 42.15 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 476.025 42.94 476.355 ;
      VIA 42.15 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 476.005 42.92 476.375 ;
      VIA 42.15 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 469.365 42.94 469.695 ;
      VIA 42.15 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 469.345 42.92 469.715 ;
      VIA 42.15 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 462.705 42.94 463.035 ;
      VIA 42.15 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 462.685 42.92 463.055 ;
      VIA 42.15 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 456.045 42.94 456.375 ;
      VIA 42.15 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 456.025 42.92 456.395 ;
      VIA 42.15 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 449.385 42.94 449.715 ;
      VIA 42.15 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 449.365 42.92 449.735 ;
      VIA 42.15 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 442.725 42.94 443.055 ;
      VIA 42.15 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 442.705 42.92 443.075 ;
      VIA 42.15 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 436.065 42.94 436.395 ;
      VIA 42.15 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 436.045 42.92 436.415 ;
      VIA 42.15 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 429.405 42.94 429.735 ;
      VIA 42.15 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 429.385 42.92 429.755 ;
      VIA 42.15 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 422.745 42.94 423.075 ;
      VIA 42.15 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 422.725 42.92 423.095 ;
      VIA 42.15 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 416.085 42.94 416.415 ;
      VIA 42.15 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 416.065 42.92 416.435 ;
      VIA 42.15 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 409.425 42.94 409.755 ;
      VIA 42.15 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 409.405 42.92 409.775 ;
      VIA 42.15 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 402.765 42.94 403.095 ;
      VIA 42.15 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 402.745 42.92 403.115 ;
      VIA 42.15 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 396.105 42.94 396.435 ;
      VIA 42.15 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 396.085 42.92 396.455 ;
      VIA 42.15 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 389.445 42.94 389.775 ;
      VIA 42.15 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 389.425 42.92 389.795 ;
      VIA 42.15 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 382.785 42.94 383.115 ;
      VIA 42.15 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 382.765 42.92 383.135 ;
      VIA 42.15 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 376.125 42.94 376.455 ;
      VIA 42.15 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 376.105 42.92 376.475 ;
      VIA 42.15 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 369.465 42.94 369.795 ;
      VIA 42.15 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 369.445 42.92 369.815 ;
      VIA 42.15 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 362.805 42.94 363.135 ;
      VIA 42.15 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 362.785 42.92 363.155 ;
      VIA 42.15 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 356.145 42.94 356.475 ;
      VIA 42.15 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 356.125 42.92 356.495 ;
      VIA 42.15 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 349.485 42.94 349.815 ;
      VIA 42.15 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 349.465 42.92 349.835 ;
      VIA 42.15 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 342.825 42.94 343.155 ;
      VIA 42.15 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 342.805 42.92 343.175 ;
      VIA 42.15 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 336.165 42.94 336.495 ;
      VIA 42.15 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 336.145 42.92 336.515 ;
      VIA 42.15 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 329.505 42.94 329.835 ;
      VIA 42.15 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 329.485 42.92 329.855 ;
      VIA 42.15 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 322.845 42.94 323.175 ;
      VIA 42.15 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 322.825 42.92 323.195 ;
      VIA 42.15 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 316.185 42.94 316.515 ;
      VIA 42.15 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 316.165 42.92 316.535 ;
      VIA 42.15 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 309.525 42.94 309.855 ;
      VIA 42.15 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 309.505 42.92 309.875 ;
      VIA 42.15 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 302.865 42.94 303.195 ;
      VIA 42.15 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 302.845 42.92 303.215 ;
      VIA 42.15 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 296.205 42.94 296.535 ;
      VIA 42.15 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 296.185 42.92 296.555 ;
      VIA 42.15 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 289.545 42.94 289.875 ;
      VIA 42.15 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 289.525 42.92 289.895 ;
      VIA 42.15 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 282.885 42.94 283.215 ;
      VIA 42.15 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 282.865 42.92 283.235 ;
      VIA 42.15 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 276.225 42.94 276.555 ;
      VIA 42.15 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 276.205 42.92 276.575 ;
      VIA 42.15 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 269.565 42.94 269.895 ;
      VIA 42.15 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 269.545 42.92 269.915 ;
      VIA 42.15 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 262.905 42.94 263.235 ;
      VIA 42.15 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 262.885 42.92 263.255 ;
      VIA 42.15 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 256.245 42.94 256.575 ;
      VIA 42.15 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 256.225 42.92 256.595 ;
      VIA 42.15 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 249.585 42.94 249.915 ;
      VIA 42.15 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 249.565 42.92 249.935 ;
      VIA 42.15 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 242.925 42.94 243.255 ;
      VIA 42.15 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 242.905 42.92 243.275 ;
      VIA 42.15 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 236.265 42.94 236.595 ;
      VIA 42.15 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 236.245 42.92 236.615 ;
      VIA 42.15 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 229.605 42.94 229.935 ;
      VIA 42.15 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 229.585 42.92 229.955 ;
      VIA 42.15 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 222.945 42.94 223.275 ;
      VIA 42.15 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 222.925 42.92 223.295 ;
      VIA 42.15 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 216.285 42.94 216.615 ;
      VIA 42.15 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 216.265 42.92 216.635 ;
      VIA 42.15 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 209.625 42.94 209.955 ;
      VIA 42.15 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 209.605 42.92 209.975 ;
      VIA 42.15 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 202.965 42.94 203.295 ;
      VIA 42.15 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 202.945 42.92 203.315 ;
      VIA 42.15 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 196.305 42.94 196.635 ;
      VIA 42.15 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 196.285 42.92 196.655 ;
      VIA 42.15 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 189.645 42.94 189.975 ;
      VIA 42.15 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 189.625 42.92 189.995 ;
      VIA 42.15 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 182.985 42.94 183.315 ;
      VIA 42.15 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 182.965 42.92 183.335 ;
      VIA 42.15 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 176.325 42.94 176.655 ;
      VIA 42.15 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 176.305 42.92 176.675 ;
      VIA 42.15 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 169.665 42.94 169.995 ;
      VIA 42.15 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 169.645 42.92 170.015 ;
      VIA 42.15 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 163.005 42.94 163.335 ;
      VIA 42.15 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 162.985 42.92 163.355 ;
      VIA 42.15 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 156.345 42.94 156.675 ;
      VIA 42.15 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 156.325 42.92 156.695 ;
      VIA 42.15 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 149.685 42.94 150.015 ;
      VIA 42.15 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 149.665 42.92 150.035 ;
      VIA 42.15 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 143.025 42.94 143.355 ;
      VIA 42.15 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 143.005 42.92 143.375 ;
      VIA 42.15 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 136.365 42.94 136.695 ;
      VIA 42.15 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 136.345 42.92 136.715 ;
      VIA 42.15 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 129.705 42.94 130.035 ;
      VIA 42.15 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 129.685 42.92 130.055 ;
      VIA 42.15 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 123.045 42.94 123.375 ;
      VIA 42.15 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 123.025 42.92 123.395 ;
      VIA 42.15 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 116.385 42.94 116.715 ;
      VIA 42.15 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 116.365 42.92 116.735 ;
      VIA 42.15 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 109.725 42.94 110.055 ;
      VIA 42.15 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 109.705 42.92 110.075 ;
      VIA 42.15 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 103.065 42.94 103.395 ;
      VIA 42.15 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 103.045 42.92 103.415 ;
      VIA 42.15 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 96.405 42.94 96.735 ;
      VIA 42.15 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 96.385 42.92 96.755 ;
      VIA 42.15 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 89.745 42.94 90.075 ;
      VIA 42.15 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 89.725 42.92 90.095 ;
      VIA 42.15 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 83.085 42.94 83.415 ;
      VIA 42.15 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 83.065 42.92 83.435 ;
      VIA 42.15 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 76.425 42.94 76.755 ;
      VIA 42.15 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 76.405 42.92 76.775 ;
      VIA 42.15 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 69.765 42.94 70.095 ;
      VIA 42.15 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 69.745 42.92 70.115 ;
      VIA 42.15 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 63.105 42.94 63.435 ;
      VIA 42.15 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 63.085 42.92 63.455 ;
      VIA 42.15 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 56.445 42.94 56.775 ;
      VIA 42.15 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 56.425 42.92 56.795 ;
      VIA 42.15 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 49.785 42.94 50.115 ;
      VIA 42.15 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 49.765 42.92 50.135 ;
      VIA 42.15 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 43.125 42.94 43.455 ;
      VIA 42.15 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 43.105 42.92 43.475 ;
      VIA 42.15 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 36.465 42.94 36.795 ;
      VIA 42.15 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 36.445 42.92 36.815 ;
      VIA 42.15 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 29.805 42.94 30.135 ;
      VIA 42.15 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 29.785 42.92 30.155 ;
      VIA 42.15 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 23.145 42.94 23.475 ;
      VIA 42.15 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 23.125 42.92 23.495 ;
      VIA 42.15 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 16.485 42.94 16.815 ;
      VIA 42.15 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 16.465 42.92 16.835 ;
      VIA 42.15 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 9.825 42.94 10.155 ;
      VIA 42.15 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 9.805 42.92 10.175 ;
      VIA 42.15 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.36 3.165 42.94 3.495 ;
      VIA 42.15 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.38 3.145 42.92 3.515 ;
      VIA 42.15 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 42.15 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 775.725 15.8 776.055 ;
      VIA 15.01 775.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 775.705 15.78 776.075 ;
      VIA 15.01 775.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 775.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 769.065 15.8 769.395 ;
      VIA 15.01 769.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 769.045 15.78 769.415 ;
      VIA 15.01 769.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 769.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 762.405 15.8 762.735 ;
      VIA 15.01 762.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 762.385 15.78 762.755 ;
      VIA 15.01 762.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 762.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 755.745 15.8 756.075 ;
      VIA 15.01 755.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 755.725 15.78 756.095 ;
      VIA 15.01 755.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 755.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 749.085 15.8 749.415 ;
      VIA 15.01 749.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 749.065 15.78 749.435 ;
      VIA 15.01 749.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 749.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 742.425 15.8 742.755 ;
      VIA 15.01 742.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 742.405 15.78 742.775 ;
      VIA 15.01 742.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 742.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 735.765 15.8 736.095 ;
      VIA 15.01 735.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 735.745 15.78 736.115 ;
      VIA 15.01 735.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 735.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 729.105 15.8 729.435 ;
      VIA 15.01 729.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 729.085 15.78 729.455 ;
      VIA 15.01 729.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 729.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 722.445 15.8 722.775 ;
      VIA 15.01 722.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 722.425 15.78 722.795 ;
      VIA 15.01 722.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 722.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 715.785 15.8 716.115 ;
      VIA 15.01 715.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 715.765 15.78 716.135 ;
      VIA 15.01 715.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 715.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 709.125 15.8 709.455 ;
      VIA 15.01 709.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 709.105 15.78 709.475 ;
      VIA 15.01 709.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 709.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 702.465 15.8 702.795 ;
      VIA 15.01 702.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 702.445 15.78 702.815 ;
      VIA 15.01 702.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 702.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 695.805 15.8 696.135 ;
      VIA 15.01 695.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 695.785 15.78 696.155 ;
      VIA 15.01 695.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 695.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 689.145 15.8 689.475 ;
      VIA 15.01 689.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 689.125 15.78 689.495 ;
      VIA 15.01 689.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 689.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 682.485 15.8 682.815 ;
      VIA 15.01 682.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 682.465 15.78 682.835 ;
      VIA 15.01 682.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 682.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 675.825 15.8 676.155 ;
      VIA 15.01 675.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 675.805 15.78 676.175 ;
      VIA 15.01 675.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 675.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 669.165 15.8 669.495 ;
      VIA 15.01 669.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 669.145 15.78 669.515 ;
      VIA 15.01 669.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 669.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 662.505 15.8 662.835 ;
      VIA 15.01 662.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 662.485 15.78 662.855 ;
      VIA 15.01 662.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 662.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 655.845 15.8 656.175 ;
      VIA 15.01 656.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 655.825 15.78 656.195 ;
      VIA 15.01 656.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 656.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 649.185 15.8 649.515 ;
      VIA 15.01 649.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 649.165 15.78 649.535 ;
      VIA 15.01 649.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 649.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 642.525 15.8 642.855 ;
      VIA 15.01 642.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 642.505 15.78 642.875 ;
      VIA 15.01 642.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 642.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 635.865 15.8 636.195 ;
      VIA 15.01 636.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 635.845 15.78 636.215 ;
      VIA 15.01 636.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 636.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 629.205 15.8 629.535 ;
      VIA 15.01 629.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 629.185 15.78 629.555 ;
      VIA 15.01 629.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 629.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 622.545 15.8 622.875 ;
      VIA 15.01 622.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 622.525 15.78 622.895 ;
      VIA 15.01 622.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 622.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 615.885 15.8 616.215 ;
      VIA 15.01 616.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 615.865 15.78 616.235 ;
      VIA 15.01 616.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 616.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 609.225 15.8 609.555 ;
      VIA 15.01 609.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 609.205 15.78 609.575 ;
      VIA 15.01 609.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 609.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 602.565 15.8 602.895 ;
      VIA 15.01 602.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 602.545 15.78 602.915 ;
      VIA 15.01 602.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 602.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 595.905 15.8 596.235 ;
      VIA 15.01 596.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 595.885 15.78 596.255 ;
      VIA 15.01 596.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 596.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 589.245 15.8 589.575 ;
      VIA 15.01 589.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 589.225 15.78 589.595 ;
      VIA 15.01 589.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 589.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 582.585 15.8 582.915 ;
      VIA 15.01 582.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 582.565 15.78 582.935 ;
      VIA 15.01 582.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 582.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 575.925 15.8 576.255 ;
      VIA 15.01 576.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 575.905 15.78 576.275 ;
      VIA 15.01 576.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 576.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 569.265 15.8 569.595 ;
      VIA 15.01 569.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 569.245 15.78 569.615 ;
      VIA 15.01 569.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 569.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 562.605 15.8 562.935 ;
      VIA 15.01 562.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 562.585 15.78 562.955 ;
      VIA 15.01 562.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 562.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 555.945 15.8 556.275 ;
      VIA 15.01 556.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 555.925 15.78 556.295 ;
      VIA 15.01 556.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 556.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 549.285 15.8 549.615 ;
      VIA 15.01 549.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 549.265 15.78 549.635 ;
      VIA 15.01 549.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 549.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 542.625 15.8 542.955 ;
      VIA 15.01 542.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 542.605 15.78 542.975 ;
      VIA 15.01 542.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 542.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 535.965 15.8 536.295 ;
      VIA 15.01 536.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 535.945 15.78 536.315 ;
      VIA 15.01 536.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 536.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 529.305 15.8 529.635 ;
      VIA 15.01 529.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 529.285 15.78 529.655 ;
      VIA 15.01 529.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 529.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 522.645 15.8 522.975 ;
      VIA 15.01 522.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 522.625 15.78 522.995 ;
      VIA 15.01 522.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 522.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 515.985 15.8 516.315 ;
      VIA 15.01 516.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 515.965 15.78 516.335 ;
      VIA 15.01 516.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 516.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 509.325 15.8 509.655 ;
      VIA 15.01 509.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 509.305 15.78 509.675 ;
      VIA 15.01 509.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 509.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 502.665 15.8 502.995 ;
      VIA 15.01 502.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 502.645 15.78 503.015 ;
      VIA 15.01 502.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 502.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 496.005 15.8 496.335 ;
      VIA 15.01 496.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 495.985 15.78 496.355 ;
      VIA 15.01 496.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 496.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 489.345 15.8 489.675 ;
      VIA 15.01 489.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 489.325 15.78 489.695 ;
      VIA 15.01 489.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 489.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 482.685 15.8 483.015 ;
      VIA 15.01 482.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 482.665 15.78 483.035 ;
      VIA 15.01 482.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 482.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 476.025 15.8 476.355 ;
      VIA 15.01 476.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 476.005 15.78 476.375 ;
      VIA 15.01 476.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 476.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 469.365 15.8 469.695 ;
      VIA 15.01 469.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 469.345 15.78 469.715 ;
      VIA 15.01 469.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 469.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 462.705 15.8 463.035 ;
      VIA 15.01 462.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 462.685 15.78 463.055 ;
      VIA 15.01 462.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 462.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 456.045 15.8 456.375 ;
      VIA 15.01 456.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 456.025 15.78 456.395 ;
      VIA 15.01 456.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 456.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 449.385 15.8 449.715 ;
      VIA 15.01 449.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 449.365 15.78 449.735 ;
      VIA 15.01 449.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 449.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 442.725 15.8 443.055 ;
      VIA 15.01 442.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 442.705 15.78 443.075 ;
      VIA 15.01 442.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 442.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 436.065 15.8 436.395 ;
      VIA 15.01 436.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 436.045 15.78 436.415 ;
      VIA 15.01 436.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 436.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 429.405 15.8 429.735 ;
      VIA 15.01 429.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 429.385 15.78 429.755 ;
      VIA 15.01 429.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 429.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 422.745 15.8 423.075 ;
      VIA 15.01 422.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 422.725 15.78 423.095 ;
      VIA 15.01 422.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 422.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 416.085 15.8 416.415 ;
      VIA 15.01 416.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 416.065 15.78 416.435 ;
      VIA 15.01 416.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 416.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 409.425 15.8 409.755 ;
      VIA 15.01 409.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 409.405 15.78 409.775 ;
      VIA 15.01 409.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 409.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 402.765 15.8 403.095 ;
      VIA 15.01 402.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 402.745 15.78 403.115 ;
      VIA 15.01 402.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 402.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 396.105 15.8 396.435 ;
      VIA 15.01 396.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 396.085 15.78 396.455 ;
      VIA 15.01 396.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 396.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 389.445 15.8 389.775 ;
      VIA 15.01 389.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 389.425 15.78 389.795 ;
      VIA 15.01 389.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 389.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 382.785 15.8 383.115 ;
      VIA 15.01 382.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 382.765 15.78 383.135 ;
      VIA 15.01 382.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 382.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 376.125 15.8 376.455 ;
      VIA 15.01 376.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 376.105 15.78 376.475 ;
      VIA 15.01 376.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 376.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 369.465 15.8 369.795 ;
      VIA 15.01 369.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 369.445 15.78 369.815 ;
      VIA 15.01 369.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 369.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 362.805 15.8 363.135 ;
      VIA 15.01 362.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 362.785 15.78 363.155 ;
      VIA 15.01 362.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 362.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 356.145 15.8 356.475 ;
      VIA 15.01 356.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 356.125 15.78 356.495 ;
      VIA 15.01 356.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 356.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 349.485 15.8 349.815 ;
      VIA 15.01 349.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 349.465 15.78 349.835 ;
      VIA 15.01 349.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 349.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 342.825 15.8 343.155 ;
      VIA 15.01 342.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 342.805 15.78 343.175 ;
      VIA 15.01 342.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 342.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 336.165 15.8 336.495 ;
      VIA 15.01 336.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 336.145 15.78 336.515 ;
      VIA 15.01 336.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 336.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 329.505 15.8 329.835 ;
      VIA 15.01 329.67 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 329.485 15.78 329.855 ;
      VIA 15.01 329.67 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 329.67 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 322.845 15.8 323.175 ;
      VIA 15.01 323.01 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 322.825 15.78 323.195 ;
      VIA 15.01 323.01 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 323.01 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 316.185 15.8 316.515 ;
      VIA 15.01 316.35 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 316.165 15.78 316.535 ;
      VIA 15.01 316.35 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 316.35 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 309.525 15.8 309.855 ;
      VIA 15.01 309.69 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 309.505 15.78 309.875 ;
      VIA 15.01 309.69 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 309.69 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 302.865 15.8 303.195 ;
      VIA 15.01 303.03 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 302.845 15.78 303.215 ;
      VIA 15.01 303.03 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 303.03 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 296.205 15.8 296.535 ;
      VIA 15.01 296.37 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 296.185 15.78 296.555 ;
      VIA 15.01 296.37 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 296.37 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 289.545 15.8 289.875 ;
      VIA 15.01 289.71 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 289.525 15.78 289.895 ;
      VIA 15.01 289.71 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 289.71 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 282.885 15.8 283.215 ;
      VIA 15.01 283.05 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 282.865 15.78 283.235 ;
      VIA 15.01 283.05 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 283.05 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 276.225 15.8 276.555 ;
      VIA 15.01 276.39 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 276.205 15.78 276.575 ;
      VIA 15.01 276.39 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 276.39 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 269.565 15.8 269.895 ;
      VIA 15.01 269.73 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 269.545 15.78 269.915 ;
      VIA 15.01 269.73 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 269.73 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 262.905 15.8 263.235 ;
      VIA 15.01 263.07 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 262.885 15.78 263.255 ;
      VIA 15.01 263.07 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 263.07 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 256.245 15.8 256.575 ;
      VIA 15.01 256.41 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 256.225 15.78 256.595 ;
      VIA 15.01 256.41 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 256.41 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 249.585 15.8 249.915 ;
      VIA 15.01 249.75 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 249.565 15.78 249.935 ;
      VIA 15.01 249.75 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 249.75 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 242.925 15.8 243.255 ;
      VIA 15.01 243.09 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 242.905 15.78 243.275 ;
      VIA 15.01 243.09 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 243.09 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 236.265 15.8 236.595 ;
      VIA 15.01 236.43 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 236.245 15.78 236.615 ;
      VIA 15.01 236.43 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 236.43 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 229.605 15.8 229.935 ;
      VIA 15.01 229.77 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 229.585 15.78 229.955 ;
      VIA 15.01 229.77 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 229.77 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 222.945 15.8 223.275 ;
      VIA 15.01 223.11 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 222.925 15.78 223.295 ;
      VIA 15.01 223.11 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 223.11 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 216.285 15.8 216.615 ;
      VIA 15.01 216.45 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 216.265 15.78 216.635 ;
      VIA 15.01 216.45 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 216.45 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 209.625 15.8 209.955 ;
      VIA 15.01 209.79 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 209.605 15.78 209.975 ;
      VIA 15.01 209.79 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 209.79 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 202.965 15.8 203.295 ;
      VIA 15.01 203.13 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 202.945 15.78 203.315 ;
      VIA 15.01 203.13 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 203.13 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 196.305 15.8 196.635 ;
      VIA 15.01 196.47 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 196.285 15.78 196.655 ;
      VIA 15.01 196.47 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 196.47 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 189.645 15.8 189.975 ;
      VIA 15.01 189.81 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 189.625 15.78 189.995 ;
      VIA 15.01 189.81 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 189.81 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 182.985 15.8 183.315 ;
      VIA 15.01 183.15 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 182.965 15.78 183.335 ;
      VIA 15.01 183.15 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 183.15 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 176.325 15.8 176.655 ;
      VIA 15.01 176.49 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 176.305 15.78 176.675 ;
      VIA 15.01 176.49 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 176.49 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 169.665 15.8 169.995 ;
      VIA 15.01 169.83 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 169.645 15.78 170.015 ;
      VIA 15.01 169.83 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 169.83 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 163.005 15.8 163.335 ;
      VIA 15.01 163.17 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 162.985 15.78 163.355 ;
      VIA 15.01 163.17 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 163.17 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 156.345 15.8 156.675 ;
      VIA 15.01 156.51 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 156.325 15.78 156.695 ;
      VIA 15.01 156.51 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 156.51 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 149.685 15.8 150.015 ;
      VIA 15.01 149.85 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 149.665 15.78 150.035 ;
      VIA 15.01 149.85 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 149.85 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 143.025 15.8 143.355 ;
      VIA 15.01 143.19 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 143.005 15.78 143.375 ;
      VIA 15.01 143.19 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 143.19 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 136.365 15.8 136.695 ;
      VIA 15.01 136.53 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 136.345 15.78 136.715 ;
      VIA 15.01 136.53 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 136.53 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 129.705 15.8 130.035 ;
      VIA 15.01 129.87 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 129.685 15.78 130.055 ;
      VIA 15.01 129.87 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 129.87 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 123.045 15.8 123.375 ;
      VIA 15.01 123.21 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 123.025 15.78 123.395 ;
      VIA 15.01 123.21 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 123.21 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 116.385 15.8 116.715 ;
      VIA 15.01 116.55 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 116.365 15.78 116.735 ;
      VIA 15.01 116.55 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 116.55 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 109.725 15.8 110.055 ;
      VIA 15.01 109.89 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 109.705 15.78 110.075 ;
      VIA 15.01 109.89 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 109.89 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 103.065 15.8 103.395 ;
      VIA 15.01 103.23 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 103.045 15.78 103.415 ;
      VIA 15.01 103.23 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 103.23 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 96.405 15.8 96.735 ;
      VIA 15.01 96.57 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 96.385 15.78 96.755 ;
      VIA 15.01 96.57 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 96.57 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 89.745 15.8 90.075 ;
      VIA 15.01 89.91 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 89.725 15.78 90.095 ;
      VIA 15.01 89.91 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 89.91 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 83.085 15.8 83.415 ;
      VIA 15.01 83.25 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 83.065 15.78 83.435 ;
      VIA 15.01 83.25 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 83.25 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 76.425 15.8 76.755 ;
      VIA 15.01 76.59 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 76.405 15.78 76.775 ;
      VIA 15.01 76.59 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 76.59 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 69.765 15.8 70.095 ;
      VIA 15.01 69.93 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 69.745 15.78 70.115 ;
      VIA 15.01 69.93 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 69.93 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 63.105 15.8 63.435 ;
      VIA 15.01 63.27 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 63.085 15.78 63.455 ;
      VIA 15.01 63.27 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 63.27 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 56.445 15.8 56.775 ;
      VIA 15.01 56.61 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 56.425 15.78 56.795 ;
      VIA 15.01 56.61 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 56.61 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 49.785 15.8 50.115 ;
      VIA 15.01 49.95 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 49.765 15.78 50.135 ;
      VIA 15.01 49.95 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 49.95 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 43.125 15.8 43.455 ;
      VIA 15.01 43.29 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 43.105 15.78 43.475 ;
      VIA 15.01 43.29 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 43.29 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 36.465 15.8 36.795 ;
      VIA 15.01 36.63 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 36.445 15.78 36.815 ;
      VIA 15.01 36.63 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 36.63 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 29.805 15.8 30.135 ;
      VIA 15.01 29.97 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 29.785 15.78 30.155 ;
      VIA 15.01 29.97 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 29.97 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 23.145 15.8 23.475 ;
      VIA 15.01 23.31 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 23.125 15.78 23.495 ;
      VIA 15.01 23.31 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 23.31 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 16.485 15.8 16.815 ;
      VIA 15.01 16.65 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 16.465 15.78 16.835 ;
      VIA 15.01 16.65 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 16.65 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 9.825 15.8 10.155 ;
      VIA 15.01 9.99 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 9.805 15.78 10.175 ;
      VIA 15.01 9.99 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 9.99 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.22 3.165 15.8 3.495 ;
      VIA 15.01 3.33 ibex_ex_block_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.24 3.145 15.78 3.515 ;
      VIA 15.01 3.33 ibex_ex_block_via3_4_1600_480_1_4_400_400 ;
      VIA 15.01 3.33 ibex_ex_block_via2_3_1600_480_1_5_320_320 ;
    END
  END VSS
  PIN alu_adder_result_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 763.9 0.8 764.2 ;
    END
  END alu_adder_result_ex_o[0]
  PIN alu_adder_result_ex_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 763.9 262.08 764.2 ;
    END
  END alu_adder_result_ex_o[10]
  PIN alu_adder_result_ex_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 759.46 262.08 759.76 ;
    END
  END alu_adder_result_ex_o[11]
  PIN alu_adder_result_ex_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 675.1 0.8 675.4 ;
    END
  END alu_adder_result_ex_o[12]
  PIN alu_adder_result_ex_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 657.34 262.08 657.64 ;
    END
  END alu_adder_result_ex_o[13]
  PIN alu_adder_result_ex_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  237.77 781.755 237.91 782.24 ;
    END
  END alu_adder_result_ex_o[14]
  PIN alu_adder_result_ex_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  255.05 781.755 255.19 782.24 ;
    END
  END alu_adder_result_ex_o[15]
  PIN alu_adder_result_ex_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  138.41 781.755 138.55 782.24 ;
    END
  END alu_adder_result_ex_o[16]
  PIN alu_adder_result_ex_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 759.46 0.8 759.76 ;
    END
  END alu_adder_result_ex_o[17]
  PIN alu_adder_result_ex_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 723.94 262.08 724.24 ;
    END
  END alu_adder_result_ex_o[18]
  PIN alu_adder_result_ex_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  142.73 781.755 142.87 782.24 ;
    END
  END alu_adder_result_ex_o[19]
  PIN alu_adder_result_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  125.45 781.755 125.59 782.24 ;
    END
  END alu_adder_result_ex_o[1]
  PIN alu_adder_result_ex_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 715.06 262.08 715.36 ;
    END
  END alu_adder_result_ex_o[20]
  PIN alu_adder_result_ex_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 661.78 262.08 662.08 ;
    END
  END alu_adder_result_ex_o[21]
  PIN alu_adder_result_ex_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 683.98 262.08 684.28 ;
    END
  END alu_adder_result_ex_o[22]
  PIN alu_adder_result_ex_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 639.58 262.08 639.88 ;
    END
  END alu_adder_result_ex_o[23]
  PIN alu_adder_result_ex_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 670.66 262.08 670.96 ;
    END
  END alu_adder_result_ex_o[24]
  PIN alu_adder_result_ex_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 612.94 262.08 613.24 ;
    END
  END alu_adder_result_ex_o[25]
  PIN alu_adder_result_ex_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 630.7 262.08 631 ;
    END
  END alu_adder_result_ex_o[26]
  PIN alu_adder_result_ex_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 621.82 262.08 622.12 ;
    END
  END alu_adder_result_ex_o[27]
  PIN alu_adder_result_ex_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 728.38 262.08 728.68 ;
    END
  END alu_adder_result_ex_o[28]
  PIN alu_adder_result_ex_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 675.1 262.08 675.4 ;
    END
  END alu_adder_result_ex_o[29]
  PIN alu_adder_result_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 377.62 0.8 377.92 ;
    END
  END alu_adder_result_ex_o[2]
  PIN alu_adder_result_ex_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 719.5 262.08 719.8 ;
    END
  END alu_adder_result_ex_o[30]
  PIN alu_adder_result_ex_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 697.3 262.08 697.6 ;
    END
  END alu_adder_result_ex_o[31]
  PIN alu_adder_result_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 755.02 0.8 755.32 ;
    END
  END alu_adder_result_ex_o[3]
  PIN alu_adder_result_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 692.86 262.08 693.16 ;
    END
  END alu_adder_result_ex_o[4]
  PIN alu_adder_result_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 453.1 0.8 453.4 ;
    END
  END alu_adder_result_ex_o[5]
  PIN alu_adder_result_ex_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  116.81 781.755 116.95 782.24 ;
    END
  END alu_adder_result_ex_o[6]
  PIN alu_adder_result_ex_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  121.13 781.755 121.27 782.24 ;
    END
  END alu_adder_result_ex_o[7]
  PIN alu_adder_result_ex_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 755.02 262.08 755.32 ;
    END
  END alu_adder_result_ex_o[8]
  PIN alu_adder_result_ex_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.49 781.755 112.63 782.24 ;
    END
  END alu_adder_result_ex_o[9]
  PIN alu_instr_first_cycle_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 62.38 0.8 62.68 ;
    END
  END alu_instr_first_cycle_i
  PIN alu_operand_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 599.62 0.8 599.92 ;
    END
  END alu_operand_a_i[0]
  PIN alu_operand_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 595.18 0.8 595.48 ;
    END
  END alu_operand_a_i[10]
  PIN alu_operand_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 604.06 0.8 604.36 ;
    END
  END alu_operand_a_i[11]
  PIN alu_operand_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  4.49 781.755 4.63 782.24 ;
    END
  END alu_operand_a_i[12]
  PIN alu_operand_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  52.01 781.755 52.15 782.24 ;
    END
  END alu_operand_a_i[13]
  PIN alu_operand_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  17.45 781.755 17.59 782.24 ;
    END
  END alu_operand_a_i[14]
  PIN alu_operand_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  56.33 781.755 56.47 782.24 ;
    END
  END alu_operand_a_i[15]
  PIN alu_operand_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  60.65 781.755 60.79 782.24 ;
    END
  END alu_operand_a_i[16]
  PIN alu_operand_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  21.77 781.755 21.91 782.24 ;
    END
  END alu_operand_a_i[17]
  PIN alu_operand_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.13 781.755 13.27 782.24 ;
    END
  END alu_operand_a_i[18]
  PIN alu_operand_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  8.81 781.755 8.95 782.24 ;
    END
  END alu_operand_a_i[19]
  PIN alu_operand_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 630.7 0.8 631 ;
    END
  END alu_operand_a_i[1]
  PIN alu_operand_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 621.82 0.8 622.12 ;
    END
  END alu_operand_a_i[20]
  PIN alu_operand_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 719.5 0.8 719.8 ;
    END
  END alu_operand_a_i[21]
  PIN alu_operand_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 710.62 0.8 710.92 ;
    END
  END alu_operand_a_i[22]
  PIN alu_operand_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 568.54 0.8 568.84 ;
    END
  END alu_operand_a_i[23]
  PIN alu_operand_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 670.66 0.8 670.96 ;
    END
  END alu_operand_a_i[24]
  PIN alu_operand_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 639.58 0.8 639.88 ;
    END
  END alu_operand_a_i[25]
  PIN alu_operand_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 683.98 0.8 684.28 ;
    END
  END alu_operand_a_i[26]
  PIN alu_operand_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 555.22 0.8 555.52 ;
    END
  END alu_operand_a_i[27]
  PIN alu_operand_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 541.9 0.8 542.2 ;
    END
  END alu_operand_a_i[28]
  PIN alu_operand_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 732.82 0.8 733.12 ;
    END
  END alu_operand_a_i[29]
  PIN alu_operand_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 750.58 0.8 750.88 ;
    END
  END alu_operand_a_i[2]
  PIN alu_operand_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 723.94 0.8 724.24 ;
    END
  END alu_operand_a_i[30]
  PIN alu_operand_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 626.26 0.8 626.56 ;
    END
  END alu_operand_a_i[31]
  PIN alu_operand_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 697.3 0.8 697.6 ;
    END
  END alu_operand_a_i[3]
  PIN alu_operand_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 728.38 0.8 728.68 ;
    END
  END alu_operand_a_i[4]
  PIN alu_operand_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 688.42 0.8 688.72 ;
    END
  END alu_operand_a_i[5]
  PIN alu_operand_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 679.54 0.8 679.84 ;
    END
  END alu_operand_a_i[6]
  PIN alu_operand_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 564.1 0.8 564.4 ;
    END
  END alu_operand_a_i[7]
  PIN alu_operand_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 586.3 0.8 586.6 ;
    END
  END alu_operand_a_i[8]
  PIN alu_operand_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 577.42 0.8 577.72 ;
    END
  END alu_operand_a_i[9]
  PIN alu_operand_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 657.34 0.8 657.64 ;
    END
  END alu_operand_b_i[0]
  PIN alu_operand_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 572.98 0.8 573.28 ;
    END
  END alu_operand_b_i[10]
  PIN alu_operand_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 559.66 0.8 559.96 ;
    END
  END alu_operand_b_i[11]
  PIN alu_operand_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.25 781.755 82.39 782.24 ;
    END
  END alu_operand_b_i[12]
  PIN alu_operand_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.85 781.755 103.99 782.24 ;
    END
  END alu_operand_b_i[13]
  PIN alu_operand_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.89 781.755 91.03 782.24 ;
    END
  END alu_operand_b_i[14]
  PIN alu_operand_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.97 781.755 65.11 782.24 ;
    END
  END alu_operand_b_i[15]
  PIN alu_operand_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  69.29 781.755 69.43 782.24 ;
    END
  END alu_operand_b_i[16]
  PIN alu_operand_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  95.21 781.755 95.35 782.24 ;
    END
  END alu_operand_b_i[17]
  PIN alu_operand_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.53 781.755 99.67 782.24 ;
    END
  END alu_operand_b_i[18]
  PIN alu_operand_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.61 781.755 73.75 782.24 ;
    END
  END alu_operand_b_i[19]
  PIN alu_operand_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 390.94 0.8 391.24 ;
    END
  END alu_operand_b_i[1]
  PIN alu_operand_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 612.94 0.8 613.24 ;
    END
  END alu_operand_b_i[20]
  PIN alu_operand_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 661.78 0.8 662.08 ;
    END
  END alu_operand_b_i[21]
  PIN alu_operand_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.17 781.755 108.31 782.24 ;
    END
  END alu_operand_b_i[22]
  PIN alu_operand_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 706.18 0.8 706.48 ;
    END
  END alu_operand_b_i[23]
  PIN alu_operand_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 608.5 0.8 608.8 ;
    END
  END alu_operand_b_i[24]
  PIN alu_operand_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 519.7 0.8 520 ;
    END
  END alu_operand_b_i[25]
  PIN alu_operand_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 524.14 0.8 524.44 ;
    END
  END alu_operand_b_i[26]
  PIN alu_operand_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 533.02 0.8 533.32 ;
    END
  END alu_operand_b_i[27]
  PIN alu_operand_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 546.34 0.8 546.64 ;
    END
  END alu_operand_b_i[28]
  PIN alu_operand_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 537.46 0.8 537.76 ;
    END
  END alu_operand_b_i[29]
  PIN alu_operand_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 97.9 0.8 98.2 ;
    END
  END alu_operand_b_i[2]
  PIN alu_operand_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 550.78 0.8 551.08 ;
    END
  END alu_operand_b_i[30]
  PIN alu_operand_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 652.9 0.8 653.2 ;
    END
  END alu_operand_b_i[31]
  PIN alu_operand_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 128.98 0.8 129.28 ;
    END
  END alu_operand_b_i[3]
  PIN alu_operand_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 666.22 0.8 666.52 ;
    END
  END alu_operand_b_i[4]
  PIN alu_operand_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 346.54 0.8 346.84 ;
    END
  END alu_operand_b_i[5]
  PIN alu_operand_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 426.46 0.8 426.76 ;
    END
  END alu_operand_b_i[6]
  PIN alu_operand_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 635.14 0.8 635.44 ;
    END
  END alu_operand_b_i[7]
  PIN alu_operand_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  77.93 781.755 78.07 782.24 ;
    END
  END alu_operand_b_i[8]
  PIN alu_operand_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  86.57 781.755 86.71 782.24 ;
    END
  END alu_operand_b_i[9]
  PIN alu_operator_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  30.41 781.755 30.55 782.24 ;
    END
  END alu_operator_i[0]
  PIN alu_operator_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  26.09 781.755 26.23 782.24 ;
    END
  END alu_operator_i[1]
  PIN alu_operator_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  39.05 781.755 39.19 782.24 ;
    END
  END alu_operator_i[2]
  PIN alu_operator_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  34.73 781.755 34.87 782.24 ;
    END
  END alu_operator_i[3]
  PIN alu_operator_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  47.69 781.755 47.83 782.24 ;
    END
  END alu_operator_i[4]
  PIN alu_operator_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  43.37 781.755 43.51 782.24 ;
    END
  END alu_operator_i[5]
  PIN branch_decision_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  250.73 781.755 250.87 782.24 ;
    END
  END branch_decision_o
  PIN branch_target_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  242.09 781.755 242.23 782.24 ;
    END
  END branch_target_o[0]
  PIN branch_target_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  129.77 781.755 129.91 782.24 ;
    END
  END branch_target_o[10]
  PIN branch_target_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  172.97 781.755 173.11 782.24 ;
    END
  END branch_target_o[11]
  PIN branch_target_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  134.09 781.755 134.23 782.24 ;
    END
  END branch_target_o[12]
  PIN branch_target_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  185.93 781.755 186.07 782.24 ;
    END
  END branch_target_o[13]
  PIN branch_target_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  177.29 781.755 177.43 782.24 ;
    END
  END branch_target_o[14]
  PIN branch_target_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  164.33 781.755 164.47 782.24 ;
    END
  END branch_target_o[15]
  PIN branch_target_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  160.01 781.755 160.15 782.24 ;
    END
  END branch_target_o[16]
  PIN branch_target_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  181.61 781.755 181.75 782.24 ;
    END
  END branch_target_o[17]
  PIN branch_target_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  155.69 781.755 155.83 782.24 ;
    END
  END branch_target_o[18]
  PIN branch_target_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.37 781.755 151.51 782.24 ;
    END
  END branch_target_o[19]
  PIN branch_target_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 479.74 0.8 480.04 ;
    END
  END branch_target_o[1]
  PIN branch_target_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  220.49 781.755 220.63 782.24 ;
    END
  END branch_target_o[20]
  PIN branch_target_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  168.65 781.755 168.79 782.24 ;
    END
  END branch_target_o[21]
  PIN branch_target_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  216.17 781.755 216.31 782.24 ;
    END
  END branch_target_o[22]
  PIN branch_target_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  198.89 781.755 199.03 782.24 ;
    END
  END branch_target_o[23]
  PIN branch_target_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  194.57 781.755 194.71 782.24 ;
    END
  END branch_target_o[24]
  PIN branch_target_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  246.41 781.755 246.55 782.24 ;
    END
  END branch_target_o[25]
  PIN branch_target_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  190.25 781.755 190.39 782.24 ;
    END
  END branch_target_o[26]
  PIN branch_target_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  233.45 781.755 233.59 782.24 ;
    END
  END branch_target_o[27]
  PIN branch_target_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  229.13 781.755 229.27 782.24 ;
    END
  END branch_target_o[28]
  PIN branch_target_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  203.21 781.755 203.35 782.24 ;
    END
  END branch_target_o[29]
  PIN branch_target_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 49.06 0.8 49.36 ;
    END
  END branch_target_o[2]
  PIN branch_target_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  211.85 781.755 211.99 782.24 ;
    END
  END branch_target_o[30]
  PIN branch_target_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  207.53 781.755 207.67 782.24 ;
    END
  END branch_target_o[31]
  PIN branch_target_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 177.82 0.8 178.12 ;
    END
  END branch_target_o[3]
  PIN branch_target_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  224.81 781.755 224.95 782.24 ;
    END
  END branch_target_o[4]
  PIN branch_target_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 444.22 0.8 444.52 ;
    END
  END branch_target_o[5]
  PIN branch_target_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  147.05 781.755 147.19 782.24 ;
    END
  END branch_target_o[6]
  PIN branch_target_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 688.42 262.08 688.72 ;
    END
  END branch_target_o[7]
  PIN branch_target_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 666.22 262.08 666.52 ;
    END
  END branch_target_o[8]
  PIN branch_target_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 635.14 262.08 635.44 ;
    END
  END branch_target_o[9]
  PIN bt_a_operand_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  4.49 0 4.63 0.485 ;
    END
  END bt_a_operand_i[0]
  PIN bt_a_operand_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  8.81 0 8.95 0.485 ;
    END
  END bt_a_operand_i[10]
  PIN bt_a_operand_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.13 0 13.27 0.485 ;
    END
  END bt_a_operand_i[11]
  PIN bt_a_operand_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  17.45 0 17.59 0.485 ;
    END
  END bt_a_operand_i[12]
  PIN bt_a_operand_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  21.77 0 21.91 0.485 ;
    END
  END bt_a_operand_i[13]
  PIN bt_a_operand_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  26.09 0 26.23 0.485 ;
    END
  END bt_a_operand_i[14]
  PIN bt_a_operand_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  30.41 0 30.55 0.485 ;
    END
  END bt_a_operand_i[15]
  PIN bt_a_operand_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  34.73 0 34.87 0.485 ;
    END
  END bt_a_operand_i[16]
  PIN bt_a_operand_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  39.05 0 39.19 0.485 ;
    END
  END bt_a_operand_i[17]
  PIN bt_a_operand_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  43.37 0 43.51 0.485 ;
    END
  END bt_a_operand_i[18]
  PIN bt_a_operand_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  47.69 0 47.83 0.485 ;
    END
  END bt_a_operand_i[19]
  PIN bt_a_operand_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  52.01 0 52.15 0.485 ;
    END
  END bt_a_operand_i[1]
  PIN bt_a_operand_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  56.33 0 56.47 0.485 ;
    END
  END bt_a_operand_i[20]
  PIN bt_a_operand_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  60.65 0 60.79 0.485 ;
    END
  END bt_a_operand_i[21]
  PIN bt_a_operand_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.97 0 65.11 0.485 ;
    END
  END bt_a_operand_i[22]
  PIN bt_a_operand_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  69.29 0 69.43 0.485 ;
    END
  END bt_a_operand_i[23]
  PIN bt_a_operand_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.61 0 73.75 0.485 ;
    END
  END bt_a_operand_i[24]
  PIN bt_a_operand_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  77.93 0 78.07 0.485 ;
    END
  END bt_a_operand_i[25]
  PIN bt_a_operand_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.25 0 82.39 0.485 ;
    END
  END bt_a_operand_i[26]
  PIN bt_a_operand_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  86.57 0 86.71 0.485 ;
    END
  END bt_a_operand_i[27]
  PIN bt_a_operand_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.89 0 91.03 0.485 ;
    END
  END bt_a_operand_i[28]
  PIN bt_a_operand_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  95.21 0 95.35 0.485 ;
    END
  END bt_a_operand_i[29]
  PIN bt_a_operand_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.53 0 99.67 0.485 ;
    END
  END bt_a_operand_i[2]
  PIN bt_a_operand_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.85 0 103.99 0.485 ;
    END
  END bt_a_operand_i[30]
  PIN bt_a_operand_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.17 0 108.31 0.485 ;
    END
  END bt_a_operand_i[31]
  PIN bt_a_operand_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.49 0 112.63 0.485 ;
    END
  END bt_a_operand_i[3]
  PIN bt_a_operand_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  116.81 0 116.95 0.485 ;
    END
  END bt_a_operand_i[4]
  PIN bt_a_operand_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  121.13 0 121.27 0.485 ;
    END
  END bt_a_operand_i[5]
  PIN bt_a_operand_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  125.45 0 125.59 0.485 ;
    END
  END bt_a_operand_i[6]
  PIN bt_a_operand_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  129.77 0 129.91 0.485 ;
    END
  END bt_a_operand_i[7]
  PIN bt_a_operand_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  134.09 0 134.23 0.485 ;
    END
  END bt_a_operand_i[8]
  PIN bt_a_operand_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  138.41 0 138.55 0.485 ;
    END
  END bt_a_operand_i[9]
  PIN bt_b_operand_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  142.73 0 142.87 0.485 ;
    END
  END bt_b_operand_i[0]
  PIN bt_b_operand_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  147.05 0 147.19 0.485 ;
    END
  END bt_b_operand_i[10]
  PIN bt_b_operand_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.37 0 151.51 0.485 ;
    END
  END bt_b_operand_i[11]
  PIN bt_b_operand_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  155.69 0 155.83 0.485 ;
    END
  END bt_b_operand_i[12]
  PIN bt_b_operand_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  160.01 0 160.15 0.485 ;
    END
  END bt_b_operand_i[13]
  PIN bt_b_operand_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  164.33 0 164.47 0.485 ;
    END
  END bt_b_operand_i[14]
  PIN bt_b_operand_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  168.65 0 168.79 0.485 ;
    END
  END bt_b_operand_i[15]
  PIN bt_b_operand_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  172.97 0 173.11 0.485 ;
    END
  END bt_b_operand_i[16]
  PIN bt_b_operand_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  177.29 0 177.43 0.485 ;
    END
  END bt_b_operand_i[17]
  PIN bt_b_operand_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  181.61 0 181.75 0.485 ;
    END
  END bt_b_operand_i[18]
  PIN bt_b_operand_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  185.93 0 186.07 0.485 ;
    END
  END bt_b_operand_i[19]
  PIN bt_b_operand_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  190.25 0 190.39 0.485 ;
    END
  END bt_b_operand_i[1]
  PIN bt_b_operand_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  194.57 0 194.71 0.485 ;
    END
  END bt_b_operand_i[20]
  PIN bt_b_operand_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  198.89 0 199.03 0.485 ;
    END
  END bt_b_operand_i[21]
  PIN bt_b_operand_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  203.21 0 203.35 0.485 ;
    END
  END bt_b_operand_i[22]
  PIN bt_b_operand_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  207.53 0 207.67 0.485 ;
    END
  END bt_b_operand_i[23]
  PIN bt_b_operand_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  211.85 0 211.99 0.485 ;
    END
  END bt_b_operand_i[24]
  PIN bt_b_operand_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  216.17 0 216.31 0.485 ;
    END
  END bt_b_operand_i[25]
  PIN bt_b_operand_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  220.49 0 220.63 0.485 ;
    END
  END bt_b_operand_i[26]
  PIN bt_b_operand_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  224.81 0 224.95 0.485 ;
    END
  END bt_b_operand_i[27]
  PIN bt_b_operand_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  229.13 0 229.27 0.485 ;
    END
  END bt_b_operand_i[28]
  PIN bt_b_operand_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  233.45 0 233.59 0.485 ;
    END
  END bt_b_operand_i[29]
  PIN bt_b_operand_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  237.77 0 237.91 0.485 ;
    END
  END bt_b_operand_i[2]
  PIN bt_b_operand_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  242.09 0 242.23 0.485 ;
    END
  END bt_b_operand_i[30]
  PIN bt_b_operand_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  246.41 0 246.55 0.485 ;
    END
  END bt_b_operand_i[31]
  PIN bt_b_operand_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  250.73 0 250.87 0.485 ;
    END
  END bt_b_operand_i[3]
  PIN bt_b_operand_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  255.05 0 255.19 0.485 ;
    END
  END bt_b_operand_i[4]
  PIN bt_b_operand_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 4.66 262.08 4.96 ;
    END
  END bt_b_operand_i[5]
  PIN bt_b_operand_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 9.1 262.08 9.4 ;
    END
  END bt_b_operand_i[6]
  PIN bt_b_operand_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 13.54 262.08 13.84 ;
    END
  END bt_b_operand_i[7]
  PIN bt_b_operand_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 17.98 262.08 18.28 ;
    END
  END bt_b_operand_i[8]
  PIN bt_b_operand_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 22.42 262.08 22.72 ;
    END
  END bt_b_operand_i[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 608.5 262.08 608.8 ;
    END
  END clk_i
  PIN data_ind_timing_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 701.74 262.08 702.04 ;
    END
  END data_ind_timing_i
  PIN div_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 408.7 262.08 409 ;
    END
  END div_en_i
  PIN div_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 115.66 262.08 115.96 ;
    END
  END div_sel_i
  PIN ex_valid_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 226.66 262.08 226.96 ;
    END
  END ex_valid_o
  PIN imd_val_d_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 319.9 0.8 320.2 ;
    END
  END imd_val_d_o[0]
  PIN imd_val_d_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 448.66 0.8 448.96 ;
    END
  END imd_val_d_o[10]
  PIN imd_val_d_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 466.42 0.8 466.72 ;
    END
  END imd_val_d_o[11]
  PIN imd_val_d_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 457.54 0.8 457.84 ;
    END
  END imd_val_d_o[12]
  PIN imd_val_d_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 439.78 0.8 440.08 ;
    END
  END imd_val_d_o[13]
  PIN imd_val_d_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 617.38 0.8 617.68 ;
    END
  END imd_val_d_o[14]
  PIN imd_val_d_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 262.18 0.8 262.48 ;
    END
  END imd_val_d_o[15]
  PIN imd_val_d_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 315.46 0.8 315.76 ;
    END
  END imd_val_d_o[16]
  PIN imd_val_d_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 417.58 0.8 417.88 ;
    END
  END imd_val_d_o[17]
  PIN imd_val_d_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 266.62 0.8 266.92 ;
    END
  END imd_val_d_o[18]
  PIN imd_val_d_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 115.66 0.8 115.96 ;
    END
  END imd_val_d_o[19]
  PIN imd_val_d_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 746.14 0.8 746.44 ;
    END
  END imd_val_d_o[1]
  PIN imd_val_d_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 248.86 0.8 249.16 ;
    END
  END imd_val_d_o[20]
  PIN imd_val_d_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 182.26 0.8 182.56 ;
    END
  END imd_val_d_o[21]
  PIN imd_val_d_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 133.42 0.8 133.72 ;
    END
  END imd_val_d_o[22]
  PIN imd_val_d_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 200.02 0.8 200.32 ;
    END
  END imd_val_d_o[23]
  PIN imd_val_d_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 217.78 0.8 218.08 ;
    END
  END imd_val_d_o[24]
  PIN imd_val_d_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 106.78 0.8 107.08 ;
    END
  END imd_val_d_o[25]
  PIN imd_val_d_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 306.58 0.8 306.88 ;
    END
  END imd_val_d_o[26]
  PIN imd_val_d_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 146.74 262.08 147.04 ;
    END
  END imd_val_d_o[27]
  PIN imd_val_d_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 244.42 0.8 244.72 ;
    END
  END imd_val_d_o[28]
  PIN imd_val_d_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 35.74 0.8 36.04 ;
    END
  END imd_val_d_o[29]
  PIN imd_val_d_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 173.38 0.8 173.68 ;
    END
  END imd_val_d_o[2]
  PIN imd_val_d_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 390.94 262.08 391.24 ;
    END
  END imd_val_d_o[30]
  PIN imd_val_d_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 377.62 262.08 377.92 ;
    END
  END imd_val_d_o[31]
  PIN imd_val_d_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 737.26 262.08 737.56 ;
    END
  END imd_val_d_o[32]
  PIN imd_val_d_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 732.82 262.08 733.12 ;
    END
  END imd_val_d_o[33]
  PIN imd_val_d_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 404.26 262.08 404.56 ;
    END
  END imd_val_d_o[34]
  PIN imd_val_d_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 488.62 262.08 488.92 ;
    END
  END imd_val_d_o[35]
  PIN imd_val_d_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 461.98 262.08 462.28 ;
    END
  END imd_val_d_o[36]
  PIN imd_val_d_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 546.34 262.08 546.64 ;
    END
  END imd_val_d_o[37]
  PIN imd_val_d_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 750.58 262.08 750.88 ;
    END
  END imd_val_d_o[38]
  PIN imd_val_d_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 555.22 262.08 555.52 ;
    END
  END imd_val_d_o[39]
  PIN imd_val_d_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 253.3 0.8 253.6 ;
    END
  END imd_val_d_o[3]
  PIN imd_val_d_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 741.7 262.08 742 ;
    END
  END imd_val_d_o[40]
  PIN imd_val_d_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 604.06 262.08 604.36 ;
    END
  END imd_val_d_o[41]
  PIN imd_val_d_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 541.9 262.08 542.2 ;
    END
  END imd_val_d_o[42]
  PIN imd_val_d_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 550.78 262.08 551.08 ;
    END
  END imd_val_d_o[43]
  PIN imd_val_d_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 590.74 262.08 591.04 ;
    END
  END imd_val_d_o[44]
  PIN imd_val_d_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 710.62 262.08 710.92 ;
    END
  END imd_val_d_o[45]
  PIN imd_val_d_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 559.66 262.08 559.96 ;
    END
  END imd_val_d_o[46]
  PIN imd_val_d_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 537.46 262.08 537.76 ;
    END
  END imd_val_d_o[47]
  PIN imd_val_d_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 568.54 262.08 568.84 ;
    END
  END imd_val_d_o[48]
  PIN imd_val_d_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 746.14 262.08 746.44 ;
    END
  END imd_val_d_o[49]
  PIN imd_val_d_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 239.98 0.8 240.28 ;
    END
  END imd_val_d_o[4]
  PIN imd_val_d_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 595.18 262.08 595.48 ;
    END
  END imd_val_d_o[50]
  PIN imd_val_d_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 599.62 262.08 599.92 ;
    END
  END imd_val_d_o[51]
  PIN imd_val_d_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 572.98 262.08 573.28 ;
    END
  END imd_val_d_o[52]
  PIN imd_val_d_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 644.02 262.08 644.32 ;
    END
  END imd_val_d_o[53]
  PIN imd_val_d_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 519.7 262.08 520 ;
    END
  END imd_val_d_o[54]
  PIN imd_val_d_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 577.42 262.08 577.72 ;
    END
  END imd_val_d_o[55]
  PIN imd_val_d_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 581.86 262.08 582.16 ;
    END
  END imd_val_d_o[56]
  PIN imd_val_d_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 626.26 262.08 626.56 ;
    END
  END imd_val_d_o[57]
  PIN imd_val_d_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 515.26 262.08 515.56 ;
    END
  END imd_val_d_o[58]
  PIN imd_val_d_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 479.74 262.08 480.04 ;
    END
  END imd_val_d_o[59]
  PIN imd_val_d_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 22.42 0.8 22.72 ;
    END
  END imd_val_d_o[5]
  PIN imd_val_d_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 435.34 262.08 435.64 ;
    END
  END imd_val_d_o[60]
  PIN imd_val_d_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 497.5 262.08 497.8 ;
    END
  END imd_val_d_o[61]
  PIN imd_val_d_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 506.38 262.08 506.68 ;
    END
  END imd_val_d_o[62]
  PIN imd_val_d_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 470.86 262.08 471.16 ;
    END
  END imd_val_d_o[63]
  PIN imd_val_d_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 528.58 262.08 528.88 ;
    END
  END imd_val_d_o[64]
  PIN imd_val_d_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 679.54 262.08 679.84 ;
    END
  END imd_val_d_o[65]
  PIN imd_val_d_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 235.54 262.08 235.84 ;
    END
  END imd_val_d_o[66]
  PIN imd_val_d_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 239.98 262.08 240.28 ;
    END
  END imd_val_d_o[67]
  PIN imd_val_d_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 413.14 0.8 413.44 ;
    END
  END imd_val_d_o[6]
  PIN imd_val_d_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 9.1 0.8 9.4 ;
    END
  END imd_val_d_o[7]
  PIN imd_val_d_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 284.38 0.8 284.68 ;
    END
  END imd_val_d_o[8]
  PIN imd_val_d_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 777.22 0.8 777.52 ;
    END
  END imd_val_d_o[9]
  PIN imd_val_q_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 235.54 0.8 235.84 ;
    END
  END imd_val_q_i[0]
  PIN imd_val_q_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 648.46 0.8 648.76 ;
    END
  END imd_val_q_i[10]
  PIN imd_val_q_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 768.34 0.8 768.64 ;
    END
  END imd_val_q_i[11]
  PIN imd_val_q_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 644.02 0.8 644.32 ;
    END
  END imd_val_q_i[12]
  PIN imd_val_q_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 737.26 0.8 737.56 ;
    END
  END imd_val_q_i[13]
  PIN imd_val_q_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 435.34 0.8 435.64 ;
    END
  END imd_val_q_i[14]
  PIN imd_val_q_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 399.82 0.8 400.12 ;
    END
  END imd_val_q_i[15]
  PIN imd_val_q_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 404.26 0.8 404.56 ;
    END
  END imd_val_q_i[16]
  PIN imd_val_q_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 422.02 0.8 422.32 ;
    END
  END imd_val_q_i[17]
  PIN imd_val_q_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 257.74 0.8 258.04 ;
    END
  END imd_val_q_i[18]
  PIN imd_val_q_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 57.94 0.8 58.24 ;
    END
  END imd_val_q_i[19]
  PIN imd_val_q_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 430.9 0.8 431.2 ;
    END
  END imd_val_q_i[1]
  PIN imd_val_q_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 84.58 0.8 84.88 ;
    END
  END imd_val_q_i[20]
  PIN imd_val_q_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 231.1 0.8 231.4 ;
    END
  END imd_val_q_i[21]
  PIN imd_val_q_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 302.14 0.8 302.44 ;
    END
  END imd_val_q_i[22]
  PIN imd_val_q_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 226.66 0.8 226.96 ;
    END
  END imd_val_q_i[23]
  PIN imd_val_q_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 137.86 0.8 138.16 ;
    END
  END imd_val_q_i[24]
  PIN imd_val_q_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 26.86 0.8 27.16 ;
    END
  END imd_val_q_i[25]
  PIN imd_val_q_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 293.26 0.8 293.56 ;
    END
  END imd_val_q_i[26]
  PIN imd_val_q_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 364.3 262.08 364.6 ;
    END
  END imd_val_q_i[27]
  PIN imd_val_q_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 324.34 0.8 324.64 ;
    END
  END imd_val_q_i[28]
  PIN imd_val_q_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 328.78 0.8 329.08 ;
    END
  END imd_val_q_i[29]
  PIN imd_val_q_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 271.06 0.8 271.36 ;
    END
  END imd_val_q_i[2]
  PIN imd_val_q_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 399.82 262.08 400.12 ;
    END
  END imd_val_q_i[30]
  PIN imd_val_q_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 652.9 262.08 653.2 ;
    END
  END imd_val_q_i[31]
  PIN imd_val_q_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 26.86 262.08 27.16 ;
    END
  END imd_val_q_i[32]
  PIN imd_val_q_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 31.3 262.08 31.6 ;
    END
  END imd_val_q_i[33]
  PIN imd_val_q_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 315.46 262.08 315.76 ;
    END
  END imd_val_q_i[34]
  PIN imd_val_q_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 31.3 0.8 31.6 ;
    END
  END imd_val_q_i[35]
  PIN imd_val_q_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 279.94 0.8 280.24 ;
    END
  END imd_val_q_i[36]
  PIN imd_val_q_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 208.9 0.8 209.2 ;
    END
  END imd_val_q_i[37]
  PIN imd_val_q_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 297.7 0.8 298 ;
    END
  END imd_val_q_i[38]
  PIN imd_val_q_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 164.5 0.8 164.8 ;
    END
  END imd_val_q_i[39]
  PIN imd_val_q_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 168.94 0.8 169.24 ;
    END
  END imd_val_q_i[3]
  PIN imd_val_q_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 191.14 0.8 191.44 ;
    END
  END imd_val_q_i[40]
  PIN imd_val_q_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 275.5 0.8 275.8 ;
    END
  END imd_val_q_i[41]
  PIN imd_val_q_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 213.34 0.8 213.64 ;
    END
  END imd_val_q_i[42]
  PIN imd_val_q_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 4.66 0.8 4.96 ;
    END
  END imd_val_q_i[43]
  PIN imd_val_q_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 13.54 0.8 13.84 ;
    END
  END imd_val_q_i[44]
  PIN imd_val_q_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 160.06 0.8 160.36 ;
    END
  END imd_val_q_i[45]
  PIN imd_val_q_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 146.74 0.8 147.04 ;
    END
  END imd_val_q_i[46]
  PIN imd_val_q_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 706.18 262.08 706.48 ;
    END
  END imd_val_q_i[47]
  PIN imd_val_q_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 581.86 0.8 582.16 ;
    END
  END imd_val_q_i[48]
  PIN imd_val_q_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 648.46 262.08 648.76 ;
    END
  END imd_val_q_i[49]
  PIN imd_val_q_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 151.18 0.8 151.48 ;
    END
  END imd_val_q_i[4]
  PIN imd_val_q_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 311.02 262.08 311.32 ;
    END
  END imd_val_q_i[50]
  PIN imd_val_q_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 319.9 262.08 320.2 ;
    END
  END imd_val_q_i[51]
  PIN imd_val_q_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 248.86 262.08 249.16 ;
    END
  END imd_val_q_i[52]
  PIN imd_val_q_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 142.3 0.8 142.6 ;
    END
  END imd_val_q_i[53]
  PIN imd_val_q_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 271.06 262.08 271.36 ;
    END
  END imd_val_q_i[54]
  PIN imd_val_q_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 257.74 262.08 258.04 ;
    END
  END imd_val_q_i[55]
  PIN imd_val_q_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 262.18 262.08 262.48 ;
    END
  END imd_val_q_i[56]
  PIN imd_val_q_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 284.38 262.08 284.68 ;
    END
  END imd_val_q_i[57]
  PIN imd_val_q_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 275.5 262.08 275.8 ;
    END
  END imd_val_q_i[58]
  PIN imd_val_q_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 293.26 262.08 293.56 ;
    END
  END imd_val_q_i[59]
  PIN imd_val_q_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 71.26 0.8 71.56 ;
    END
  END imd_val_q_i[5]
  PIN imd_val_q_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 279.94 262.08 280.24 ;
    END
  END imd_val_q_i[60]
  PIN imd_val_q_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 297.7 262.08 298 ;
    END
  END imd_val_q_i[61]
  PIN imd_val_q_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 288.82 262.08 289.12 ;
    END
  END imd_val_q_i[62]
  PIN imd_val_q_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 266.62 262.08 266.92 ;
    END
  END imd_val_q_i[63]
  PIN imd_val_q_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 253.3 262.08 253.6 ;
    END
  END imd_val_q_i[64]
  PIN imd_val_q_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 586.3 262.08 586.6 ;
    END
  END imd_val_q_i[65]
  PIN imd_val_q_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 302.14 262.08 302.44 ;
    END
  END imd_val_q_i[66]
  PIN imd_val_q_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 306.58 262.08 306.88 ;
    END
  END imd_val_q_i[67]
  PIN imd_val_q_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 408.7 0.8 409 ;
    END
  END imd_val_q_i[6]
  PIN imd_val_q_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 311.02 0.8 311.32 ;
    END
  END imd_val_q_i[7]
  PIN imd_val_q_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 155.62 0.8 155.92 ;
    END
  END imd_val_q_i[8]
  PIN imd_val_q_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 772.78 0.8 773.08 ;
    END
  END imd_val_q_i[9]
  PIN imd_val_we_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 386.5 262.08 386.8 ;
    END
  END imd_val_we_o[0]
  PIN imd_val_we_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 382.06 262.08 382.36 ;
    END
  END imd_val_we_o[1]
  PIN mult_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 244.42 262.08 244.72 ;
    END
  END mult_en_i
  PIN mult_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 89.02 0.8 89.32 ;
    END
  END mult_sel_i
  PIN multdiv_operand_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 186.7 262.08 187 ;
    END
  END multdiv_operand_a_i[0]
  PIN multdiv_operand_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 168.94 262.08 169.24 ;
    END
  END multdiv_operand_a_i[10]
  PIN multdiv_operand_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 155.62 262.08 155.92 ;
    END
  END multdiv_operand_a_i[11]
  PIN multdiv_operand_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 124.54 262.08 124.84 ;
    END
  END multdiv_operand_a_i[12]
  PIN multdiv_operand_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 422.02 262.08 422.32 ;
    END
  END multdiv_operand_a_i[13]
  PIN multdiv_operand_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 426.46 262.08 426.76 ;
    END
  END multdiv_operand_a_i[14]
  PIN multdiv_operand_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 173.38 262.08 173.68 ;
    END
  END multdiv_operand_a_i[15]
  PIN multdiv_operand_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 359.86 262.08 360.16 ;
    END
  END multdiv_operand_a_i[16]
  PIN multdiv_operand_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 417.58 262.08 417.88 ;
    END
  END multdiv_operand_a_i[17]
  PIN multdiv_operand_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 128.98 262.08 129.28 ;
    END
  END multdiv_operand_a_i[18]
  PIN multdiv_operand_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 133.42 262.08 133.72 ;
    END
  END multdiv_operand_a_i[19]
  PIN multdiv_operand_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 413.14 262.08 413.44 ;
    END
  END multdiv_operand_a_i[1]
  PIN multdiv_operand_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 177.82 262.08 178.12 ;
    END
  END multdiv_operand_a_i[20]
  PIN multdiv_operand_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 204.46 262.08 204.76 ;
    END
  END multdiv_operand_a_i[21]
  PIN multdiv_operand_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 195.58 262.08 195.88 ;
    END
  END multdiv_operand_a_i[22]
  PIN multdiv_operand_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 217.78 262.08 218.08 ;
    END
  END multdiv_operand_a_i[23]
  PIN multdiv_operand_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 342.1 262.08 342.4 ;
    END
  END multdiv_operand_a_i[24]
  PIN multdiv_operand_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 191.14 262.08 191.44 ;
    END
  END multdiv_operand_a_i[25]
  PIN multdiv_operand_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 160.06 262.08 160.36 ;
    END
  END multdiv_operand_a_i[26]
  PIN multdiv_operand_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 151.18 262.08 151.48 ;
    END
  END multdiv_operand_a_i[27]
  PIN multdiv_operand_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 120.1 262.08 120.4 ;
    END
  END multdiv_operand_a_i[28]
  PIN multdiv_operand_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 137.86 262.08 138.16 ;
    END
  END multdiv_operand_a_i[29]
  PIN multdiv_operand_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 373.18 262.08 373.48 ;
    END
  END multdiv_operand_a_i[2]
  PIN multdiv_operand_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 368.74 262.08 369.04 ;
    END
  END multdiv_operand_a_i[30]
  PIN multdiv_operand_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 164.5 262.08 164.8 ;
    END
  END multdiv_operand_a_i[31]
  PIN multdiv_operand_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 142.3 262.08 142.6 ;
    END
  END multdiv_operand_a_i[3]
  PIN multdiv_operand_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 182.26 262.08 182.56 ;
    END
  END multdiv_operand_a_i[4]
  PIN multdiv_operand_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 208.9 262.08 209.2 ;
    END
  END multdiv_operand_a_i[5]
  PIN multdiv_operand_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 200.02 262.08 200.32 ;
    END
  END multdiv_operand_a_i[6]
  PIN multdiv_operand_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 222.22 262.08 222.52 ;
    END
  END multdiv_operand_a_i[7]
  PIN multdiv_operand_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 346.54 262.08 346.84 ;
    END
  END multdiv_operand_a_i[8]
  PIN multdiv_operand_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 355.42 262.08 355.72 ;
    END
  END multdiv_operand_a_i[9]
  PIN multdiv_operand_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 337.66 0.8 337.96 ;
    END
  END multdiv_operand_b_i[0]
  PIN multdiv_operand_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 350.98 0.8 351.28 ;
    END
  END multdiv_operand_b_i[10]
  PIN multdiv_operand_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 359.86 0.8 360.16 ;
    END
  END multdiv_operand_b_i[11]
  PIN multdiv_operand_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 368.74 0.8 369.04 ;
    END
  END multdiv_operand_b_i[12]
  PIN multdiv_operand_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 364.3 0.8 364.6 ;
    END
  END multdiv_operand_b_i[13]
  PIN multdiv_operand_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 386.5 0.8 386.8 ;
    END
  END multdiv_operand_b_i[14]
  PIN multdiv_operand_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 231.1 262.08 231.4 ;
    END
  END multdiv_operand_b_i[15]
  PIN multdiv_operand_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 342.1 0.8 342.4 ;
    END
  END multdiv_operand_b_i[16]
  PIN multdiv_operand_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 395.38 0.8 395.68 ;
    END
  END multdiv_operand_b_i[17]
  PIN multdiv_operand_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 373.18 0.8 373.48 ;
    END
  END multdiv_operand_b_i[18]
  PIN multdiv_operand_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 102.34 0.8 102.64 ;
    END
  END multdiv_operand_b_i[19]
  PIN multdiv_operand_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 40.18 0.8 40.48 ;
    END
  END multdiv_operand_b_i[1]
  PIN multdiv_operand_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 80.14 0.8 80.44 ;
    END
  END multdiv_operand_b_i[20]
  PIN multdiv_operand_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 195.58 0.8 195.88 ;
    END
  END multdiv_operand_b_i[21]
  PIN multdiv_operand_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 53.5 0.8 53.8 ;
    END
  END multdiv_operand_b_i[22]
  PIN multdiv_operand_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 288.82 0.8 289.12 ;
    END
  END multdiv_operand_b_i[23]
  PIN multdiv_operand_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 222.22 0.8 222.52 ;
    END
  END multdiv_operand_b_i[24]
  PIN multdiv_operand_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 93.46 0.8 93.76 ;
    END
  END multdiv_operand_b_i[25]
  PIN multdiv_operand_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 124.54 0.8 124.84 ;
    END
  END multdiv_operand_b_i[26]
  PIN multdiv_operand_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 75.7 0.8 76 ;
    END
  END multdiv_operand_b_i[27]
  PIN multdiv_operand_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 382.06 0.8 382.36 ;
    END
  END multdiv_operand_b_i[28]
  PIN multdiv_operand_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 333.22 0.8 333.52 ;
    END
  END multdiv_operand_b_i[29]
  PIN multdiv_operand_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 111.22 0.8 111.52 ;
    END
  END multdiv_operand_b_i[2]
  PIN multdiv_operand_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 395.38 262.08 395.68 ;
    END
  END multdiv_operand_b_i[30]
  PIN multdiv_operand_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 337.66 262.08 337.96 ;
    END
  END multdiv_operand_b_i[31]
  PIN multdiv_operand_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 186.7 0.8 187 ;
    END
  END multdiv_operand_b_i[3]
  PIN multdiv_operand_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 204.46 0.8 204.76 ;
    END
  END multdiv_operand_b_i[4]
  PIN multdiv_operand_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 44.62 0.8 44.92 ;
    END
  END multdiv_operand_b_i[5]
  PIN multdiv_operand_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 66.82 0.8 67.12 ;
    END
  END multdiv_operand_b_i[6]
  PIN multdiv_operand_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 120.1 0.8 120.4 ;
    END
  END multdiv_operand_b_i[7]
  PIN multdiv_operand_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 17.98 0.8 18.28 ;
    END
  END multdiv_operand_b_i[8]
  PIN multdiv_operand_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 355.42 0.8 355.72 ;
    END
  END multdiv_operand_b_i[9]
  PIN multdiv_operator_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 350.98 262.08 351.28 ;
    END
  END multdiv_operator_i[0]
  PIN multdiv_operator_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 213.34 262.08 213.64 ;
    END
  END multdiv_operator_i[1]
  PIN multdiv_ready_id_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 328.78 262.08 329.08 ;
    END
  END multdiv_ready_id_i
  PIN multdiv_signed_mode_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 324.34 262.08 324.64 ;
    END
  END multdiv_signed_mode_i[0]
  PIN multdiv_signed_mode_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 333.22 262.08 333.52 ;
    END
  END multdiv_signed_mode_i[1]
  PIN result_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 590.74 0.8 591.04 ;
    END
  END result_ex_o[0]
  PIN result_ex_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 470.86 0.8 471.16 ;
    END
  END result_ex_o[10]
  PIN result_ex_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 506.38 0.8 506.68 ;
    END
  END result_ex_o[11]
  PIN result_ex_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 715.06 0.8 715.36 ;
    END
  END result_ex_o[12]
  PIN result_ex_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 488.62 0.8 488.92 ;
    END
  END result_ex_o[13]
  PIN result_ex_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 741.7 0.8 742 ;
    END
  END result_ex_o[14]
  PIN result_ex_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 528.58 0.8 528.88 ;
    END
  END result_ex_o[15]
  PIN result_ex_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 515.26 0.8 515.56 ;
    END
  END result_ex_o[16]
  PIN result_ex_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 484.18 0.8 484.48 ;
    END
  END result_ex_o[17]
  PIN result_ex_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 701.74 0.8 702.04 ;
    END
  END result_ex_o[18]
  PIN result_ex_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 493.06 0.8 493.36 ;
    END
  END result_ex_o[19]
  PIN result_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 461.98 0.8 462.28 ;
    END
  END result_ex_o[1]
  PIN result_ex_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 510.82 0.8 511.12 ;
    END
  END result_ex_o[20]
  PIN result_ex_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 475.3 0.8 475.6 ;
    END
  END result_ex_o[21]
  PIN result_ex_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 501.94 0.8 502.24 ;
    END
  END result_ex_o[22]
  PIN result_ex_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 692.86 0.8 693.16 ;
    END
  END result_ex_o[23]
  PIN result_ex_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 497.5 0.8 497.8 ;
    END
  END result_ex_o[24]
  PIN result_ex_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 484.18 262.08 484.48 ;
    END
  END result_ex_o[25]
  PIN result_ex_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 457.54 262.08 457.84 ;
    END
  END result_ex_o[26]
  PIN result_ex_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 475.3 262.08 475.6 ;
    END
  END result_ex_o[27]
  PIN result_ex_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 466.42 262.08 466.72 ;
    END
  END result_ex_o[28]
  PIN result_ex_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 564.1 262.08 564.4 ;
    END
  END result_ex_o[29]
  PIN result_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 453.1 262.08 453.4 ;
    END
  END result_ex_o[2]
  PIN result_ex_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 533.02 262.08 533.32 ;
    END
  END result_ex_o[30]
  PIN result_ex_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 524.14 262.08 524.44 ;
    END
  END result_ex_o[31]
  PIN result_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 444.22 262.08 444.52 ;
    END
  END result_ex_o[3]
  PIN result_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 439.78 262.08 440.08 ;
    END
  END result_ex_o[4]
  PIN result_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 448.66 262.08 448.96 ;
    END
  END result_ex_o[5]
  PIN result_ex_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 430.9 262.08 431.2 ;
    END
  END result_ex_o[6]
  PIN result_ex_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 501.94 262.08 502.24 ;
    END
  END result_ex_o[7]
  PIN result_ex_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 493.06 262.08 493.36 ;
    END
  END result_ex_o[8]
  PIN result_ex_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 510.82 262.08 511.12 ;
    END
  END result_ex_o[9]
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  261.28 617.38 262.08 617.68 ;
    END
  END rst_ni
  OBS
    LAYER li1 ;
     RECT  0 0 262.08 782.24 ;
    LAYER met1 ;
     RECT  0 0 262.08 782.24 ;
    LAYER met2 ;
     RECT  0 0 262.08 782.24 ;
    LAYER met3 ;
     RECT  0 0 262.08 782.24 ;
    LAYER met4 ;
     RECT  0 0 262.08 782.24 ;
    LAYER met5 ;
     RECT  0 0 262.08 782.24 ;
  END
END ibex_ex_block
END LIBRARY
